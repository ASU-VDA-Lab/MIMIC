module real_aes_12287_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_0), .A2(n_214), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_0), .A2(n_214), .B1(n_613), .B2(n_1403), .Y(n_1402) );
INVxp33_ASAP7_75t_L g1438 ( .A(n_1), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_1), .A2(n_26), .B1(n_427), .B2(n_1462), .Y(n_1461) );
AO221x1_ASAP7_75t_L g1218 ( .A1(n_2), .A2(n_150), .B1(n_1185), .B2(n_1219), .C(n_1221), .Y(n_1218) );
OAI222xp33_ASAP7_75t_L g651 ( .A1(n_3), .A2(n_34), .B1(n_148), .B2(n_652), .C1(n_654), .C2(n_656), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_3), .A2(n_148), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g1141 ( .A(n_4), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_5), .A2(n_167), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_5), .A2(n_122), .B1(n_282), .B2(n_330), .C(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_6), .Y(n_263) );
AND2x2_ASAP7_75t_L g289 ( .A(n_6), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_6), .B(n_189), .Y(n_305) );
INVx1_ASAP7_75t_L g362 ( .A(n_6), .Y(n_362) );
OA22x2_ASAP7_75t_L g276 ( .A1(n_7), .A2(n_277), .B1(n_457), .B2(n_458), .Y(n_276) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_7), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_7), .A2(n_101), .B1(n_1185), .B2(n_1189), .Y(n_1210) );
INVxp67_ASAP7_75t_L g1444 ( .A(n_8), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_8), .A2(n_66), .B1(n_371), .B2(n_427), .Y(n_1468) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_9), .A2(n_89), .B1(n_387), .B2(n_428), .Y(n_592) );
INVx1_ASAP7_75t_L g605 ( .A(n_9), .Y(n_605) );
OAI332xp33_ASAP7_75t_L g321 ( .A1(n_10), .A2(n_322), .A3(n_331), .B1(n_341), .B2(n_345), .B3(n_352), .C1(n_358), .C2(n_363), .Y(n_321) );
INVx1_ASAP7_75t_L g450 ( .A(n_10), .Y(n_450) );
INVxp33_ASAP7_75t_L g839 ( .A(n_11), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_11), .A2(n_133), .B1(n_452), .B2(n_594), .C(n_643), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_12), .A2(n_93), .B1(n_500), .B2(n_1013), .Y(n_1012) );
INVxp67_ASAP7_75t_SL g1039 ( .A(n_12), .Y(n_1039) );
INVx1_ASAP7_75t_L g1017 ( .A(n_13), .Y(n_1017) );
AO221x2_ASAP7_75t_L g1241 ( .A1(n_14), .A2(n_166), .B1(n_1219), .B2(n_1242), .C(n_1244), .Y(n_1241) );
INVx1_ASAP7_75t_L g757 ( .A(n_15), .Y(n_757) );
OR2x2_ASAP7_75t_L g394 ( .A(n_16), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g403 ( .A(n_16), .Y(n_403) );
INVx1_ASAP7_75t_L g888 ( .A(n_17), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_18), .A2(n_235), .B1(n_962), .B2(n_964), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_18), .A2(n_235), .B1(n_982), .B2(n_983), .Y(n_981) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_19), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_20), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_21), .A2(n_129), .B1(n_427), .B2(n_442), .Y(n_1004) );
INVxp33_ASAP7_75t_SL g1027 ( .A(n_21), .Y(n_1027) );
INVx1_ASAP7_75t_L g288 ( .A(n_22), .Y(n_288) );
OR2x2_ASAP7_75t_L g304 ( .A(n_22), .B(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g344 ( .A(n_22), .Y(n_344) );
BUFx2_ASAP7_75t_L g516 ( .A(n_22), .Y(n_516) );
INVx1_ASAP7_75t_L g1015 ( .A(n_23), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_24), .A2(n_164), .B1(n_316), .B2(n_319), .C(n_530), .Y(n_1127) );
OAI22xp33_ASAP7_75t_SL g1151 ( .A1(n_24), .A2(n_164), .B1(n_661), .B2(n_887), .Y(n_1151) );
AOI22xp33_ASAP7_75t_SL g1400 ( .A1(n_25), .A2(n_92), .B1(n_387), .B2(n_580), .Y(n_1400) );
INVxp67_ASAP7_75t_L g1413 ( .A(n_25), .Y(n_1413) );
INVxp33_ASAP7_75t_L g1434 ( .A(n_26), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_27), .A2(n_153), .B1(n_543), .B2(n_609), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_27), .A2(n_153), .B1(n_780), .B2(n_1109), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_28), .A2(n_139), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_28), .A2(n_130), .B1(n_611), .B2(n_613), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_29), .A2(n_105), .B1(n_342), .B2(n_527), .C(n_983), .Y(n_1084) );
INVx1_ASAP7_75t_L g1106 ( .A(n_29), .Y(n_1106) );
INVx1_ASAP7_75t_L g509 ( .A(n_30), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_31), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_32), .A2(n_172), .B1(n_475), .B2(n_476), .C(n_479), .Y(n_474) );
INVxp33_ASAP7_75t_SL g537 ( .A(n_32), .Y(n_537) );
INVxp33_ASAP7_75t_L g901 ( .A(n_33), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_33), .A2(n_36), .B1(n_982), .B2(n_983), .Y(n_993) );
INVx1_ASAP7_75t_L g694 ( .A(n_34), .Y(n_694) );
INVxp33_ASAP7_75t_L g1124 ( .A(n_35), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_35), .A2(n_37), .B1(n_452), .B2(n_636), .C(n_1147), .Y(n_1146) );
INVxp67_ASAP7_75t_L g919 ( .A(n_36), .Y(n_919) );
INVxp33_ASAP7_75t_L g1122 ( .A(n_37), .Y(n_1122) );
INVx1_ASAP7_75t_L g860 ( .A(n_38), .Y(n_860) );
INVxp33_ASAP7_75t_SL g1125 ( .A(n_39), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_39), .A2(n_232), .B1(n_970), .B2(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1139 ( .A(n_40), .Y(n_1139) );
INVx1_ASAP7_75t_L g1222 ( .A(n_41), .Y(n_1222) );
INVx1_ASAP7_75t_L g1018 ( .A(n_42), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_43), .A2(n_184), .B1(n_560), .B2(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g817 ( .A(n_43), .Y(n_817) );
INVx1_ASAP7_75t_L g473 ( .A(n_44), .Y(n_473) );
INVx1_ASAP7_75t_L g1098 ( .A(n_45), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_45), .A2(n_137), .B1(n_1109), .B2(n_1113), .Y(n_1112) );
INVxp33_ASAP7_75t_L g953 ( .A(n_46), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_46), .A2(n_119), .B1(n_962), .B2(n_972), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_47), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_48), .A2(n_215), .B1(n_1398), .B2(n_1399), .Y(n_1397) );
INVxp33_ASAP7_75t_L g1415 ( .A(n_48), .Y(n_1415) );
OAI222xp33_ASAP7_75t_L g658 ( .A1(n_49), .A2(n_125), .B1(n_197), .B2(n_412), .C1(n_659), .C2(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g669 ( .A(n_49), .Y(n_669) );
INVxp67_ASAP7_75t_L g950 ( .A(n_50), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_50), .A2(n_70), .B1(n_642), .B2(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g912 ( .A(n_51), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_52), .A2(n_186), .B1(n_280), .B2(n_291), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_52), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_53), .A2(n_126), .B1(n_427), .B2(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g686 ( .A(n_53), .Y(n_686) );
INVxp33_ASAP7_75t_SL g704 ( .A(n_54), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_54), .A2(n_234), .B1(n_737), .B2(n_747), .C(n_749), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_55), .A2(n_82), .B1(n_639), .B2(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g675 ( .A(n_55), .Y(n_675) );
INVx1_ASAP7_75t_L g1223 ( .A(n_56), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_57), .Y(n_567) );
INVxp67_ASAP7_75t_L g1442 ( .A(n_58), .Y(n_1442) );
AOI221xp5_ASAP7_75t_L g1467 ( .A1(n_58), .A2(n_168), .B1(n_479), .B2(n_643), .C(n_885), .Y(n_1467) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_59), .B(n_556), .Y(n_555) );
INVxp33_ASAP7_75t_L g907 ( .A(n_60), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_60), .A2(n_75), .B1(n_543), .B2(n_986), .Y(n_992) );
INVx1_ASAP7_75t_L g502 ( .A(n_61), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_62), .Y(n_1093) );
AO221x1_ASAP7_75t_L g1199 ( .A1(n_63), .A2(n_107), .B1(n_1185), .B2(n_1189), .C(n_1200), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_64), .A2(n_134), .B1(n_298), .B2(n_303), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_64), .Y(n_444) );
INVx1_ASAP7_75t_L g1247 ( .A(n_65), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1446 ( .A(n_66), .Y(n_1446) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_67), .A2(n_218), .B1(n_657), .B2(n_738), .C(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g804 ( .A(n_67), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g1050 ( .A(n_68), .B(n_1051), .Y(n_1050) );
INVxp33_ASAP7_75t_L g1130 ( .A(n_69), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_69), .A2(n_207), .B1(n_879), .B2(n_1156), .Y(n_1155) );
INVxp33_ASAP7_75t_L g946 ( .A(n_70), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_71), .A2(n_138), .B1(n_475), .B2(n_504), .C(n_507), .Y(n_503) );
INVxp33_ASAP7_75t_SL g525 ( .A(n_71), .Y(n_525) );
AO221x1_ASAP7_75t_L g1192 ( .A1(n_72), .A2(n_156), .B1(n_1185), .B2(n_1189), .C(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g395 ( .A(n_73), .Y(n_395) );
INVx1_ASAP7_75t_L g438 ( .A(n_73), .Y(n_438) );
INVx1_ASAP7_75t_L g498 ( .A(n_74), .Y(n_498) );
INVxp33_ASAP7_75t_L g916 ( .A(n_75), .Y(n_916) );
INVx1_ASAP7_75t_L g926 ( .A(n_76), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_76), .A2(n_175), .B1(n_940), .B2(n_942), .Y(n_939) );
INVx1_ASAP7_75t_L g1046 ( .A(n_77), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_78), .Y(n_1058) );
INVx1_ASAP7_75t_L g1197 ( .A(n_79), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_80), .A2(n_199), .B1(n_481), .B2(n_483), .Y(n_480) );
INVxp67_ASAP7_75t_L g545 ( .A(n_80), .Y(n_545) );
INVx1_ASAP7_75t_L g1378 ( .A(n_81), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_81), .A2(n_182), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
INVx1_ASAP7_75t_L g671 ( .A(n_82), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g1439 ( .A1(n_83), .A2(n_110), .B1(n_530), .B2(n_531), .C(n_842), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1464 ( .A1(n_83), .A2(n_110), .B1(n_1007), .B2(n_1465), .Y(n_1464) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_84), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_84), .A2(n_194), .B1(n_475), .B2(n_479), .C(n_562), .Y(n_877) );
INVxp33_ASAP7_75t_SL g835 ( .A(n_85), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_85), .A2(n_102), .B1(n_762), .B2(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g1059 ( .A(n_86), .Y(n_1059) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_86), .A2(n_160), .B1(n_1079), .B2(n_1081), .C(n_1082), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_87), .A2(n_145), .B1(n_969), .B2(n_970), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_87), .A2(n_145), .B1(n_986), .B2(n_988), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_88), .A2(n_206), .B1(n_1185), .B2(n_1189), .Y(n_1215) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_89), .A2(n_596), .B(n_597), .C(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g494 ( .A(n_90), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_90), .A2(n_209), .B1(n_530), .B2(n_531), .C(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g1056 ( .A(n_91), .Y(n_1056) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_91), .A2(n_147), .B1(n_282), .B2(n_1071), .C(n_1072), .Y(n_1070) );
INVxp33_ASAP7_75t_L g1412 ( .A(n_92), .Y(n_1412) );
INVxp33_ASAP7_75t_L g1031 ( .A(n_93), .Y(n_1031) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_94), .Y(n_775) );
INVx1_ASAP7_75t_L g1005 ( .A(n_95), .Y(n_1005) );
OAI22xp33_ASAP7_75t_SL g794 ( .A1(n_96), .A2(n_195), .B1(n_561), .B2(n_741), .Y(n_794) );
INVx1_ASAP7_75t_L g821 ( .A(n_96), .Y(n_821) );
INVx1_ASAP7_75t_L g856 ( .A(n_97), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_97), .A2(n_159), .B1(n_427), .B2(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1137 ( .A(n_98), .Y(n_1137) );
INVx1_ASAP7_75t_L g1202 ( .A(n_99), .Y(n_1202) );
AO22x2_ASAP7_75t_L g1367 ( .A1(n_99), .A2(n_1202), .B1(n_1368), .B2(n_1417), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_99), .A2(n_1424), .B1(n_1428), .B2(n_1471), .Y(n_1423) );
INVx1_ASAP7_75t_L g255 ( .A(n_100), .Y(n_255) );
INVxp33_ASAP7_75t_SL g840 ( .A(n_102), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_103), .Y(n_589) );
INVx1_ASAP7_75t_L g718 ( .A(n_104), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_104), .A2(n_193), .B1(n_737), .B2(n_738), .C(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g1107 ( .A(n_105), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_106), .A2(n_190), .B1(n_1173), .B2(n_1181), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_108), .A2(n_144), .B1(n_583), .B2(n_780), .C(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g824 ( .A(n_108), .Y(n_824) );
INVx1_ASAP7_75t_L g1201 ( .A(n_109), .Y(n_1201) );
INVx1_ASAP7_75t_L g1449 ( .A(n_111), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_112), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_113), .Y(n_783) );
INVx1_ASAP7_75t_L g1380 ( .A(n_114), .Y(n_1380) );
INVx1_ASAP7_75t_L g758 ( .A(n_115), .Y(n_758) );
INVx1_ASAP7_75t_L g461 ( .A(n_116), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_116), .A2(n_173), .B1(n_1185), .B2(n_1189), .Y(n_1184) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_117), .A2(n_170), .B1(n_642), .B2(n_643), .C(n_644), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_117), .A2(n_126), .B1(n_681), .B2(n_683), .C(n_685), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_118), .A2(n_246), .B1(n_1173), .B2(n_1181), .Y(n_1216) );
INVxp67_ASAP7_75t_L g933 ( .A(n_119), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_120), .A2(n_205), .B1(n_308), .B2(n_315), .C(n_319), .Y(n_307) );
OAI222xp33_ASAP7_75t_L g406 ( .A1(n_120), .A2(n_134), .B1(n_205), .B2(n_407), .C1(n_412), .C2(n_414), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_121), .A2(n_176), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g1028 ( .A1(n_121), .A2(n_176), .B1(n_319), .B2(n_530), .C(n_531), .Y(n_1028) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_122), .A2(n_583), .B(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_123), .A2(n_127), .B1(n_443), .B2(n_657), .Y(n_1388) );
AOI22xp33_ASAP7_75t_SL g1401 ( .A1(n_123), .A2(n_127), .B1(n_330), .B2(n_987), .Y(n_1401) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_124), .A2(n_136), .B1(n_634), .B2(n_636), .C(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g673 ( .A(n_124), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_125), .Y(n_677) );
INVx1_ASAP7_75t_L g1245 ( .A(n_128), .Y(n_1245) );
INVxp33_ASAP7_75t_L g1023 ( .A(n_129), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_130), .A2(n_142), .B1(n_445), .B2(n_564), .Y(n_563) );
INVxp33_ASAP7_75t_SL g1372 ( .A(n_131), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_131), .A2(n_143), .B1(n_613), .B2(n_720), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_132), .A2(n_201), .B1(n_527), .B2(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_132), .A2(n_216), .B1(n_560), .B2(n_761), .Y(n_760) );
INVxp33_ASAP7_75t_L g837 ( .A(n_133), .Y(n_837) );
INVx1_ASAP7_75t_L g1455 ( .A(n_135), .Y(n_1455) );
INVx1_ASAP7_75t_L g679 ( .A(n_136), .Y(n_679) );
INVx1_ASAP7_75t_L g1096 ( .A(n_137), .Y(n_1096) );
INVxp33_ASAP7_75t_SL g523 ( .A(n_138), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_139), .A2(n_142), .B1(n_522), .B2(n_609), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_140), .A2(n_452), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g604 ( .A(n_140), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_141), .Y(n_650) );
INVxp67_ASAP7_75t_SL g1375 ( .A(n_143), .Y(n_1375) );
INVx1_ASAP7_75t_L g826 ( .A(n_144), .Y(n_826) );
INVx1_ASAP7_75t_L g1019 ( .A(n_146), .Y(n_1019) );
INVx1_ASAP7_75t_L g1063 ( .A(n_147), .Y(n_1063) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_149), .A2(n_245), .B1(n_316), .B2(n_530), .C(n_842), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_149), .A2(n_245), .B1(n_661), .B2(n_887), .Y(n_886) );
INVxp33_ASAP7_75t_SL g1381 ( .A(n_151), .Y(n_1381) );
AOI22xp33_ASAP7_75t_SL g1392 ( .A1(n_151), .A2(n_174), .B1(n_330), .B2(n_987), .Y(n_1392) );
INVx1_ASAP7_75t_L g712 ( .A(n_152), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g1115 ( .A(n_154), .B(n_1116), .Y(n_1115) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_155), .Y(n_788) );
INVx1_ASAP7_75t_L g830 ( .A(n_156), .Y(n_830) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_157), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_157), .B(n_255), .Y(n_1180) );
AND3x2_ASAP7_75t_L g1188 ( .A(n_157), .B(n_255), .C(n_1177), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_158), .Y(n_575) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_159), .Y(n_848) );
INVx1_ASAP7_75t_L g1060 ( .A(n_160), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_161), .A2(n_200), .B1(n_564), .B2(n_570), .C(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g599 ( .A(n_161), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_162), .Y(n_346) );
INVx2_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
XNOR2x2_ASAP7_75t_L g700 ( .A(n_165), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g618 ( .A(n_167), .Y(n_618) );
INVxp33_ASAP7_75t_L g1447 ( .A(n_168), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_169), .Y(n_353) );
INVx1_ASAP7_75t_L g688 ( .A(n_170), .Y(n_688) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_171), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_171), .A2(n_222), .B1(n_475), .B2(n_479), .C(n_1154), .Y(n_1153) );
INVxp67_ASAP7_75t_L g541 ( .A(n_172), .Y(n_541) );
INVxp33_ASAP7_75t_SL g1373 ( .A(n_174), .Y(n_1373) );
INVx1_ASAP7_75t_L g921 ( .A(n_175), .Y(n_921) );
INVx1_ASAP7_75t_L g1450 ( .A(n_177), .Y(n_1450) );
INVx1_ASAP7_75t_L g1177 ( .A(n_178), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1010 ( .A1(n_179), .A2(n_239), .B1(n_443), .B2(n_479), .C(n_1011), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1036 ( .A(n_179), .Y(n_1036) );
INVx1_ASAP7_75t_L g715 ( .A(n_180), .Y(n_715) );
INVx1_ASAP7_75t_L g706 ( .A(n_181), .Y(n_706) );
INVx1_ASAP7_75t_L g1376 ( .A(n_182), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_183), .Y(n_323) );
INVx1_ASAP7_75t_L g819 ( .A(n_184), .Y(n_819) );
INVx1_ASAP7_75t_L g863 ( .A(n_185), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_186), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_187), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_188), .Y(n_799) );
INVx1_ASAP7_75t_L g270 ( .A(n_189), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_189), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g1209 ( .A1(n_191), .A2(n_208), .B1(n_1173), .B2(n_1181), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_192), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_193), .A2(n_196), .B1(n_720), .B2(n_722), .Y(n_719) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_194), .Y(n_855) );
INVx1_ASAP7_75t_L g815 ( .A(n_195), .Y(n_815) );
INVx1_ASAP7_75t_L g743 ( .A(n_196), .Y(n_743) );
INVx1_ASAP7_75t_L g668 ( .A(n_197), .Y(n_668) );
INVx1_ASAP7_75t_L g1194 ( .A(n_198), .Y(n_1194) );
INVxp67_ASAP7_75t_L g535 ( .A(n_199), .Y(n_535) );
INVx1_ASAP7_75t_L g623 ( .A(n_200), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_201), .A2(n_223), .B1(n_477), .B2(n_564), .Y(n_763) );
INVxp33_ASAP7_75t_L g1437 ( .A(n_202), .Y(n_1437) );
AOI221xp5_ASAP7_75t_L g1460 ( .A1(n_202), .A2(n_203), .B1(n_636), .B2(n_637), .C(n_972), .Y(n_1460) );
INVxp33_ASAP7_75t_L g1435 ( .A(n_203), .Y(n_1435) );
INVx1_ASAP7_75t_L g861 ( .A(n_204), .Y(n_861) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_207), .Y(n_1134) );
INVx1_ASAP7_75t_L g495 ( .A(n_209), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_210), .Y(n_335) );
INVx1_ASAP7_75t_L g1454 ( .A(n_211), .Y(n_1454) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_212), .A2(n_248), .B1(n_371), .B2(n_637), .C(n_972), .Y(n_1003) );
INVxp33_ASAP7_75t_L g1026 ( .A(n_212), .Y(n_1026) );
INVx1_ASAP7_75t_L g1178 ( .A(n_213), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_213), .B(n_1176), .Y(n_1183) );
INVxp67_ASAP7_75t_SL g1406 ( .A(n_215), .Y(n_1406) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_216), .Y(n_729) );
INVx1_ASAP7_75t_L g489 ( .A(n_217), .Y(n_489) );
INVx1_ASAP7_75t_L g813 ( .A(n_218), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_219), .Y(n_1457) );
INVx1_ASAP7_75t_L g1158 ( .A(n_220), .Y(n_1158) );
AO22x1_ASAP7_75t_L g1235 ( .A1(n_221), .A2(n_233), .B1(n_1189), .B2(n_1236), .Y(n_1235) );
INVxp33_ASAP7_75t_L g1131 ( .A(n_222), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_223), .Y(n_727) );
INVx1_ASAP7_75t_L g1062 ( .A(n_224), .Y(n_1062) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_224), .A2(n_1075), .B(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g1142 ( .A(n_225), .Y(n_1142) );
INVx2_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_227), .Y(n_1055) );
AO22x1_ASAP7_75t_L g1237 ( .A1(n_228), .A2(n_238), .B1(n_1173), .B2(n_1181), .Y(n_1237) );
XNOR2x1_ASAP7_75t_L g629 ( .A(n_229), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g486 ( .A(n_230), .Y(n_486) );
XNOR2x2_ASAP7_75t_L g769 ( .A(n_231), .B(n_770), .Y(n_769) );
INVxp33_ASAP7_75t_L g1120 ( .A(n_232), .Y(n_1120) );
INVxp33_ASAP7_75t_SL g708 ( .A(n_234), .Y(n_708) );
OAI22x1_ASAP7_75t_SL g895 ( .A1(n_236), .A2(n_896), .B1(n_994), .B2(n_995), .Y(n_895) );
INVx1_ASAP7_75t_L g994 ( .A(n_236), .Y(n_994) );
INVx1_ASAP7_75t_L g710 ( .A(n_237), .Y(n_710) );
INVxp33_ASAP7_75t_SL g1033 ( .A(n_239), .Y(n_1033) );
INVx1_ASAP7_75t_L g864 ( .A(n_240), .Y(n_864) );
BUFx3_ASAP7_75t_L g376 ( .A(n_241), .Y(n_376) );
INVx1_ASAP7_75t_L g383 ( .A(n_241), .Y(n_383) );
BUFx3_ASAP7_75t_L g378 ( .A(n_242), .Y(n_378) );
INVx1_ASAP7_75t_L g389 ( .A(n_242), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_243), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_244), .Y(n_776) );
XNOR2xp5_ASAP7_75t_L g1429 ( .A(n_247), .B(n_1430), .Y(n_1429) );
INVxp33_ASAP7_75t_L g1024 ( .A(n_248), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_271), .B(n_1163), .Y(n_249) );
INVx3_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_253), .B(n_259), .Y(n_1422) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_SL g1427 ( .A(n_254), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_254), .B(n_256), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_256), .B(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g956 ( .A(n_261), .B(n_516), .Y(n_956) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g615 ( .A(n_262), .B(n_270), .Y(n_615) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g342 ( .A(n_263), .B(n_343), .Y(n_342) );
INVx8_ASAP7_75t_L g952 ( .A(n_264), .Y(n_952) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
OR2x2_ASAP7_75t_L g303 ( .A(n_265), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g334 ( .A(n_265), .Y(n_334) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_265), .Y(n_354) );
INVx2_ASAP7_75t_SL g550 ( .A(n_265), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_265), .A2(n_337), .B1(n_575), .B2(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g687 ( .A(n_265), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_265), .A2(n_337), .B1(n_650), .B2(n_694), .Y(n_693) );
OR2x6_ASAP7_75t_L g955 ( .A(n_265), .B(n_945), .Y(n_955) );
INVx2_ASAP7_75t_SL g1453 ( .A(n_265), .Y(n_1453) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
INVx1_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
AND2x4_ASAP7_75t_L g302 ( .A(n_267), .B(n_296), .Y(n_302) );
INVx1_ASAP7_75t_L g340 ( .A(n_267), .Y(n_340) );
AND2x2_ASAP7_75t_L g367 ( .A(n_267), .B(n_268), .Y(n_367) );
INVx1_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
INVx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
INVx1_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_268), .B(n_284), .Y(n_327) );
INVx1_ASAP7_75t_L g339 ( .A(n_268), .Y(n_339) );
AND2x4_ASAP7_75t_L g941 ( .A(n_269), .B(n_313), .Y(n_941) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g942 ( .A(n_270), .B(n_602), .Y(n_942) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_270), .B(n_602), .Y(n_1410) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_696), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_627), .B1(n_628), .B2(n_695), .Y(n_272) );
INVx1_ASAP7_75t_L g695 ( .A(n_273), .Y(n_695) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_459), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g457 ( .A(n_277), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_306), .C(n_368), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_297), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g596 ( .A(n_281), .Y(n_596) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_287), .Y(n_281) );
AND2x2_ASAP7_75t_L g528 ( .A(n_282), .B(n_287), .Y(n_528) );
AND2x2_ASAP7_75t_L g672 ( .A(n_282), .B(n_287), .Y(n_672) );
AND2x2_ASAP7_75t_L g709 ( .A(n_282), .B(n_287), .Y(n_709) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_282), .B(n_287), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_283), .Y(n_609) );
INVx1_ASAP7_75t_L g682 ( .A(n_283), .Y(n_682) );
INVx1_ASAP7_75t_L g691 ( .A(n_283), .Y(n_691) );
AND2x4_ASAP7_75t_L g944 ( .A(n_283), .B(n_945), .Y(n_944) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_283), .Y(n_987) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_283), .B(n_289), .Y(n_1097) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x6_ASAP7_75t_L g292 ( .A(n_287), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g299 ( .A(n_287), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g364 ( .A(n_287), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g521 ( .A(n_287), .B(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g526 ( .A(n_287), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g619 ( .A(n_287), .B(n_613), .Y(n_619) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g359 ( .A(n_288), .Y(n_359) );
INVx2_ASAP7_75t_L g1092 ( .A(n_289), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_289), .B(n_612), .Y(n_1094) );
INVx1_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
INVx1_ASAP7_75t_L g361 ( .A(n_290), .Y(n_361) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_292), .A2(n_502), .B1(n_520), .B2(n_523), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_292), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_292), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_292), .A2(n_521), .B1(n_782), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_292), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_292), .A2(n_836), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_292), .A2(n_1120), .B1(n_1121), .B2(n_1122), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_292), .A2(n_521), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_293), .B(n_314), .Y(n_320) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_294), .Y(n_613) );
BUFx2_ASAP7_75t_L g625 ( .A(n_294), .Y(n_625) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_294), .Y(n_724) );
BUFx3_ASAP7_75t_L g732 ( .A(n_294), .Y(n_732) );
AND2x4_ASAP7_75t_L g936 ( .A(n_294), .B(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g984 ( .A(n_294), .Y(n_984) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_299), .A2(n_364), .B1(n_604), .B2(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g350 ( .A(n_300), .Y(n_350) );
INVx2_ASAP7_75t_L g684 ( .A(n_300), .Y(n_684) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g522 ( .A(n_301), .Y(n_522) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_301), .Y(n_544) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx1_ASAP7_75t_L g949 ( .A(n_302), .Y(n_949) );
INVx1_ASAP7_75t_L g1101 ( .A(n_302), .Y(n_1101) );
AND2x4_ASAP7_75t_L g513 ( .A(n_303), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g598 ( .A(n_303), .Y(n_598) );
INVx3_ASAP7_75t_L g314 ( .A(n_304), .Y(n_314) );
INVx1_ASAP7_75t_L g1069 ( .A(n_305), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_321), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g530 ( .A(n_309), .Y(n_530) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2x1_ASAP7_75t_SL g310 ( .A(n_311), .B(n_314), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g1079 ( .A(n_311), .B(n_1080), .Y(n_1079) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_313), .Y(n_622) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_314), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g600 ( .A(n_314), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g621 ( .A(n_314), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g624 ( .A(n_314), .B(n_625), .Y(n_624) );
BUFx4f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_316), .Y(n_531) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x6_ASAP7_75t_L g1081 ( .A(n_318), .B(n_1068), .Y(n_1081) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g532 ( .A(n_320), .Y(n_532) );
BUFx2_ASAP7_75t_L g842 ( .A(n_320), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_328), .B2(n_329), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_323), .A2(n_335), .B1(n_430), .B2(n_433), .C(n_436), .Y(n_429) );
INVx2_ASAP7_75t_L g540 ( .A(n_324), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_324), .A2(n_1137), .B1(n_1138), .B2(n_1139), .Y(n_1136) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g726 ( .A(n_325), .Y(n_726) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g859 ( .A(n_326), .Y(n_859) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g349 ( .A(n_327), .Y(n_349) );
INVx1_ASAP7_75t_L g812 ( .A(n_327), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_328), .A2(n_332), .B1(n_420), .B2(n_426), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_329), .A2(n_853), .B1(n_855), .B2(n_856), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_329), .A2(n_858), .B1(n_860), .B2(n_861), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_329), .A2(n_1442), .B1(n_1443), .B2(n_1444), .Y(n_1441) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g728 ( .A(n_330), .Y(n_728) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_330), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_335), .B2(n_336), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_333), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_534) );
OAI22xp33_ASAP7_75t_L g803 ( .A1(n_333), .A2(n_775), .B1(n_804), .B2(n_805), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_333), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_818) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
BUFx3_ASAP7_75t_L g551 ( .A(n_337), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_337), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_685) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g808 ( .A(n_339), .B(n_340), .Y(n_808) );
INVx1_ASAP7_75t_L g602 ( .A(n_340), .Y(n_602) );
OAI33xp33_ASAP7_75t_L g533 ( .A1(n_341), .A2(n_534), .A3(n_538), .B1(n_546), .B2(n_547), .B3(n_552), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_341), .A2(n_714), .B1(n_725), .B2(n_733), .Y(n_713) );
OAI33xp33_ASAP7_75t_L g802 ( .A1(n_341), .A2(n_552), .A3(n_803), .B1(n_809), .B2(n_814), .B3(n_818), .Y(n_802) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_341), .Y(n_844) );
OAI33xp33_ASAP7_75t_L g1029 ( .A1(n_341), .A2(n_733), .A3(n_1030), .B1(n_1035), .B2(n_1040), .B3(n_1043), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1440 ( .A1(n_341), .A2(n_733), .A3(n_1441), .B1(n_1445), .B2(n_1448), .B3(n_1451), .Y(n_1440) );
OR2x6_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g945 ( .A(n_343), .Y(n_945) );
INVx2_ASAP7_75t_L g456 ( .A(n_344), .Y(n_456) );
BUFx2_ASAP7_75t_L g665 ( .A(n_344), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_350), .B2(n_351), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_346), .A2(n_355), .B1(n_385), .B2(n_390), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_347), .A2(n_715), .B1(n_716), .B2(n_718), .C(n_719), .Y(n_714) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g692 ( .A(n_350), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_350), .A2(n_1443), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_351), .A2(n_353), .B1(n_371), .B2(n_379), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_354), .B1(n_355), .B2(n_356), .Y(n_352) );
INVx1_ASAP7_75t_L g847 ( .A(n_354), .Y(n_847) );
BUFx2_ASAP7_75t_L g1032 ( .A(n_354), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_356), .A2(n_846), .B1(n_863), .B2(n_864), .Y(n_862) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g536 ( .A(n_357), .Y(n_536) );
INVx2_ASAP7_75t_L g820 ( .A(n_357), .Y(n_820) );
INVx6_ASAP7_75t_L g553 ( .A(n_358), .Y(n_553) );
INVx5_ASAP7_75t_L g734 ( .A(n_358), .Y(n_734) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g1077 ( .A(n_360), .Y(n_1077) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g938 ( .A(n_361), .Y(n_938) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_364), .A2(n_553), .B1(n_614), .B2(n_679), .C1(n_680), .C2(n_689), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_365), .B(n_1088), .Y(n_1087) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g527 ( .A(n_366), .Y(n_527) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_367), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_406), .A3(n_418), .B(n_454), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_384), .B(n_394), .C(n_396), .Y(n_369) );
INVx4_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g568 ( .A(n_372), .Y(n_568) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g482 ( .A(n_373), .Y(n_482) );
INVx2_ASAP7_75t_L g506 ( .A(n_373), .Y(n_506) );
INVx1_ASAP7_75t_L g579 ( .A(n_373), .Y(n_579) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_373), .Y(n_647) );
INVx2_ASAP7_75t_SL g881 ( .A(n_373), .Y(n_881) );
INVx2_ASAP7_75t_L g906 ( .A(n_373), .Y(n_906) );
INVx1_ASAP7_75t_L g963 ( .A(n_373), .Y(n_963) );
INVx6_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g413 ( .A(n_374), .B(n_400), .Y(n_413) );
BUFx2_ASAP7_75t_L g594 ( .A(n_374), .Y(n_594) );
AND2x4_ASAP7_75t_L g913 ( .A(n_374), .B(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g1014 ( .A(n_374), .Y(n_1014) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g388 ( .A(n_376), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g393 ( .A(n_376), .B(n_378), .Y(n_393) );
INVx1_ASAP7_75t_L g411 ( .A(n_377), .Y(n_411) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g382 ( .A(n_378), .B(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_382), .Y(n_446) );
INVx2_ASAP7_75t_L g492 ( .A(n_382), .Y(n_492) );
INVx1_ASAP7_75t_L g501 ( .A(n_382), .Y(n_501) );
INVx1_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_387), .Y(n_1109) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_388), .Y(n_478) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_388), .Y(n_562) );
INVx2_ASAP7_75t_SL g584 ( .A(n_388), .Y(n_584) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_388), .Y(n_642) );
BUFx2_ASAP7_75t_L g655 ( .A(n_388), .Y(n_655) );
BUFx2_ASAP7_75t_L g885 ( .A(n_388), .Y(n_885) );
AND2x6_ASAP7_75t_L g908 ( .A(n_388), .B(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_388), .Y(n_1154) );
INVx1_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_391), .Y(n_920) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g471 ( .A(n_392), .B(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g475 ( .A(n_392), .Y(n_475) );
INVx2_ASAP7_75t_SL g635 ( .A(n_392), .Y(n_635) );
AND2x4_ASAP7_75t_L g648 ( .A(n_392), .B(n_573), .Y(n_648) );
BUFx4f_ASAP7_75t_L g972 ( .A(n_392), .Y(n_972) );
INVx1_ASAP7_75t_L g1148 ( .A(n_392), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_393), .Y(n_405) );
INVx2_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
OR2x2_ASAP7_75t_L g488 ( .A(n_394), .B(n_423), .Y(n_488) );
OR2x2_ASAP7_75t_L g491 ( .A(n_394), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g401 ( .A(n_395), .Y(n_401) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_397), .A2(n_469), .B1(n_473), .B2(n_474), .C(n_480), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_397), .A2(n_864), .B1(n_875), .B2(n_877), .C(n_878), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_397), .A2(n_471), .B1(n_1010), .B2(n_1012), .C(n_1015), .Y(n_1009) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_397), .A2(n_469), .B1(n_1142), .B2(n_1153), .C(n_1155), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1466 ( .A1(n_397), .A2(n_1455), .B1(n_1467), .B2(n_1468), .C(n_1469), .Y(n_1466) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_404), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g414 ( .A(n_399), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g408 ( .A(n_400), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g496 ( .A(n_400), .B(n_416), .Y(n_496) );
BUFx2_ASAP7_75t_L g573 ( .A(n_400), .Y(n_573) );
AND2x4_ASAP7_75t_L g660 ( .A(n_400), .B(n_409), .Y(n_660) );
AND2x4_ASAP7_75t_L g662 ( .A(n_400), .B(n_416), .Y(n_662) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AND2x4_ASAP7_75t_L g453 ( .A(n_402), .B(n_438), .Y(n_453) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g437 ( .A(n_403), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g905 ( .A(n_403), .Y(n_905) );
INVx1_ASAP7_75t_L g910 ( .A(n_403), .Y(n_910) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_403), .Y(n_915) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_404), .Y(n_643) );
INVx1_ASAP7_75t_L g790 ( .A(n_404), .Y(n_790) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g929 ( .A(n_405), .B(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g967 ( .A(n_405), .Y(n_967) );
BUFx6f_ASAP7_75t_L g1391 ( .A(n_405), .Y(n_1391) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_408), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_408), .A2(n_496), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_408), .Y(n_1007) );
INVxp67_ASAP7_75t_L g570 ( .A(n_409), .Y(n_570) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g925 ( .A(n_411), .Y(n_925) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g515 ( .A(n_413), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g571 ( .A(n_416), .Y(n_571) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x6_ASAP7_75t_L g927 ( .A(n_417), .B(n_910), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_429), .B1(n_439), .B2(n_447), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_420), .A2(n_590), .B1(n_1089), .B2(n_1093), .C(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g449 ( .A(n_422), .Y(n_449) );
INVx2_ASAP7_75t_L g560 ( .A(n_422), .Y(n_560) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g752 ( .A(n_423), .Y(n_752) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AND2x2_ASAP7_75t_L g432 ( .A(n_424), .B(n_425), .Y(n_432) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
BUFx3_ASAP7_75t_L g780 ( .A(n_428), .Y(n_780) );
INVx1_ASAP7_75t_L g793 ( .A(n_428), .Y(n_793) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_430), .A2(n_448), .B1(n_449), .B2(n_450), .C(n_451), .Y(n_447) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx4f_ASAP7_75t_L g565 ( .A(n_432), .Y(n_565) );
INVx2_ASAP7_75t_L g577 ( .A(n_432), .Y(n_577) );
INVx1_ASAP7_75t_L g653 ( .A(n_432), .Y(n_653) );
BUFx2_ASAP7_75t_L g742 ( .A(n_432), .Y(n_742) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g744 ( .A(n_435), .Y(n_744) );
INVx3_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g587 ( .A(n_437), .Y(n_587) );
INVx2_ASAP7_75t_SL g644 ( .A(n_437), .Y(n_644) );
INVx1_ASAP7_75t_L g778 ( .A(n_437), .Y(n_778) );
INVx1_ASAP7_75t_L g1387 ( .A(n_437), .Y(n_1387) );
INVx1_ASAP7_75t_L g898 ( .A(n_438), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_444), .B2(n_445), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_441), .A2(n_498), .B1(n_499), .B2(n_502), .C(n_503), .Y(n_497) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g510 ( .A(n_443), .B(n_472), .Y(n_510) );
INVx2_ASAP7_75t_SL g1463 ( .A(n_443), .Y(n_1463) );
INVx1_ASAP7_75t_L g640 ( .A(n_445), .Y(n_640) );
INVx1_ASAP7_75t_L g1156 ( .A(n_445), .Y(n_1156) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_446), .Y(n_657) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_446), .Y(n_737) );
AND2x6_ASAP7_75t_L g917 ( .A(n_446), .B(n_904), .Y(n_917) );
INVx1_ASAP7_75t_L g975 ( .A(n_446), .Y(n_975) );
OAI221xp5_ASAP7_75t_L g1105 ( .A1(n_449), .A2(n_590), .B1(n_1106), .B2(n_1107), .C(n_1108), .Y(n_1105) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g507 ( .A(n_453), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_453), .Y(n_637) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_453), .Y(n_753) );
INVx2_ASAP7_75t_SL g785 ( .A(n_453), .Y(n_785) );
AND2x4_ASAP7_75t_L g977 ( .A(n_453), .B(n_516), .Y(n_977) );
AND2x4_ASAP7_75t_L g1396 ( .A(n_453), .B(n_516), .Y(n_1396) );
OAI31xp33_ASAP7_75t_SL g735 ( .A1(n_454), .A2(n_736), .A3(n_746), .B(n_754), .Y(n_735) );
CKINVDCx8_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g466 ( .A(n_456), .Y(n_466) );
AND2x4_ASAP7_75t_L g614 ( .A(n_456), .B(n_615), .Y(n_614) );
OR2x6_ASAP7_75t_L g960 ( .A(n_456), .B(n_587), .Y(n_960) );
AND2x4_ASAP7_75t_L g980 ( .A(n_456), .B(n_615), .Y(n_980) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_456), .B(n_1387), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_456), .B(n_1077), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_554), .B1(n_555), .B2(n_626), .Y(n_459) );
INVx1_ASAP7_75t_SL g626 ( .A(n_460), .Y(n_626) );
XNOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_517), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B1(n_511), .B2(n_512), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g556 ( .A1(n_466), .A2(n_557), .B(n_595), .C(n_606), .Y(n_556) );
NAND5xp2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_485), .C(n_493), .D(n_497), .E(n_508), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g876 ( .A(n_471), .Y(n_876) );
BUFx6f_ASAP7_75t_L g1469 ( .A(n_471), .Y(n_1469) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_472), .A2(n_559), .B(n_563), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_472), .A2(n_487), .B1(n_650), .B2(n_651), .C(n_658), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_472), .A2(n_760), .B(n_763), .Y(n_759) );
OAI21xp33_ASAP7_75t_L g791 ( .A1(n_472), .A2(n_792), .B(n_794), .Y(n_791) );
AND2x2_ASAP7_75t_L g873 ( .A(n_472), .B(n_562), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_473), .A2(n_486), .B1(n_548), .B2(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g639 ( .A(n_478), .Y(n_639) );
INVx1_ASAP7_75t_L g748 ( .A(n_478), .Y(n_748) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_489), .B2(n_490), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_487), .A2(n_860), .B1(n_863), .B2(n_871), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_487), .A2(n_490), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_487), .A2(n_510), .B1(n_1137), .B2(n_1141), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_487), .A2(n_490), .B1(n_1450), .B2(n_1454), .Y(n_1470) );
INVx6_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_489), .A2(n_509), .B1(n_539), .B2(n_542), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_490), .A2(n_861), .B1(n_883), .B2(n_884), .C(n_886), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_490), .A2(n_1139), .B1(n_1146), .B2(n_1149), .C(n_1151), .Y(n_1145) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g581 ( .A(n_492), .Y(n_581) );
INVx1_ASAP7_75t_L g762 ( .A(n_492), .Y(n_762) );
INVx3_ASAP7_75t_L g1008 ( .A(n_496), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_498), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_524) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g970 ( .A(n_501), .Y(n_970) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_506), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_510), .A2(n_1003), .B1(n_1004), .B2(n_1005), .C(n_1006), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_510), .A2(n_1449), .B1(n_1460), .B2(n_1461), .C(n_1464), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_512), .A2(n_1000), .B1(n_1001), .B2(n_1019), .Y(n_999) );
AOI21xp33_ASAP7_75t_SL g1456 ( .A1(n_512), .A2(n_1457), .B(n_1458), .Y(n_1456) );
INVx5_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g889 ( .A(n_513), .Y(n_889) );
INVx2_ASAP7_75t_L g1159 ( .A(n_513), .Y(n_1159) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_529), .C(n_533), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g676 ( .A(n_521), .Y(n_676) );
BUFx2_ASAP7_75t_L g705 ( .A(n_521), .Y(n_705) );
BUFx2_ASAP7_75t_L g836 ( .A(n_521), .Y(n_836) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_521), .Y(n_1121) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_522), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_526), .A2(n_712), .B(n_713), .Y(n_711) );
BUFx2_ASAP7_75t_L g801 ( .A(n_526), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_526), .A2(n_672), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_526), .A2(n_528), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_526), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_526), .A2(n_1126), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_528), .A2(n_598), .B1(n_788), .B2(n_826), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g1445 ( .A1(n_536), .A2(n_549), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_541), .B1(n_542), .B2(n_545), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g816 ( .A(n_543), .Y(n_816) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g717 ( .A(n_544), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_544), .A2(n_776), .B1(n_810), .B2(n_813), .Y(n_809) );
INVx2_ASAP7_75t_L g1071 ( .A(n_544), .Y(n_1071) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI322xp5_ASAP7_75t_L g607 ( .A1(n_553), .A2(n_589), .A3(n_608), .B1(n_610), .B2(n_614), .C1(n_616), .C2(n_619), .Y(n_607) );
AOI33xp33_ASAP7_75t_L g978 ( .A1(n_553), .A2(n_979), .A3(n_981), .B1(n_985), .B2(n_992), .B3(n_993), .Y(n_978) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .C(n_574), .D(n_588), .Y(n_557) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g969 ( .A(n_562), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_564), .A2(n_751), .B1(n_782), .B2(n_783), .C(n_784), .Y(n_781) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g750 ( .A(n_565), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_569), .C(n_572), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_567), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_SL g787 ( .A1(n_568), .A2(n_572), .B(n_788), .C(n_789), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g755 ( .A1(n_572), .A2(n_594), .B(n_643), .C(n_710), .Y(n_755) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI211xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_578), .C(n_582), .Y(n_574) );
BUFx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g591 ( .A(n_577), .Y(n_591) );
INVx1_ASAP7_75t_L g739 ( .A(n_579), .Y(n_739) );
BUFx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g1114 ( .A(n_581), .Y(n_1114) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_592), .C(n_593), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_598), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_598), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_600), .A2(n_621), .B1(n_624), .B2(n_668), .C(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g766 ( .A(n_600), .Y(n_766) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_620), .Y(n_606) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g721 ( .A(n_612), .Y(n_721) );
BUFx2_ASAP7_75t_L g982 ( .A(n_612), .Y(n_982) );
BUFx6f_ASAP7_75t_L g1407 ( .A(n_613), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g768 ( .A(n_621), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_624), .A2(n_757), .B1(n_758), .B2(n_765), .C(n_767), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_624), .A2(n_765), .B1(n_767), .B2(n_798), .C(n_799), .Y(n_827) );
INVx1_ASAP7_75t_L g935 ( .A(n_625), .Y(n_935) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_666), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_649), .B(n_663), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_638), .B1(n_641), .B2(n_645), .C(n_648), .Y(n_632) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g745 ( .A(n_644), .Y(n_745) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx4_ASAP7_75t_L g797 ( .A(n_660), .Y(n_797) );
INVx2_ASAP7_75t_L g887 ( .A(n_660), .Y(n_887) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_662), .A2(n_796), .B1(n_798), .B2(n_799), .Y(n_795) );
INVx2_ASAP7_75t_SL g1465 ( .A(n_662), .Y(n_1465) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI31xp33_ASAP7_75t_SL g771 ( .A1(n_664), .A2(n_772), .A3(n_779), .B(n_786), .Y(n_771) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g868 ( .A(n_665), .Y(n_868) );
AND2x4_ASAP7_75t_L g897 ( .A(n_665), .B(n_898), .Y(n_897) );
AND2x4_ASAP7_75t_L g1382 ( .A(n_665), .B(n_898), .Y(n_1382) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .C(n_674), .D(n_678), .Y(n_666) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_684), .Y(n_1138) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_892), .B1(n_1161), .B2(n_1162), .Y(n_696) );
INVx1_ASAP7_75t_L g1162 ( .A(n_697), .Y(n_1162) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_828), .B1(n_890), .B2(n_891), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_699), .Y(n_890) );
XOR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_769), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_702), .B(n_711), .C(n_735), .D(n_764), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_706), .A2(n_712), .B1(n_750), .B2(n_751), .C(n_753), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g740 ( .A1(n_715), .A2(n_741), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_740) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g1075 ( .A(n_721), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_721), .Y(n_1403) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .C(n_730), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_726), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_814) );
OAI22xp5_ASAP7_75t_SL g1035 ( .A1(n_728), .A2(n_1036), .B1(n_1037), .B2(n_1039), .Y(n_1035) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_732), .B(n_1091), .Y(n_1090) );
OAI33xp33_ASAP7_75t_L g843 ( .A1(n_733), .A2(n_844), .A3(n_845), .B1(n_852), .B2(n_857), .B3(n_862), .Y(n_843) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_733), .A2(n_844), .A3(n_1129), .B1(n_1132), .B2(n_1136), .B3(n_1140), .Y(n_1128) );
CKINVDCx8_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g774 ( .A(n_742), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_744), .A2(n_774), .B1(n_775), .B2(n_776), .C(n_777), .Y(n_773) );
INVx1_ASAP7_75t_L g1150 ( .A(n_744), .Y(n_1150) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .C(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_800), .C(n_822), .D(n_827), .Y(n_770) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_783), .A2(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND3xp33_ASAP7_75t_SL g786 ( .A(n_787), .B(n_791), .C(n_795), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g1011 ( .A(n_790), .Y(n_1011) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g1073 ( .A(n_806), .Y(n_1073) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OR2x6_ASAP7_75t_L g1067 ( .A(n_807), .B(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g850 ( .A(n_808), .Y(n_850) );
INVx2_ASAP7_75t_L g1034 ( .A(n_808), .Y(n_1034) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_808), .Y(n_1045) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g854 ( .A(n_812), .Y(n_854) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g891 ( .A(n_828), .Y(n_891) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
XNOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_865), .Y(n_831) );
NOR3xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_841), .C(n_843), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_838), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_848), .B1(n_849), .B2(n_851), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_846), .A2(n_849), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_846), .A2(n_849), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_849), .A2(n_1452), .B1(n_1454), .B2(n_1455), .Y(n_1451) );
BUFx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_853), .A2(n_1133), .B1(n_1134), .B2(n_1135), .Y(n_1132) );
BUFx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
BUFx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g1038 ( .A(n_859), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_869), .B1(n_888), .B2(n_889), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_866), .A2(n_1144), .B1(n_1158), .B2(n_1159), .Y(n_1143) );
INVx5_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
AOI221x1_ASAP7_75t_SL g1051 ( .A1(n_867), .A2(n_897), .B1(n_1052), .B2(n_1064), .C(n_1102), .Y(n_1051) );
AOI31xp33_ASAP7_75t_L g1458 ( .A1(n_867), .A2(n_1459), .A3(n_1466), .B(n_1470), .Y(n_1458) );
BUFx8_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g1000 ( .A(n_868), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_874), .C(n_882), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1161 ( .A(n_892), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_1048), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_996), .B2(n_1047), .Y(n_893) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g995 ( .A(n_896), .Y(n_995) );
AO211x2_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_899), .B(n_931), .C(n_957), .Y(n_896) );
NAND4xp25_ASAP7_75t_L g899 ( .A(n_900), .B(n_911), .C(n_918), .D(n_928), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_902), .B1(n_907), .B2(n_908), .Y(n_900) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_903), .A2(n_908), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_903), .A2(n_908), .B1(n_1372), .B2(n_1373), .Y(n_1371) );
AND2x4_ASAP7_75t_L g903 ( .A(n_904), .B(n_906), .Y(n_903) );
INVx1_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g930 ( .A(n_909), .Y(n_930) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B1(n_916), .B2(n_917), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_912), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_913), .A2(n_917), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_913), .A2(n_917), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
AND2x4_ASAP7_75t_L g923 ( .A(n_914), .B(n_924), .Y(n_923) );
AND2x2_ASAP7_75t_SL g1377 ( .A(n_914), .B(n_924), .Y(n_1377) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AOI222xp33_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_920), .B1(n_921), .B2(n_922), .C1(n_926), .C2(n_927), .Y(n_918) );
AOI222xp33_ASAP7_75t_L g1057 ( .A1(n_922), .A2(n_927), .B1(n_964), .B2(n_1058), .C1(n_1059), .C2(n_1060), .Y(n_1057) );
BUFx4f_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AOI222xp33_ASAP7_75t_L g1374 ( .A1(n_927), .A2(n_1147), .B1(n_1375), .B2(n_1376), .C1(n_1377), .C2(n_1378), .Y(n_1374) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_928), .Y(n_1053) );
INVx5_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
CKINVDCx8_ASAP7_75t_R g1370 ( .A(n_929), .Y(n_1370) );
AOI31xp33_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_943), .A3(n_951), .B(n_956), .Y(n_931) );
AOI211xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B(n_936), .C(n_939), .Y(n_932) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI211xp5_ASAP7_75t_L g1405 ( .A1(n_936), .A2(n_1406), .B(n_1407), .C(n_1408), .Y(n_1405) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g1409 ( .A(n_941), .Y(n_1409) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_944), .A2(n_946), .B1(n_947), .B2(n_950), .Y(n_943) );
AOI22xp33_ASAP7_75t_SL g1411 ( .A1(n_944), .A2(n_947), .B1(n_1412), .B2(n_1413), .Y(n_1411) );
AND2x4_ASAP7_75t_L g947 ( .A(n_945), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_949), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g1414 ( .A1(n_952), .A2(n_1380), .B1(n_1415), .B2(n_1416), .Y(n_1414) );
INVx4_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx5_ASAP7_75t_L g1416 ( .A(n_955), .Y(n_1416) );
AOI31xp33_ASAP7_75t_L g1404 ( .A1(n_956), .A2(n_1405), .A3(n_1411), .B(n_1414), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_978), .Y(n_957) );
AOI33xp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_961), .A3(n_968), .B1(n_971), .B2(n_973), .B3(n_976), .Y(n_958) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_960), .Y(n_959) );
INVx2_ASAP7_75t_L g1104 ( .A(n_960), .Y(n_1104) );
BUFx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx2_ASAP7_75t_L g1399 ( .A(n_967), .Y(n_1399) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
BUFx4f_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx4_ASAP7_75t_L g1110 ( .A(n_977), .Y(n_1110) );
BUFx3_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AOI33xp33_ASAP7_75t_L g1395 ( .A1(n_980), .A2(n_1396), .A3(n_1397), .B1(n_1400), .B2(n_1401), .B3(n_1402), .Y(n_1395) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
BUFx3_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx2_ASAP7_75t_SL g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1047 ( .A(n_997), .Y(n_1047) );
XOR2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1046), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1020), .Y(n_998) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1009), .C(n_1016), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_1005), .A2(n_1018), .B1(n_1037), .B2(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1014), .Y(n_1390) );
INVx2_ASAP7_75t_SL g1398 ( .A(n_1014), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_1015), .A2(n_1017), .B1(n_1032), .B2(n_1044), .Y(n_1043) );
NOR3xp33_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1028), .C(n_1029), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B1(n_1033), .B2(n_1034), .Y(n_1030) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1443 ( .A(n_1038), .Y(n_1443) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_1042), .Y(n_1041) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AO22x2_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1050), .B1(n_1115), .B2(n_1160), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND4xp25_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .C(n_1057), .D(n_1061), .Y(n_1052) );
AOI222xp33_ASAP7_75t_L g1085 ( .A1(n_1055), .A2(n_1086), .B1(n_1089), .B2(n_1090), .C1(n_1093), .C2(n_1094), .Y(n_1085) );
OAI21xp5_ASAP7_75t_SL g1072 ( .A1(n_1058), .A2(n_1073), .B(n_1074), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1085), .C(n_1095), .Y(n_1064) );
NOR3xp33_ASAP7_75t_SL g1065 ( .A(n_1066), .B(n_1070), .C(n_1078), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1068), .Y(n_1080) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1068), .Y(n_1088) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_1077), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1091), .B(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_1096), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1095) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_1103), .A2(n_1105), .B1(n_1110), .B2(n_1111), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1115), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1143), .Y(n_1116) );
NOR3xp33_ASAP7_75t_SL g1117 ( .A(n_1118), .B(n_1127), .C(n_1128), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1123), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1152), .C(n_1157), .Y(n_1144) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1364), .B1(n_1366), .B2(n_1418), .C(n_1423), .Y(n_1163) );
NOR3xp33_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1304), .C(n_1342), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1240), .B1(n_1285), .B2(n_1293), .Y(n_1165) );
NOR3xp33_ASAP7_75t_SL g1166 ( .A(n_1167), .B(n_1250), .C(n_1253), .Y(n_1166) );
A2O1A1Ixp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1203), .B(n_1211), .C(n_1225), .Y(n_1167) );
O2A1O1Ixp33_ASAP7_75t_L g1360 ( .A1(n_1168), .A2(n_1170), .B(n_1361), .C(n_1362), .Y(n_1360) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1169), .B(n_1207), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1190), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1170), .B(n_1230), .Y(n_1296) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1170), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1170), .B(n_1259), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1170), .B(n_1263), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1170), .B(n_1217), .Y(n_1357) );
INVx4_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1171), .B(n_1214), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1171), .B(n_1205), .Y(n_1252) );
INVx3_ASAP7_75t_L g1261 ( .A(n_1171), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1171), .B(n_1257), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1171), .B(n_1190), .Y(n_1278) );
NOR2xp67_ASAP7_75t_SL g1280 ( .A(n_1171), .B(n_1239), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1171), .B(n_1207), .Y(n_1311) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_1171), .B(n_1329), .C(n_1338), .Y(n_1340) );
AOI211xp5_ASAP7_75t_L g1344 ( .A1(n_1171), .A2(n_1272), .B(n_1345), .C(n_1346), .Y(n_1344) );
AND2x4_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1184), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1179), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1175), .B(n_1180), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1178), .Y(n_1187) );
AND2x4_ASAP7_75t_L g1181 ( .A(n_1179), .B(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1180), .B(n_1183), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1472 ( .A(n_1182), .Y(n_1472) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1185), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1188), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1186), .B(n_1188), .Y(n_1236) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1187), .B(n_1188), .Y(n_1189) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1189), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1190), .B(n_1208), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1190), .B(n_1296), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1190), .B(n_1311), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1199), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1191), .B(n_1206), .Y(n_1257) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1192), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1192), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1192), .B(n_1199), .Y(n_1284) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1195), .B1(n_1197), .B2(n_1198), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_1195), .A2(n_1198), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_1195), .A2(n_1222), .B1(n_1223), .B2(n_1224), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1246 ( .A(n_1195), .Y(n_1246) );
BUFx6f_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1224 ( .A(n_1198), .Y(n_1224) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1198), .Y(n_1249) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1199), .Y(n_1206) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1203), .B(n_1270), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1207), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1205), .B(n_1296), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1205), .B(n_1311), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1206), .B(n_1230), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1206), .B(n_1207), .Y(n_1239) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1206), .Y(n_1341) );
OAI322xp33_ASAP7_75t_L g1355 ( .A1(n_1206), .A2(n_1232), .A3(n_1239), .B1(n_1263), .B2(n_1356), .C1(n_1358), .C2(n_1359), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1207), .B(n_1252), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1207), .B(n_1264), .Y(n_1273) );
BUFx3_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1208), .Y(n_1230) );
AOI222xp33_ASAP7_75t_L g1279 ( .A1(n_1208), .A2(n_1234), .B1(n_1259), .B2(n_1280), .C1(n_1281), .C2(n_1283), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1208), .B(n_1257), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1208), .B(n_1284), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1217), .Y(n_1211) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_1212), .A2(n_1255), .B1(n_1258), .B2(n_1260), .Y(n_1254) );
A2O1A1Ixp33_ASAP7_75t_L g1293 ( .A1(n_1212), .A2(n_1294), .B(n_1297), .C(n_1303), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1212), .B(n_1218), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1212), .B(n_1350), .Y(n_1349) );
INVx3_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_1213), .B(n_1251), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1213), .B(n_1233), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1213), .B(n_1271), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1213), .B(n_1292), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_1214), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1214), .B(n_1234), .Y(n_1259) );
INVx1_ASAP7_75t_SL g1277 ( .A(n_1214), .Y(n_1277) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1214), .Y(n_1317) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1214), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1214), .B(n_1233), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1217), .B(n_1233), .Y(n_1232) );
AND2x4_ASAP7_75t_SL g1271 ( .A(n_1217), .B(n_1233), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1217), .B(n_1234), .Y(n_1322) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1218), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1218), .B(n_1233), .Y(n_1303) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1229), .B1(n_1231), .B2(n_1238), .C(n_1240), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1228), .Y(n_1226) );
OAI211xp5_ASAP7_75t_SL g1253 ( .A1(n_1227), .A2(n_1254), .B(n_1265), .C(n_1279), .Y(n_1253) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1227), .Y(n_1282) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1227), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1227), .B(n_1241), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1227), .B(n_1259), .Y(n_1346) );
O2A1O1Ixp33_ASAP7_75t_L g1347 ( .A1(n_1227), .A2(n_1348), .B(n_1351), .C(n_1352), .Y(n_1347) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1228), .Y(n_1326) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1229), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1230), .B(n_1257), .Y(n_1256) );
NOR2x1_ASAP7_75t_L g1263 ( .A(n_1230), .B(n_1264), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1230), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1233), .B(n_1298), .Y(n_1337) );
CKINVDCx6p67_ASAP7_75t_R g1233 ( .A(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1234), .B(n_1277), .Y(n_1276) );
OR2x6_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1237), .Y(n_1234) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
OAI31xp33_ASAP7_75t_L g1305 ( .A1(n_1241), .A2(n_1306), .A3(n_1315), .B(n_1327), .Y(n_1305) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_1245), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g1365 ( .A(n_1248), .Y(n_1365) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1251), .Y(n_1351) );
OAI31xp33_ASAP7_75t_SL g1313 ( .A1(n_1255), .A2(n_1308), .A3(n_1310), .B(n_1314), .Y(n_1313) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1255), .A2(n_1321), .B(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1257), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_1258), .A2(n_1261), .B1(n_1287), .B2(n_1289), .Y(n_1286) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1259), .B(n_1357), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1262), .Y(n_1260) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1261), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_1261), .A2(n_1298), .B1(n_1299), .B2(n_1301), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1261), .B(n_1300), .Y(n_1331) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1264), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1268), .B1(n_1269), .B2(n_1272), .C(n_1274), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1268), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1268), .Y(n_1312) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1271), .Y(n_1343) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1276), .B(n_1282), .Y(n_1281) );
OAI21xp5_ASAP7_75t_SL g1353 ( .A1(n_1276), .A2(n_1300), .B(n_1321), .Y(n_1353) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1280), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1281), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1283), .B(n_1288), .Y(n_1292) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1284), .Y(n_1336) );
AOI21xp33_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1290), .B(n_1291), .Y(n_1285) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OAI21xp33_ASAP7_75t_L g1323 ( .A1(n_1302), .A2(n_1324), .B(n_1326), .Y(n_1323) );
NAND2xp5_ASAP7_75t_SL g1304 ( .A(n_1305), .B(n_1332), .Y(n_1304) );
A2O1A1Ixp33_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1309), .B(n_1312), .C(n_1313), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
A2O1A1Ixp33_ASAP7_75t_L g1352 ( .A1(n_1312), .A2(n_1318), .B(n_1350), .C(n_1353), .Y(n_1352) );
OAI211xp5_ASAP7_75t_SL g1315 ( .A1(n_1316), .A2(n_1318), .B(n_1320), .C(n_1323), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1322), .B(n_1325), .Y(n_1324) );
AOI21xp33_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1330), .B(n_1331), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AOI32xp33_ASAP7_75t_L g1332 ( .A1(n_1333), .A2(n_1337), .A3(n_1338), .B1(n_1339), .B2(n_1341), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1336), .Y(n_1334) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
OAI211xp5_ASAP7_75t_SL g1342 ( .A1(n_1343), .A2(n_1344), .B(n_1347), .C(n_1354), .Y(n_1342) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1346), .Y(n_1362) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NOR3xp33_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1360), .C(n_1363), .Y(n_1354) );
BUFx2_ASAP7_75t_SL g1364 ( .A(n_1365), .Y(n_1364) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1368), .Y(n_1417) );
AOI211x1_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1382), .B(n_1383), .C(n_1404), .Y(n_1368) );
NAND4xp25_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1371), .C(n_1374), .D(n_1379), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1395), .Y(n_1383) );
AOI33xp33_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1388), .A3(n_1389), .B1(n_1392), .B2(n_1393), .B3(n_1394), .Y(n_1384) );
INVx3_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
CKINVDCx14_ASAP7_75t_R g1418 ( .A(n_1419), .Y(n_1418) );
BUFx2_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_1426), .Y(n_1425) );
OAI21xp5_ASAP7_75t_L g1471 ( .A1(n_1427), .A2(n_1472), .B(n_1473), .Y(n_1471) );
INVxp33_ASAP7_75t_SL g1428 ( .A(n_1429), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1456), .Y(n_1430) );
NOR3xp33_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1439), .C(n_1440), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1436), .Y(n_1432) );
INVx3_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
endmodule