module fake_jpeg_24013_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_45)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_21),
.B1(n_14),
.B2(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_61),
.B1(n_69),
.B2(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_43),
.C(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_34),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_66),
.B1(n_38),
.B2(n_20),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_63),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_17),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_35),
.B1(n_29),
.B2(n_28),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_83),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_35),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_60),
.B(n_23),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.B1(n_65),
.B2(n_53),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_18),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_61),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_93),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_50),
.C(n_67),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_97),
.C(n_80),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_98),
.B(n_72),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_32),
.B1(n_22),
.B2(n_14),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_15),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_19),
.B1(n_23),
.B2(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_82),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_83),
.B(n_71),
.C(n_77),
.D(n_79),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_106),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_80),
.C(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_93),
.B1(n_88),
.B2(n_94),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_98),
.B1(n_81),
.B2(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_114),
.C(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_91),
.A3(n_84),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_100),
.B(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_113),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_104),
.Y(n_120)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_115),
.B(n_113),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_2),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_4),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_123),
.B(n_120),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_132),
.A3(n_128),
.B1(n_126),
.B2(n_125),
.C1(n_127),
.C2(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_133),
.B(n_132),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_5),
.Y(n_137)
);


endmodule