module fake_netlist_1_10933_n_500 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_139, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_145, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_500);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_139;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_145;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_500;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_479;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_486;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_283;
wire n_435;
wire n_216;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_25), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_41), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_139), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_26), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_39), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_29), .Y(n_160) );
INVxp33_ASAP7_75t_SL g161 ( .A(n_93), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_98), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_95), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_118), .Y(n_164) );
CKINVDCx14_ASAP7_75t_R g165 ( .A(n_124), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_60), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_67), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_134), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_3), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_107), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_49), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_138), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_103), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_54), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_113), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_81), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_90), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_116), .Y(n_182) );
BUFx2_ASAP7_75t_SL g183 ( .A(n_85), .Y(n_183) );
INVx1_ASAP7_75t_SL g184 ( .A(n_78), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_100), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_61), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_108), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_92), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_71), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_106), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_16), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_10), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_126), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_31), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_36), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_135), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_59), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_130), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_35), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_127), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_110), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_75), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_122), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_19), .Y(n_206) );
NOR2xp67_ASAP7_75t_L g207 ( .A(n_147), .B(n_87), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_68), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_73), .Y(n_209) );
BUFx5_ASAP7_75t_L g210 ( .A(n_76), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_24), .Y(n_211) );
INVxp67_ASAP7_75t_SL g212 ( .A(n_50), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_45), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_88), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_3), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_82), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_77), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_125), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_105), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_4), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_0), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_109), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_46), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_2), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_9), .Y(n_228) );
BUFx2_ASAP7_75t_SL g229 ( .A(n_117), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_65), .Y(n_230) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_33), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_84), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_91), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_151), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_28), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_15), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_169), .B(n_0), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_232), .B(n_1), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_223), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_196), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_191), .B(n_5), .Y(n_244) );
CKINVDCx8_ASAP7_75t_R g245 ( .A(n_183), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_157), .B(n_5), .Y(n_246) );
BUFx8_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_170), .A2(n_80), .B(n_143), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_194), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_210), .B(n_6), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_173), .B(n_6), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_234), .B(n_7), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_224), .B(n_8), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_179), .B(n_9), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_181), .B(n_10), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_193), .B(n_11), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_228), .Y(n_259) );
BUFx4f_ASAP7_75t_L g260 ( .A(n_259), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_238), .A2(n_161), .B1(n_236), .B2(n_227), .Y(n_261) );
INVx5_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_257), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_240), .Y(n_264) );
AND2x6_ASAP7_75t_L g265 ( .A(n_244), .B(n_152), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_241), .B(n_220), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_247), .B(n_153), .Y(n_267) );
INVx5_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_247), .B(n_197), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_237), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_249), .B(n_154), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_245), .Y(n_272) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_238), .B(n_160), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_242), .Y(n_274) );
AND2x6_ASAP7_75t_L g275 ( .A(n_252), .B(n_156), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_237), .Y(n_276) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_253), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_231), .B1(n_165), .B2(n_229), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_277), .B(n_255), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_270), .B(n_251), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_277), .B(n_258), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_276), .A2(n_256), .B(n_250), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_272), .B(n_239), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_279), .B(n_158), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_260), .B(n_248), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_272), .B(n_11), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_263), .B(n_164), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_269), .B(n_166), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_261), .A2(n_162), .B1(n_172), .B2(n_155), .Y(n_292) );
NAND2x1p5_ASAP7_75t_L g293 ( .A(n_263), .B(n_184), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_278), .B(n_159), .Y(n_294) );
NAND2x1_ASAP7_75t_L g295 ( .A(n_265), .B(n_163), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_265), .B(n_168), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_291), .B(n_267), .Y(n_298) );
OAI22x1_ASAP7_75t_L g299 ( .A1(n_284), .A2(n_212), .B1(n_275), .B2(n_265), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_292), .B(n_273), .C(n_266), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_281), .B(n_275), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_205), .B1(n_189), .B2(n_200), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_286), .A2(n_171), .B(n_167), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_293), .B(n_176), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_280), .A2(n_175), .B(n_174), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_203), .B(n_235), .C(n_230), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_283), .A2(n_178), .B(n_177), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_297), .A2(n_182), .B(n_180), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_294), .A2(n_186), .B(n_185), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_305), .A2(n_296), .B(n_187), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_307), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_302), .A2(n_290), .B(n_289), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_301), .B(n_287), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_311), .A2(n_296), .B(n_188), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_303), .A2(n_213), .B1(n_190), .B2(n_192), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_312), .A2(n_199), .B(n_198), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_300), .A2(n_218), .B1(n_202), .B2(n_204), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_308), .A2(n_208), .B(n_201), .Y(n_324) );
BUFx12f_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_298), .B(n_207), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_309), .A2(n_217), .B(n_226), .C(n_225), .Y(n_328) );
AO21x1_ASAP7_75t_L g329 ( .A1(n_313), .A2(n_215), .B(n_214), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_306), .A2(n_222), .B1(n_219), .B2(n_209), .C(n_211), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_303), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_304), .A2(n_12), .B(n_13), .C(n_14), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_323), .A2(n_210), .B(n_243), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
OA21x2_ASAP7_75t_L g335 ( .A1(n_319), .A2(n_233), .B(n_221), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
AO31x2_ASAP7_75t_L g337 ( .A1(n_329), .A2(n_254), .A3(n_206), .B(n_13), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_314), .A2(n_206), .B(n_17), .Y(n_338) );
AO31x2_ASAP7_75t_L g339 ( .A1(n_321), .A2(n_14), .A3(n_18), .B(n_20), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_332), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_318), .B(n_21), .Y(n_342) );
INVx6_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_327), .B(n_22), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_328), .A2(n_268), .B(n_262), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_320), .B(n_23), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_326), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_330), .Y(n_350) );
BUFx8_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_331), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_317), .B(n_27), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_315), .B(n_268), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_316), .A2(n_30), .B(n_32), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_317), .B(n_145), .Y(n_357) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_319), .A2(n_34), .B(n_37), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_315), .B(n_38), .Y(n_359) );
BUFx10_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_40), .B(n_42), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_351), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_354), .B(n_43), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_353), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_353), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_354), .B(n_44), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_338), .A2(n_349), .B(n_345), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_360), .Y(n_370) );
AOI21x1_ASAP7_75t_L g371 ( .A1(n_358), .A2(n_47), .B(n_48), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_342), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_356), .A2(n_51), .B(n_52), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_340), .A2(n_53), .B(n_55), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_350), .B(n_56), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_350), .B(n_57), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_341), .B(n_142), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_357), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_349), .B(n_58), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_341), .B(n_352), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_344), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
BUFx4f_ASAP7_75t_L g385 ( .A(n_341), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_348), .B(n_141), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_359), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_333), .A2(n_62), .B(n_63), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_64), .B(n_66), .Y(n_390) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_346), .A2(n_69), .B(n_70), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_343), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_347), .A2(n_72), .B(n_74), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_335), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_334), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_334), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_334), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_334), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_334), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_334), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_364), .B(n_79), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_362), .B(n_86), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_398), .B(n_89), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_399), .B(n_94), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_401), .B(n_96), .Y(n_409) );
BUFx6f_ASAP7_75t_SL g410 ( .A(n_363), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_364), .B(n_97), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_402), .B(n_99), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_402), .B(n_101), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_364), .B(n_102), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_367), .B(n_104), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_400), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_403), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_111), .B1(n_112), .B2(n_114), .C(n_115), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_397), .B(n_140), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_119), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_383), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_372), .A2(n_120), .B(n_121), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_382), .B(n_123), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_373), .B(n_131), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_379), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_374), .A2(n_378), .B1(n_377), .B2(n_388), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
INVx2_ASAP7_75t_R g440 ( .A(n_436), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_410), .B(n_387), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_419), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_404), .A2(n_395), .B1(n_381), .B2(n_376), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_421), .B(n_393), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_418), .B(n_391), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_417), .B(n_393), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_437), .B(n_390), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_428), .B(n_389), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_423), .B(n_371), .C(n_375), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_439), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_429), .B(n_433), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_404), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_435), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_438), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_441), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_457), .B(n_430), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_454), .B(n_432), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_456), .A2(n_414), .B1(n_411), .B2(n_415), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_456), .B(n_431), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_454), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_449), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_443), .B(n_413), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_444), .B(n_413), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_450), .B(n_446), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_440), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_465), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_461), .B(n_459), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_460), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_469), .B(n_448), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_465), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_464), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_466), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_464), .B(n_452), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_463), .B(n_445), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_470), .B(n_458), .Y(n_480) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_479), .A2(n_442), .B(n_455), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_477), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_472), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_473), .Y(n_484) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_476), .A2(n_480), .B(n_478), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_482), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_481), .B(n_471), .C(n_475), .Y(n_487) );
OAI21xp33_ASAP7_75t_SL g488 ( .A1(n_485), .A2(n_477), .B(n_474), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_483), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_484), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_488), .A2(n_490), .B1(n_486), .B2(n_487), .C(n_489), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_491), .B(n_422), .C(n_453), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_492), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_493), .A2(n_447), .B1(n_434), .B2(n_451), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_494), .A2(n_468), .B1(n_467), .B2(n_462), .Y(n_495) );
OAI21x1_ASAP7_75t_SL g496 ( .A1(n_495), .A2(n_427), .B(n_468), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_496), .A2(n_408), .B1(n_412), .B2(n_409), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_497), .Y(n_498) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_498), .A2(n_427), .B(n_425), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_499), .A2(n_406), .B(n_407), .Y(n_500) );
endmodule