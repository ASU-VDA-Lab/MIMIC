module fake_jpeg_26790_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_54),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_70),
.B1(n_22),
.B2(n_31),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_71),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_25),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_72),
.B(n_17),
.C(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_68),
.B1(n_22),
.B2(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_24),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_0),
.Y(n_72)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_86),
.B1(n_53),
.B2(n_62),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_25),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_83),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_42),
.C(n_37),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_98),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_82),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_57),
.A3(n_55),
.B1(n_48),
.B2(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_106),
.B1(n_58),
.B2(n_19),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_45),
.B1(n_26),
.B2(n_30),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_95),
.B1(n_99),
.B2(n_53),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_50),
.B1(n_61),
.B2(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_21),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_105),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_17),
.Y(n_98)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_17),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_23),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_0),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_131),
.B1(n_94),
.B2(n_74),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_65),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_123),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_88),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_58),
.B1(n_20),
.B2(n_19),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_125),
.B1(n_132),
.B2(n_66),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_75),
.B1(n_98),
.B2(n_89),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_93),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

OAI22x1_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_29),
.B1(n_37),
.B2(n_64),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_37),
.C(n_29),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_106),
.C(n_73),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_73),
.B1(n_83),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_64),
.B1(n_49),
.B2(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_140),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_145),
.B(n_147),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_102),
.B1(n_92),
.B2(n_80),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_120),
.B1(n_126),
.B2(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_49),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_153),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_1),
.C(n_2),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_1),
.C(n_4),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_114),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_128),
.C(n_131),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_157),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_66),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_110),
.B(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_108),
.B(n_66),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_117),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_163),
.B1(n_174),
.B2(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_107),
.B1(n_125),
.B2(n_133),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_143),
.C(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_181),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_133),
.B(n_108),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_169),
.B(n_156),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_116),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_120),
.B1(n_118),
.B2(n_126),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_132),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_152),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_135),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_192),
.C(n_172),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_135),
.B(n_138),
.C(n_158),
.D(n_147),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_194),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_136),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_191),
.B1(n_195),
.B2(n_198),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_193),
.C(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_167),
.B(n_177),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_140),
.C(n_149),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_157),
.A3(n_156),
.B1(n_137),
.B2(n_159),
.C1(n_112),
.C2(n_141),
.Y(n_193)
);

OA21x2_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_1),
.B(n_4),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_141),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_168),
.B1(n_171),
.B2(n_175),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_16),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_160),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_205),
.C(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_199),
.B1(n_196),
.B2(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_170),
.C(n_178),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_180),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_209),
.B(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_208),
.B1(n_183),
.B2(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_163),
.B1(n_167),
.B2(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_178),
.B1(n_160),
.B2(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_185),
.B1(n_197),
.B2(n_8),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_7),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_5),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_219),
.B1(n_221),
.B2(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_225),
.B(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_216),
.B(n_220),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_8),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_11),
.B(n_12),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_213),
.C(n_205),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_10),
.B(n_11),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_206),
.B(n_201),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_234),
.B(n_222),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_232),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_202),
.B1(n_210),
.B2(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_231),
.B1(n_12),
.B2(n_14),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_224),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_204),
.B(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_239),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_238),
.Y(n_244)
);

OAI221xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_219),
.B1(n_218),
.B2(n_221),
.C(n_14),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_227),
.C(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_14),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_240),
.A2(n_227),
.B(n_230),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_245),
.B(n_15),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_12),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_15),
.B(n_244),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_248),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_242),
.B(n_15),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);


endmodule