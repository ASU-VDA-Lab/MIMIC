module fake_jpeg_28156_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_57),
.B1(n_36),
.B2(n_45),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_18),
.B(n_16),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_43),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_68),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_22),
.B1(n_16),
.B2(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_45),
.B1(n_39),
.B2(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_40),
.B1(n_42),
.B2(n_38),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_82),
.B1(n_95),
.B2(n_51),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_45),
.B1(n_42),
.B2(n_28),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_17),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_78),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_83),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_94),
.Y(n_104)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_23),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_91),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_51),
.B1(n_58),
.B2(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_41),
.B1(n_38),
.B2(n_46),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_108),
.B1(n_55),
.B2(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_112),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_117),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_66),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_94),
.B1(n_90),
.B2(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_58),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_110),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_122),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_126),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_84),
.C(n_93),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_92),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_115),
.B1(n_116),
.B2(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_108),
.B1(n_115),
.B2(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_98),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_46),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_102),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_133),
.B1(n_121),
.B2(n_132),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_116),
.B(n_104),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_150),
.B1(n_142),
.B2(n_155),
.C(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_152),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_102),
.B(n_101),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_114),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_114),
.B(n_94),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_147),
.C(n_152),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_157),
.C(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_121),
.C(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_163),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_162),
.B1(n_153),
.B2(n_140),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_137),
.C(n_125),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_124),
.B1(n_135),
.B2(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_75),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_168),
.B(n_161),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_171),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_153),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_175),
.B1(n_166),
.B2(n_4),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_140),
.C(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_8),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_166),
.B1(n_9),
.B2(n_6),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_15),
.B(n_8),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_174),
.B1(n_171),
.B2(n_178),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_176),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_189),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_9),
.B(n_12),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_183),
.C(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_192),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_184),
.B1(n_5),
.B2(n_50),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_5),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_193),
.C(n_50),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_197),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_196),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);


endmodule