module fake_netlist_1_10171_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_0), .B(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_2), .B(n_7), .Y(n_16) );
A2O1A1Ixp33_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_1), .B(n_3), .C(n_4), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_13), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_16), .B(n_14), .Y(n_20) );
OA21x2_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_12), .B(n_19), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_21), .Y(n_25) );
XOR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_1), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_23), .Y(n_27) );
OAI21xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_25), .B(n_23), .Y(n_28) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_26), .B(n_3), .Y(n_29) );
INVx3_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_11), .Y(n_32) );
NAND4xp25_ASAP7_75t_L g33 ( .A(n_29), .B(n_11), .C(n_19), .D(n_9), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_28), .B1(n_19), .B2(n_10), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_35), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .B1(n_31), .B2(n_8), .Y(n_37) );
endmodule