module fake_jpeg_21229_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_2),
.B(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_54),
.C(n_47),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_4),
.C(n_5),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_52),
.B(n_44),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_15),
.B(n_27),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_45),
.B1(n_60),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_79),
.B1(n_78),
.B2(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_45),
.B1(n_54),
.B2(n_49),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_57),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_67),
.B1(n_60),
.B2(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_89),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_51),
.B(n_50),
.C(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_92),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_9),
.B(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_20),
.B1(n_32),
.B2(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_6),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_102),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_98),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.C(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_95),
.B1(n_104),
.B2(n_99),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_97),
.C(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_112),
.C(n_111),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_100),
.B1(n_109),
.B2(n_115),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_117),
.B1(n_109),
.B2(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_14),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_21),
.B(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_24),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_41),
.Y(n_125)
);


endmodule