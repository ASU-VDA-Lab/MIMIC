module fake_jpeg_3504_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_0),
.CON(n_75),
.SN(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_66),
.B1(n_60),
.B2(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_72),
.B1(n_77),
.B2(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_60),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_67),
.B1(n_54),
.B2(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_98),
.B1(n_102),
.B2(n_58),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_54),
.B1(n_63),
.B2(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_72),
.B1(n_55),
.B2(n_47),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_73),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_73),
.B1(n_58),
.B2(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_53),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_57),
.B1(n_53),
.B2(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_62),
.B1(n_56),
.B2(n_65),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_112),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_98),
.B(n_95),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_22),
.B(n_45),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_126),
.B(n_1),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_118),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_68),
.C(n_64),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_128),
.B1(n_119),
.B2(n_31),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_28),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_29),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_91),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_23),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_3),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_151),
.B(n_33),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_113),
.C(n_116),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_144),
.C(n_37),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_145),
.B(n_9),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_122),
.C(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_4),
.B(n_5),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_149),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_34),
.B(n_42),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_11),
.B(n_12),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_140),
.B(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_46),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.C(n_144),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_177),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_178),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_169),
.Y(n_177)
);

AOI32xp33_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_138),
.A3(n_134),
.B1(n_132),
.B2(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_167),
.C(n_166),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_171),
.C(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_158),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_179),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_156),
.B(n_172),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_190),
.B(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_192),
.B(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_185),
.B1(n_157),
.B2(n_180),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_176),
.B(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_163),
.B(n_141),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_16),
.B(n_19),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_25),
.B1(n_32),
.B2(n_35),
.C(n_36),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_38),
.Y(n_198)
);


endmodule