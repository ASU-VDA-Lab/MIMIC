module fake_jpeg_19094_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_7;
wire n_66;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_26)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_16),
.C(n_9),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_21),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

OAI211xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_28),
.B(n_13),
.C(n_8),
.Y(n_44)
);

XNOR2x1_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_11),
.Y(n_45)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.C(n_34),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_7),
.B(n_20),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_46),
.CI(n_11),
.CON(n_53),
.SN(n_53)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_48),
.B(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_11),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_20),
.B(n_31),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_24),
.B(n_11),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_0),
.Y(n_60)
);

OAI321xp33_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_50),
.A3(n_54),
.B1(n_58),
.B2(n_16),
.C(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_23),
.B1(n_6),
.B2(n_4),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_64),
.B1(n_23),
.B2(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_6),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_1),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_10),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_10),
.C(n_9),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.C(n_1),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_3),
.B(n_4),
.Y(n_76)
);


endmodule