module fake_aes_6612_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_2), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_12), .B(n_0), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_8), .B(n_13), .Y(n_16) );
O2A1O1Ixp33_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_2), .B(n_3), .C(n_5), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_17), .A2(n_9), .B1(n_10), .B2(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_18), .B(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AOI21xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_20), .B(n_13), .Y(n_23) );
CKINVDCx14_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
AOI21xp33_ASAP7_75t_SL g25 ( .A1(n_22), .A2(n_20), .B(n_5), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_11), .B1(n_6), .B2(n_3), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_11), .B1(n_24), .B2(n_27), .Y(n_29) );
endmodule