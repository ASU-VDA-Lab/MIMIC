module fake_jpeg_27022_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_10),
.B(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_49),
.B1(n_25),
.B2(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_23),
.B1(n_38),
.B2(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_20),
.B1(n_30),
.B2(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_36),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_74),
.B(n_78),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_63),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_28),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_23),
.B1(n_36),
.B2(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_78),
.B1(n_52),
.B2(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_26),
.B(n_30),
.C(n_25),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_24),
.B(n_17),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_75),
.Y(n_105)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_24),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_104),
.B(n_79),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_85),
.A2(n_90),
.B1(n_99),
.B2(n_17),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_52),
.B1(n_40),
.B2(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_27),
.C(n_33),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_33),
.C(n_27),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_18),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_22),
.Y(n_136)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_125),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_117),
.B(n_119),
.Y(n_150)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_81),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_140),
.B(n_94),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_59),
.B(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_129),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_124),
.B1(n_2),
.B2(n_3),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_67),
.B1(n_77),
.B2(n_76),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_138),
.B1(n_87),
.B2(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_134),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_73),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_137),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_94),
.B1(n_92),
.B2(n_100),
.Y(n_145)
);

NOR2x1_ASAP7_75t_R g134 ( 
.A(n_99),
.B(n_29),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_27),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_107),
.B1(n_110),
.B2(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_21),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_108),
.B1(n_84),
.B2(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_27),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_29),
.B(n_1),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_142),
.A2(n_145),
.B(n_148),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_118),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_157),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_97),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_88),
.B1(n_110),
.B2(n_86),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_170),
.B1(n_115),
.B2(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_169),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_86),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_166),
.B(n_2),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_111),
.C(n_109),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.C(n_122),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_109),
.C(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_134),
.B1(n_117),
.B2(n_114),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_123),
.B1(n_129),
.B2(n_125),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_176),
.B(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_126),
.B1(n_122),
.B2(n_115),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_191),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_113),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_188),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_11),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_199),
.B(n_202),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_3),
.C(n_4),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_200),
.C(n_166),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_141),
.B1(n_172),
.B2(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_6),
.C(n_7),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_6),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_142),
.B(n_7),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_154),
.C(n_144),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_206),
.B(n_208),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_158),
.C(n_155),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_148),
.B(n_150),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_213),
.B1(n_184),
.B2(n_182),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_186),
.B1(n_184),
.B2(n_197),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_169),
.B1(n_147),
.B2(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_150),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_154),
.C(n_168),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_176),
.C(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_203),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_178),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_188),
.C(n_175),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_234),
.C(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_192),
.C(n_177),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_196),
.Y(n_236)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_148),
.B1(n_190),
.B2(n_202),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_243),
.B1(n_212),
.B2(n_210),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_194),
.B1(n_200),
.B2(n_9),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_252),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_205),
.B(n_226),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_213),
.C(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_254),
.C(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_220),
.C(n_217),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_219),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_209),
.C(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_262),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_209),
.CI(n_223),
.CON(n_260),
.SN(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_204),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_255),
.B1(n_210),
.B2(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_243),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_240),
.B1(n_246),
.B2(n_238),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_272),
.B1(n_242),
.B2(n_244),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_240),
.B1(n_238),
.B2(n_245),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_237),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_8),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_251),
.B(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_244),
.B1(n_258),
.B2(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_221),
.CI(n_248),
.CON(n_281),
.SN(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_284),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_253),
.C(n_221),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_270),
.C(n_285),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_204),
.B(n_253),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_7),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_8),
.B(n_9),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_264),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_278),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_289),
.C(n_267),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_297),
.Y(n_306)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_305),
.B(n_304),
.C(n_294),
.D(n_296),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_281),
.B(n_284),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_8),
.Y(n_311)
);


endmodule