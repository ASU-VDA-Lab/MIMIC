module fake_jpeg_2215_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_25),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_23),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_24),
.B1(n_19),
.B2(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_27),
.B1(n_16),
.B2(n_18),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_22),
.C(n_20),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.C(n_0),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_17),
.C(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.C(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx24_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_45),
.C(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_14),
.C(n_13),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.C(n_4),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_12),
.C(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_2),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_5),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_50),
.B(n_6),
.Y(n_53)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_5),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_7),
.Y(n_55)
);


endmodule