module fake_jpeg_22551_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_14),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_31),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_58),
.B(n_68),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_62),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_31),
.C(n_21),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_56),
.Y(n_85)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_55),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_21),
.Y(n_56)
);

NOR4xp25_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_24),
.B2(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_71),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_22),
.C(n_16),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_5),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_91),
.B1(n_92),
.B2(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_27),
.B1(n_26),
.B2(n_19),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_97),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_7),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_50),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_93),
.C(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_113),
.C(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_58),
.B(n_52),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_75),
.B(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_68),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_95),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_74),
.C(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_57),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_121),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_74),
.C(n_60),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_79),
.C(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_60),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_83),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_83),
.B1(n_64),
.B2(n_77),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_131),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_86),
.B(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_141),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_102),
.B(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.C(n_133),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_92),
.B(n_46),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_111),
.B1(n_119),
.B2(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_136),
.B1(n_120),
.B2(n_108),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_80),
.B(n_75),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_46),
.B(n_59),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_135),
.C(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_83),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_97),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_77),
.C(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_115),
.C(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_135),
.B1(n_126),
.B2(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

AO221x1_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_103),
.B1(n_81),
.B2(n_130),
.C(n_64),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_120),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_127),
.B(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_108),
.B(n_114),
.C(n_101),
.D(n_109),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.C(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_162),
.B1(n_164),
.B2(n_160),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_164),
.B(n_141),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_123),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_126),
.C(n_140),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_152),
.C(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_151),
.C(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_145),
.C(n_155),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_174),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_156),
.B1(n_130),
.B2(n_136),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_181),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_161),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_169),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_165),
.B(n_154),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_173),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_185),
.A3(n_179),
.B1(n_84),
.B2(n_90),
.C1(n_109),
.C2(n_50),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_179),
.A3(n_84),
.B1(n_14),
.B2(n_11),
.C1(n_64),
.C2(n_9),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_178),
.C(n_180),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.B(n_11),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_9),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule