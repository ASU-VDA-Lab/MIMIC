module fake_jpeg_2071_n_565 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_565);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_11),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_60),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_19),
.B(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_62),
.Y(n_145)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_46),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_10),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_46),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_78),
.Y(n_116)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_19),
.B(n_10),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_80),
.B(n_104),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_13),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_89),
.Y(n_119)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_92),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_97),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_13),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_98),
.B(n_48),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_21),
.B(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_105),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_118),
.B1(n_124),
.B2(n_134),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_36),
.B1(n_49),
.B2(n_28),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_122),
.A2(n_130),
.B1(n_158),
.B2(n_165),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_32),
.B1(n_43),
.B2(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_73),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_30),
.B1(n_49),
.B2(n_23),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_55),
.A2(n_32),
.B1(n_43),
.B2(n_42),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_59),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_139),
.A2(n_151),
.B1(n_163),
.B2(n_25),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_146)
);

AO22x2_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_65),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_56),
.A2(n_49),
.B1(n_38),
.B2(n_31),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_67),
.A2(n_21),
.B1(n_27),
.B2(n_26),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_66),
.A2(n_28),
.B1(n_25),
.B2(n_38),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_79),
.A2(n_24),
.B(n_22),
.C(n_28),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_168),
.B(n_23),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_69),
.A2(n_48),
.B1(n_47),
.B2(n_24),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_95),
.B1(n_38),
.B2(n_31),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

AND2x4_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_93),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_170),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_174),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_114),
.B(n_105),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_175),
.B(n_177),
.Y(n_277)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_180),
.B(n_184),
.Y(n_234)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_181),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_185),
.A2(n_20),
.B(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_186),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_62),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_187),
.B(n_204),
.Y(n_252)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_188),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_118),
.B1(n_119),
.B2(n_71),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_189),
.A2(n_191),
.B1(n_198),
.B2(n_217),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_150),
.B1(n_157),
.B2(n_149),
.Y(n_244)
);

NAND2xp67_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_31),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_209),
.Y(n_276)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_195),
.A2(n_211),
.B1(n_221),
.B2(n_222),
.Y(n_247)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_104),
.B1(n_102),
.B2(n_101),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_30),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_203),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_109),
.B(n_160),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_205),
.B(n_206),
.Y(n_243)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_207),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_140),
.B(n_75),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_0),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_212),
.Y(n_233)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_126),
.B(n_91),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_92),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_164),
.B(n_57),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_151),
.A2(n_81),
.B1(n_96),
.B2(n_76),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_147),
.B(n_98),
.C(n_47),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_126),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_92),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_121),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_146),
.A2(n_88),
.B1(n_61),
.B2(n_84),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_20),
.B(n_1),
.Y(n_259)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_224),
.A2(n_229),
.B1(n_230),
.B2(n_0),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_137),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_141),
.B(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_228),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_126),
.B(n_14),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_131),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_193),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_175),
.A2(n_161),
.B1(n_157),
.B2(n_149),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_244),
.B1(n_251),
.B2(n_260),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_192),
.A2(n_108),
.B(n_142),
.C(n_144),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_248),
.A2(n_271),
.B(n_4),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_175),
.A2(n_148),
.B1(n_143),
.B2(n_136),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_172),
.A2(n_142),
.B1(n_131),
.B2(n_135),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_253),
.A2(n_258),
.B1(n_182),
.B2(n_222),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_135),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_177),
.B(n_143),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_148),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_274),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_178),
.A2(n_136),
.B1(n_137),
.B2(n_121),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_223),
.A2(n_20),
.B1(n_1),
.B2(n_0),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_171),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_270),
.B1(n_282),
.B2(n_260),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_178),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_14),
.B(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_170),
.A2(n_190),
.B1(n_191),
.B2(n_197),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_190),
.B1(n_174),
.B2(n_173),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_188),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_170),
.A2(n_4),
.B(n_5),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_179),
.B(n_221),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_284),
.B(n_288),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_285),
.A2(n_289),
.B1(n_314),
.B2(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_286),
.B(n_298),
.Y(n_348)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_190),
.B1(n_194),
.B2(n_227),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_233),
.B(n_216),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_301),
.Y(n_334)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_181),
.B1(n_176),
.B2(n_206),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_296),
.A2(n_313),
.B1(n_330),
.B2(n_269),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_302),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_275),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_169),
.B(n_212),
.C(n_230),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_229),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_303),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_211),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_309),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_325),
.Y(n_332)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_233),
.B(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_207),
.C(n_199),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_328),
.C(n_235),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_236),
.A2(n_224),
.B1(n_196),
.B2(n_203),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_241),
.Y(n_316)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_247),
.A2(n_4),
.B1(n_5),
.B2(n_14),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_319),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_231),
.B(n_18),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_255),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_241),
.B(n_263),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g323 ( 
.A(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_240),
.B(n_4),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_326),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_239),
.B(n_231),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_249),
.B(n_5),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_265),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_329),
.B1(n_232),
.B2(n_280),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_238),
.B(n_15),
.C(n_16),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_240),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_264),
.A2(n_15),
.B1(n_17),
.B2(n_244),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_323),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_248),
.B(n_242),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_362),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_276),
.B(n_249),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g409 ( 
.A1(n_339),
.A2(n_360),
.B(n_371),
.Y(n_409)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_309),
.A2(n_250),
.A3(n_251),
.B1(n_268),
.B2(n_278),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_250),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_365),
.C(n_372),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_308),
.A2(n_259),
.B1(n_271),
.B2(n_243),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_343),
.A2(n_345),
.B1(n_352),
.B2(n_368),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_308),
.A2(n_259),
.B1(n_267),
.B2(n_257),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_270),
.B1(n_245),
.B2(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_359),
.B(n_298),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_297),
.A2(n_246),
.B(n_263),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_299),
.B(n_312),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_278),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_285),
.A2(n_283),
.B(n_261),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_366),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_305),
.B(n_262),
.C(n_266),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_262),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_292),
.B(n_261),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_337),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_291),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_322),
.A2(n_232),
.B(n_266),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_280),
.C(n_245),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_351),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_388),
.Y(n_423)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_377),
.A2(n_360),
.B(n_336),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_354),
.A2(n_313),
.B1(n_299),
.B2(n_292),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_400),
.B1(n_335),
.B2(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_348),
.A2(n_317),
.B(n_287),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_382),
.A2(n_385),
.B(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_321),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_398),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_SL g385 ( 
.A(n_332),
.B(n_327),
.C(n_289),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_391),
.C(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_390),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_353),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_361),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_290),
.C(n_284),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_399),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_324),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_304),
.C(n_293),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_403),
.C(n_339),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_320),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_396),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_397),
.B(n_334),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_354),
.A2(n_333),
.B1(n_357),
.B2(n_362),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_355),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_401),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_340),
.B(n_295),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_402),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_294),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_366),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_364),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_345),
.A2(n_296),
.B1(n_314),
.B2(n_318),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_410),
.Y(n_416)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_400),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_392),
.A2(n_333),
.B1(n_357),
.B2(n_334),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_412),
.A2(n_421),
.B1(n_437),
.B2(n_438),
.Y(n_461)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_419),
.A2(n_426),
.B1(n_428),
.B2(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_422),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_392),
.A2(n_336),
.B1(n_340),
.B2(n_338),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_336),
.B1(n_352),
.B2(n_364),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_427),
.A2(n_433),
.B(n_434),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_380),
.A2(n_335),
.B1(n_338),
.B2(n_369),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_341),
.Y(n_430)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_372),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_441),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_390),
.A2(n_358),
.B(n_356),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_370),
.B(n_316),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_358),
.Y(n_435)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_380),
.A2(n_374),
.B1(n_373),
.B2(n_370),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_378),
.A2(n_374),
.B1(n_373),
.B2(n_349),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_378),
.A2(n_349),
.B1(n_347),
.B2(n_307),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_407),
.A2(n_347),
.B1(n_315),
.B2(n_310),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_412),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_389),
.B(n_329),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_391),
.C(n_403),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_424),
.C(n_422),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_331),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_470),
.Y(n_478)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_420),
.B(n_397),
.CI(n_384),
.CON(n_454),
.SN(n_454)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_469),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_394),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_458),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_438),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_430),
.B1(n_436),
.B2(n_426),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_398),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_467),
.Y(n_480)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_415),
.Y(n_463)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_418),
.B(n_383),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_418),
.B(n_377),
.CI(n_409),
.CON(n_469),
.SN(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_385),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_416),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_472),
.Y(n_495)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_448),
.A2(n_428),
.B(n_419),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_461),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_475),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_417),
.B1(n_414),
.B2(n_434),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_479),
.A2(n_445),
.B1(n_462),
.B2(n_471),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_441),
.C(n_425),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_481),
.B(n_484),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_468),
.A2(n_421),
.B1(n_440),
.B2(n_439),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_492),
.B1(n_496),
.B2(n_457),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_413),
.C(n_375),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_448),
.A2(n_427),
.B(n_414),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_493),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_413),
.C(n_437),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_494),
.C(n_462),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_452),
.A2(n_410),
.B1(n_431),
.B2(n_444),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_443),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_381),
.C(n_444),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_449),
.A2(n_393),
.B1(n_408),
.B2(n_399),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_504),
.Y(n_518)
);

AOI22x1_ASAP7_75t_L g527 ( 
.A1(n_498),
.A2(n_454),
.B1(n_387),
.B2(n_477),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_452),
.Y(n_499)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_499),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_496),
.Y(n_502)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_470),
.C(n_447),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_447),
.C(n_445),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_507),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_476),
.B(n_457),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_479),
.B1(n_482),
.B2(n_483),
.Y(n_515)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_511),
.Y(n_526)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_473),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_490),
.A2(n_472),
.B1(n_453),
.B2(n_411),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_512),
.A2(n_488),
.B1(n_487),
.B2(n_480),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_491),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_17),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_515),
.Y(n_531)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_514),
.A2(n_489),
.B1(n_488),
.B2(n_487),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_524),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_485),
.B1(n_474),
.B2(n_484),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_522),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_505),
.A2(n_485),
.B1(n_469),
.B2(n_486),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_499),
.A2(n_469),
.B1(n_481),
.B2(n_454),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_506),
.Y(n_538)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_527),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_323),
.B1(n_477),
.B2(n_306),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_528),
.A2(n_510),
.B1(n_513),
.B2(n_529),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_497),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_523),
.A2(n_501),
.B(n_522),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_532),
.A2(n_525),
.B(n_521),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_518),
.B(n_504),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_533),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_539),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_510),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_521),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_518),
.B(n_523),
.C(n_519),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_542),
.B(n_543),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_530),
.B(n_515),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_544),
.A2(n_545),
.B(n_548),
.Y(n_554)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_536),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_535),
.B(n_526),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_526),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_552),
.A2(n_547),
.B(n_538),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_550),
.A2(n_541),
.B1(n_531),
.B2(n_540),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_555),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_549),
.B(n_541),
.C(n_539),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_528),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_546),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_558),
.B(n_555),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_559),
.A2(n_554),
.B(n_553),
.Y(n_561)
);

BUFx24_ASAP7_75t_SL g562 ( 
.A(n_560),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_561),
.Y(n_563)
);

BUFx24_ASAP7_75t_SL g564 ( 
.A(n_563),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_557),
.C(n_527),
.Y(n_565)
);


endmodule