module fake_jpeg_24126_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_38),
.B(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_34),
.B1(n_29),
.B2(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

NOR2x1_ASAP7_75t_R g102 ( 
.A(n_52),
.B(n_72),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_31),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_18),
.C(n_31),
.Y(n_60)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_31),
.CI(n_32),
.CON(n_87),
.SN(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_35),
.B1(n_16),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_69),
.B1(n_74),
.B2(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_73),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_16),
.B1(n_17),
.B2(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_34),
.B1(n_28),
.B2(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_22),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_40),
.B1(n_45),
.B2(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_99),
.B1(n_117),
.B2(n_65),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_120),
.Y(n_137)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_115),
.Y(n_132)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_108),
.B1(n_113),
.B2(n_75),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_45),
.B1(n_28),
.B2(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_107),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_45),
.B(n_51),
.C(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_112),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_24),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_57),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_22),
.B1(n_48),
.B2(n_30),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_53),
.B(n_30),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_56),
.B(n_30),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_55),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_118),
.C(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_59),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_144),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_60),
.B1(n_55),
.B2(n_82),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_136),
.B1(n_152),
.B2(n_100),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_91),
.B1(n_143),
.B2(n_101),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_52),
.B1(n_65),
.B2(n_72),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_72),
.B(n_1),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_151),
.B(n_94),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_143),
.Y(n_153)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_83),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_118),
.B(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_105),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_56),
.B1(n_67),
.B2(n_3),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_68),
.B1(n_67),
.B2(n_3),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_154),
.B(n_160),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_166),
.C(n_168),
.Y(n_188)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_159),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_163),
.B(n_164),
.Y(n_190)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_171),
.B1(n_111),
.B2(n_147),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_87),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_87),
.C(n_106),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_182),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_112),
.B1(n_86),
.B2(n_113),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_172),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_151),
.B1(n_135),
.B2(n_125),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_123),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_181),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_91),
.A3(n_103),
.B1(n_86),
.B2(n_93),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_110),
.C(n_96),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_122),
.C(n_132),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_15),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_126),
.B(n_0),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_186),
.Y(n_198)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_185),
.Y(n_210)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_147),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_137),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_193),
.B(n_156),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_208),
.C(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_186),
.B1(n_139),
.B2(n_130),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_204),
.B1(n_172),
.B2(n_160),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_203),
.B1(n_212),
.B2(n_215),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_137),
.B1(n_136),
.B2(n_145),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_168),
.A2(n_164),
.B1(n_161),
.B2(n_176),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_132),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_206),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_141),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_198),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_141),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_144),
.B1(n_148),
.B2(n_138),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_138),
.C(n_133),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_220),
.B(n_216),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_154),
.A2(n_2),
.B(n_3),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_240),
.B(n_247),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_209),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_233),
.B(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_171),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_196),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_195),
.B1(n_203),
.B2(n_202),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_243),
.B1(n_246),
.B2(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_159),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_241),
.B(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_165),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_162),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_183),
.B(n_170),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_4),
.B(n_5),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_153),
.C(n_184),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_193),
.C(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_191),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_256),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_224),
.A2(n_215),
.B1(n_200),
.B2(n_190),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_224),
.B1(n_240),
.B2(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_232),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_204),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_257),
.A2(n_259),
.B1(n_264),
.B2(n_266),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_192),
.B(n_207),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_261),
.Y(n_285)
);

OAI22x1_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_220),
.B1(n_206),
.B2(n_208),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_205),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_222),
.C(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_201),
.B1(n_185),
.B2(n_199),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_11),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_11),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_234),
.B(n_4),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_9),
.Y(n_289)
);

AOI22x1_ASAP7_75t_SL g271 ( 
.A1(n_221),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_268),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_245),
.B1(n_236),
.B2(n_235),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_279),
.B1(n_283),
.B2(n_286),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_249),
.B(n_263),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_277),
.A2(n_10),
.B(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_282),
.C(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_230),
.B1(n_227),
.B2(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_229),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_287),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_231),
.C(n_229),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_226),
.B1(n_7),
.B2(n_8),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_261),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_251),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_286)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_299),
.C(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_294),
.C(n_299),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_253),
.C(n_256),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_253),
.C(n_267),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_266),
.B1(n_271),
.B2(n_265),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_305),
.B1(n_272),
.B2(n_301),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_10),
.B(n_275),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_298),
.B(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_285),
.B1(n_279),
.B2(n_280),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_280),
.C(n_285),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_314),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_284),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_10),
.B1(n_272),
.B2(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_311),
.B(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_300),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_292),
.Y(n_324)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_307),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_331),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_312),
.B1(n_309),
.B2(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_334),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_307),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_331),
.B(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_308),
.B(n_333),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_335),
.C(n_325),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_340),
.C(n_323),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_321),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_321),
.Y(n_345)
);


endmodule