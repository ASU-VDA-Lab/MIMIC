module fake_jpeg_29838_n_500 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_500);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_85),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_88),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_94),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_29),
.B(n_9),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_47),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_110),
.B(n_118),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_111),
.B(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_61),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_32),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_139),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_41),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_122),
.B(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_45),
.C(n_43),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_23),
.C(n_48),
.Y(n_169)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_57),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_49),
.B(n_27),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_30),
.B1(n_45),
.B2(n_43),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_48),
.B1(n_20),
.B2(n_23),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_120),
.B1(n_89),
.B2(n_90),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_27),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_78),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_52),
.B(n_42),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_0),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_39),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_160),
.B(n_15),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_162),
.B(n_173),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_163),
.Y(n_231)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g265 ( 
.A(n_164),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_112),
.A2(n_63),
.B1(n_79),
.B2(n_70),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_184),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_112),
.A2(n_70),
.B1(n_30),
.B2(n_18),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_179),
.Y(n_253)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

CKINVDCx11_ASAP7_75t_R g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_136),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_58),
.B1(n_71),
.B2(n_69),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_102),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_176),
.B(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_30),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_113),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_73),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_108),
.B(n_17),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_182),
.B(n_186),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_31),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_16),
.Y(n_186)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_99),
.B(n_65),
.C(n_59),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_140),
.C(n_124),
.Y(n_223)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_100),
.A2(n_48),
.B1(n_20),
.B2(n_62),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_192),
.A2(n_203),
.B1(n_208),
.B2(n_215),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

BUFx16f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_146),
.B1(n_140),
.B2(n_124),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx12_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_205),
.Y(n_249)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_156),
.B1(n_107),
.B2(n_146),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_12),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_95),
.B1(n_86),
.B2(n_13),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_142),
.B(n_17),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_214),
.Y(n_256)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_127),
.B(n_16),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_147),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_215)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_221),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_135),
.B1(n_156),
.B2(n_116),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_220),
.A2(n_166),
.B1(n_163),
.B2(n_165),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_248),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_254),
.B1(n_264),
.B2(n_166),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_117),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_185),
.A2(n_117),
.B1(n_116),
.B2(n_114),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_185),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_180),
.B(n_0),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_187),
.B(n_6),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_1),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_175),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_185),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_169),
.C(n_189),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_266),
.B(n_282),
.C(n_235),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_226),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_267),
.B(n_268),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_160),
.Y(n_268)
);

AO21x2_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_257),
.B(n_263),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_272),
.A2(n_265),
.B1(n_240),
.B2(n_250),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_197),
.C(n_161),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_274),
.B(n_304),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_191),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_277),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_278),
.B(n_280),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_279),
.A2(n_292),
.B1(n_300),
.B2(n_238),
.Y(n_312)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_194),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_170),
.C(n_172),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_203),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_202),
.B(n_194),
.C(n_179),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_238),
.B(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_233),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_293),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_232),
.A2(n_211),
.B1(n_207),
.B2(n_204),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_290),
.A2(n_243),
.B1(n_241),
.B2(n_235),
.Y(n_315)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_291),
.B(n_295),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_247),
.A2(n_216),
.B1(n_190),
.B2(n_206),
.Y(n_292)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_201),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_305),
.Y(n_333)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

CKINVDCx12_ASAP7_75t_R g298 ( 
.A(n_231),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_298),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_256),
.B(n_164),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_299),
.B(n_302),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_247),
.A2(n_213),
.B1(n_199),
.B2(n_209),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_227),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_301),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_261),
.B(n_195),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_255),
.A2(n_195),
.B(n_165),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_307),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_163),
.C(n_3),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_1),
.Y(n_305)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_252),
.B(n_251),
.Y(n_317)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_223),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_320),
.C(n_321),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_264),
.B(n_219),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_311),
.A2(n_318),
.B(n_343),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_284),
.B1(n_270),
.B2(n_290),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_315),
.A2(n_344),
.B1(n_284),
.B2(n_296),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_324),
.B(n_303),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_271),
.B(n_252),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_245),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_282),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_328),
.B(n_330),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_241),
.C(n_228),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_273),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_332),
.A2(n_335),
.B(n_288),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_225),
.C(n_240),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_268),
.A2(n_262),
.B(n_260),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_270),
.A2(n_225),
.B1(n_237),
.B2(n_262),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_293),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_350),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_229),
.B1(n_4),
.B2(n_5),
.Y(n_404)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_325),
.B(n_316),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_352),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_319),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_364),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_323),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_354),
.A2(n_355),
.B(n_304),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_356),
.B(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_276),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_362),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_374),
.B1(n_312),
.B2(n_322),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_267),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_314),
.B(n_281),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_363),
.B(n_365),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_319),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_333),
.B(n_295),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_333),
.B(n_280),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_366),
.B(n_372),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_283),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_368),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_289),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_370),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_343),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_310),
.B(n_307),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_375),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_313),
.B(n_294),
.Y(n_372)
);

CKINVDCx10_ASAP7_75t_R g373 ( 
.A(n_326),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_285),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_319),
.A2(n_310),
.B(n_332),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_311),
.B(n_330),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_377),
.A2(n_386),
.B(n_392),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_399),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_335),
.B1(n_344),
.B2(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_380),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_308),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_401),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_321),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_385),
.B(n_394),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_376),
.A2(n_324),
.B(n_318),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_328),
.C(n_320),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_364),
.C(n_353),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_355),
.A2(n_340),
.B(n_286),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_352),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_340),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_397),
.B(n_403),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_358),
.A2(n_315),
.B1(n_306),
.B2(n_291),
.Y(n_398)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_398),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_360),
.A2(n_287),
.B1(n_275),
.B2(n_260),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_297),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_228),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_404),
.A2(n_352),
.B1(n_229),
.B2(n_5),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_411),
.C(n_416),
.Y(n_436)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_370),
.C(n_346),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_379),
.A2(n_365),
.B(n_371),
.Y(n_412)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_351),
.B1(n_366),
.B2(n_354),
.Y(n_414)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_374),
.C(n_371),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_349),
.C(n_362),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_419),
.C(n_386),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_395),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_423),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_375),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_421),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_396),
.A2(n_350),
.B1(n_369),
.B2(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

HB1xp67_ASAP7_75t_SL g424 ( 
.A(n_392),
.Y(n_424)
);

XNOR2x1_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_404),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_383),
.Y(n_427)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_427),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_400),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_402),
.Y(n_438)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_401),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_441),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_439),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_382),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_408),
.C(n_407),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_413),
.A2(n_402),
.B1(n_393),
.B2(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_403),
.C(n_400),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_447),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_406),
.A2(n_400),
.B1(n_384),
.B2(n_389),
.Y(n_446)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_405),
.A2(n_3),
.B1(n_399),
.B2(n_421),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_455),
.Y(n_469)
);

A2O1A1O1Ixp25_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_420),
.B(n_412),
.C(n_419),
.D(n_409),
.Y(n_450)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_416),
.C(n_408),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_451),
.B(n_462),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g455 ( 
.A1(n_429),
.A2(n_420),
.B(n_405),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_410),
.Y(n_456)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_431),
.Y(n_457)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_457),
.Y(n_466)
);

INVx11_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_426),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_436),
.C(n_441),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_465),
.B(n_470),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_437),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_471),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_459),
.C(n_452),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_458),
.Y(n_471)
);

XNOR2x1_ASAP7_75t_SL g473 ( 
.A(n_450),
.B(n_442),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_446),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_463),
.A2(n_453),
.B1(n_456),
.B2(n_440),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_475),
.B(n_478),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_467),
.A2(n_443),
.B(n_455),
.Y(n_477)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_477),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_444),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_479),
.B(n_415),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_430),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_483),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_447),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_482),
.A2(n_469),
.B(n_473),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_464),
.B(n_434),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_487),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_476),
.A2(n_469),
.B(n_435),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_415),
.Y(n_491)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_491),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_479),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_492),
.A2(n_484),
.B(n_485),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_490),
.B(n_494),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_496),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_482),
.B(n_480),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_498),
.A2(n_492),
.B(n_466),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_499),
.Y(n_500)
);


endmodule