module fake_jpeg_29761_n_452 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_60),
.Y(n_103)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_87),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_99),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_36),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_35),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_48),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_21),
.C(n_36),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_113),
.B(n_42),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_39),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_118),
.B(n_48),
.Y(n_201)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_44),
.B1(n_29),
.B2(n_30),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_140),
.B1(n_27),
.B2(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_64),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_69),
.A2(n_30),
.B1(n_17),
.B2(n_15),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_99),
.B1(n_87),
.B2(n_84),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_39),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_26),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_70),
.A2(n_35),
.B1(n_46),
.B2(n_45),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_45),
.B1(n_98),
.B2(n_48),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_51),
.Y(n_183)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_165),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_186),
.B1(n_152),
.B2(n_109),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_85),
.B1(n_28),
.B2(n_42),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_101),
.A2(n_83),
.B1(n_57),
.B2(n_56),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_177),
.Y(n_211)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_103),
.A2(n_93),
.B1(n_90),
.B2(n_88),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_180),
.B1(n_184),
.B2(n_189),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_103),
.A2(n_71),
.B1(n_82),
.B2(n_67),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_196),
.B1(n_197),
.B2(n_141),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_185),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_118),
.A2(n_63),
.B1(n_86),
.B2(n_52),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_116),
.A2(n_99),
.B1(n_87),
.B2(n_66),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_24),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_190),
.Y(n_222)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_108),
.A2(n_84),
.B1(n_66),
.B2(n_46),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_24),
.Y(n_190)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_192),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_199),
.B1(n_156),
.B2(n_141),
.Y(n_204)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_200),
.B1(n_201),
.B2(n_137),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_133),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_195),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_138),
.B1(n_131),
.B2(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_132),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_154),
.B1(n_124),
.B2(n_143),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_157),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_220),
.C(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_221),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_155),
.B(n_134),
.C(n_130),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_48),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_152),
.B1(n_154),
.B2(n_124),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_215),
.B1(n_216),
.B2(n_181),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_157),
.B(n_142),
.C(n_104),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_143),
.B1(n_128),
.B2(n_127),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_200),
.B1(n_170),
.B2(n_168),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_136),
.C(n_120),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_190),
.B(n_117),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_182),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_238),
.A2(n_242),
.B1(n_219),
.B2(n_224),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_164),
.B1(n_180),
.B2(n_183),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_239),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_183),
.B1(n_173),
.B2(n_185),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_184),
.B(n_201),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_245),
.B(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_165),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_163),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_210),
.C(n_225),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_198),
.B1(n_169),
.B2(n_192),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_250),
.B(n_255),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_171),
.B(n_160),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_253),
.B(n_230),
.Y(n_290)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

BUFx4f_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_159),
.B1(n_158),
.B2(n_166),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_259),
.B1(n_267),
.B2(n_214),
.Y(n_291)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_172),
.B1(n_162),
.B2(n_191),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_194),
.B(n_145),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_193),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_210),
.A2(n_188),
.B(n_175),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_31),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_222),
.A2(n_31),
.B1(n_15),
.B2(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_31),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_232),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_211),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_220),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_278),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_276),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_210),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_288),
.C(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_205),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

AO22x1_ASAP7_75t_SL g284 ( 
.A1(n_241),
.A2(n_216),
.B1(n_203),
.B2(n_207),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_207),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_239),
.B1(n_248),
.B2(n_255),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_268),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_238),
.B1(n_260),
.B2(n_257),
.Y(n_308)
);

AO21x2_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_224),
.B(n_219),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_261),
.B(n_262),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_241),
.A2(n_228),
.B1(n_218),
.B2(n_212),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_254),
.B1(n_258),
.B2(n_250),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_230),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_244),
.B(n_232),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_297),
.B(n_237),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_304),
.B(n_305),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_307),
.B1(n_317),
.B2(n_291),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_243),
.B(n_261),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_242),
.B(n_264),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_319),
.B1(n_292),
.B2(n_286),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_267),
.C(n_246),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.C(n_311),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_251),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

AOI21x1_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_259),
.B(n_258),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_313),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_273),
.A2(n_265),
.B(n_228),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_214),
.B1(n_236),
.B2(n_227),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_236),
.B1(n_212),
.B2(n_229),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_229),
.C(n_235),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_275),
.C(n_269),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_279),
.B(n_269),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_290),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_326),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_278),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_308),
.B1(n_319),
.B2(n_303),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_333),
.C(n_340),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_287),
.C(n_285),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_284),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_337),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_285),
.C(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_292),
.C(n_276),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_350),
.C(n_346),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_346),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_345),
.A2(n_31),
.B1(n_15),
.B2(n_3),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_298),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_306),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_295),
.C(n_237),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_352),
.B(n_362),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_371),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_356),
.A2(n_358),
.B1(n_333),
.B2(n_350),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_322),
.C(n_298),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_370),
.C(n_335),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_303),
.B1(n_313),
.B2(n_305),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_316),
.B1(n_307),
.B2(n_302),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_372),
.B1(n_338),
.B2(n_331),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_323),
.B(n_304),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_336),
.A2(n_300),
.B(n_314),
.C(n_306),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_369),
.B(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

XNOR2x2_ASAP7_75t_SL g367 ( 
.A(n_344),
.B(n_336),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_367),
.B(n_9),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_318),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_340),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_328),
.A2(n_317),
.B(n_295),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_318),
.C(n_286),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_293),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_330),
.A2(n_286),
.B1(n_293),
.B2(n_218),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_373),
.A2(n_339),
.B1(n_334),
.B2(n_341),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_374),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_355),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_377),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_376),
.A2(n_358),
.B1(n_356),
.B2(n_365),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_369),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_383),
.B1(n_387),
.B2(n_389),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_353),
.B1(n_364),
.B2(n_351),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_390),
.C(n_364),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_359),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_382),
.B(n_384),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_337),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_352),
.A2(n_347),
.B1(n_334),
.B2(n_325),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_357),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

AOI21x1_ASAP7_75t_SL g392 ( 
.A1(n_376),
.A2(n_365),
.B(n_367),
.Y(n_392)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_401),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_395),
.B(n_402),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_379),
.A2(n_365),
.B1(n_373),
.B2(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_397),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_377),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_375),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_351),
.C(n_353),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_0),
.C(n_1),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_385),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_10),
.B1(n_13),
.B2(n_4),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_404),
.A2(n_378),
.B1(n_390),
.B2(n_381),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_408),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_389),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_411),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_406),
.B(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_414),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_6),
.B1(n_13),
.B2(n_4),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_417),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_5),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_392),
.A2(n_6),
.B(n_11),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_418),
.A2(n_398),
.B(n_12),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_393),
.B(n_405),
.Y(n_421)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_421),
.A2(n_411),
.B(n_418),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_402),
.C(n_395),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_422),
.B(n_424),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_413),
.B(n_404),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_426),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_396),
.C(n_403),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_399),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_427),
.B(n_12),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_420),
.B(n_419),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_435),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_434),
.A2(n_430),
.B(n_424),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_416),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_409),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_438),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_437),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_417),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_431),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_443),
.A2(n_429),
.B1(n_427),
.B2(n_14),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_444),
.A2(n_445),
.B(n_446),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_439),
.A2(n_437),
.B(n_429),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_444),
.A2(n_442),
.B(n_440),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_447),
.B(n_0),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_450),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_3),
.B1(n_441),
.B2(n_449),
.Y(n_452)
);


endmodule