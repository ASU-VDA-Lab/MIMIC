module fake_jpeg_960_n_685 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_685);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_685;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_60),
.Y(n_185)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_71),
.Y(n_130)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_33),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_89),
.Y(n_151)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_88),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_35),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_93),
.Y(n_144)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_105),
.Y(n_153)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_24),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_24),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_103),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_0),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_106),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_111),
.Y(n_170)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_32),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_39),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_115),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_122),
.B(n_126),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

CKINVDCx11_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_47),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_38),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_62),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_137),
.B(n_203),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_55),
.C(n_52),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_44),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_52),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_143),
.B(n_195),
.Y(n_264)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_146),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_55),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_147),
.B(n_175),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_63),
.A2(n_49),
.B1(n_51),
.B2(n_40),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_154),
.A2(n_23),
.B1(n_101),
.B2(n_129),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_161),
.B(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_40),
.Y(n_175)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_70),
.A2(n_49),
.B1(n_42),
.B2(n_22),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_179),
.A2(n_209),
.B1(n_1),
.B2(n_2),
.Y(n_281)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_81),
.A2(n_54),
.B(n_41),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_189),
.A2(n_191),
.B(n_54),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_75),
.B(n_48),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_104),
.A2(n_121),
.B(n_128),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_67),
.B(n_48),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_94),
.B(n_45),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_78),
.B(n_45),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_92),
.A2(n_106),
.B1(n_123),
.B2(n_119),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_210),
.Y(n_284)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_98),
.Y(n_211)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_99),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_118),
.Y(n_226)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_112),
.Y(n_218)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_100),
.B(n_44),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

BUFx16f_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_225),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_227),
.Y(n_365)
);

CKINVDCx12_ASAP7_75t_R g229 ( 
.A(n_222),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_229),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_38),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_230),
.B(n_235),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_131),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

INVx6_ASAP7_75t_SL g234 ( 
.A(n_222),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_234),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_130),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_237),
.B(n_242),
.Y(n_315)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_240),
.Y(n_332)
);

CKINVDCx9p33_ASAP7_75t_R g241 ( 
.A(n_144),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_241),
.Y(n_321)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_174),
.B(n_41),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_247),
.B(n_251),
.Y(n_319)
);

CKINVDCx12_ASAP7_75t_R g248 ( 
.A(n_173),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_179),
.A2(n_42),
.B1(n_22),
.B2(n_37),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_249),
.A2(n_280),
.B(n_298),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_203),
.Y(n_250)
);

NAND2x1_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_151),
.B(n_166),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_151),
.B(n_37),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_257),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_255),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_153),
.B(n_25),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_153),
.B(n_25),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_262),
.Y(n_324)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

CKINVDCx9p33_ASAP7_75t_R g263 ( 
.A(n_147),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_198),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_275),
.Y(n_326)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_268),
.A2(n_296),
.B1(n_217),
.B2(n_168),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_155),
.Y(n_269)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_134),
.Y(n_270)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_134),
.Y(n_274)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_145),
.B(n_23),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_182),
.Y(n_276)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_276),
.Y(n_345)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_182),
.Y(n_278)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_278),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_143),
.B(n_0),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_279),
.B(n_285),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_195),
.A2(n_42),
.B1(n_124),
.B2(n_3),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_281),
.A2(n_295),
.B1(n_305),
.B2(n_139),
.Y(n_343)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_145),
.B(n_2),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_177),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_199),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_132),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_290),
.Y(n_357)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_149),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_141),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_291),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_152),
.B(n_16),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_301),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_294),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_209),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_140),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_198),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_297),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_160),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_163),
.B(n_7),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_300),
.A2(n_185),
.B1(n_172),
.B2(n_148),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_157),
.B(n_8),
.Y(n_301)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_159),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_303),
.Y(n_340)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_159),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_162),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_187),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_183),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_156),
.B1(n_201),
.B2(n_186),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_308),
.A2(n_311),
.B(n_343),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_263),
.A2(n_165),
.B(n_185),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_258),
.A2(n_180),
.B1(n_171),
.B2(n_164),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_339),
.B1(n_349),
.B2(n_351),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_256),
.A2(n_224),
.B(n_220),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_328),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_250),
.A2(n_176),
.B1(n_196),
.B2(n_202),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_250),
.A2(n_181),
.B(n_207),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_330),
.B(n_334),
.C(n_231),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_268),
.A2(n_238),
.B1(n_241),
.B2(n_291),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_274),
.B1(n_278),
.B2(n_276),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_149),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_252),
.A2(n_219),
.A3(n_214),
.B1(n_135),
.B2(n_133),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_240),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_237),
.A2(n_207),
.B1(n_193),
.B2(n_181),
.Y(n_339)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_237),
.A2(n_193),
.B1(n_217),
.B2(n_168),
.Y(n_349)
);

OAI22x1_ASAP7_75t_L g351 ( 
.A1(n_234),
.A2(n_204),
.B1(n_187),
.B2(n_184),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_354),
.A2(n_358),
.B1(n_359),
.B2(n_273),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_233),
.A2(n_139),
.B1(n_204),
.B2(n_13),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_270),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_264),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_296),
.A2(n_299),
.B1(n_267),
.B2(n_304),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_350),
.B(n_299),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_368),
.B(n_378),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_372),
.A2(n_375),
.B1(n_393),
.B2(n_408),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_325),
.B(n_333),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_374),
.B(n_377),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_261),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_381),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_228),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_326),
.B(n_243),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_379),
.A2(n_340),
.B1(n_321),
.B2(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_307),
.B(n_314),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

AO22x1_ASAP7_75t_SL g383 ( 
.A1(n_315),
.A2(n_254),
.B1(n_261),
.B2(n_244),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_383),
.B(n_392),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_355),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_389),
.Y(n_418)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_387),
.Y(n_425)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_347),
.B(n_266),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_390),
.B(n_398),
.Y(n_430)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_316),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_315),
.A2(n_302),
.B1(n_303),
.B2(n_239),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_315),
.B(n_225),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_401),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_314),
.B(n_254),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_404),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_286),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_319),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_399),
.B(n_406),
.Y(n_442)
);

BUFx12_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_316),
.B(n_236),
.Y(n_404)
);

INVx13_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_405),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_284),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_407),
.B(n_413),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_354),
.A2(n_244),
.B1(n_239),
.B2(n_236),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_308),
.Y(n_420)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_284),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_246),
.C(n_231),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_341),
.C(n_330),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_412),
.A2(n_327),
.B(n_328),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_417),
.A2(n_427),
.B(n_445),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_438),
.C(n_441),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_346),
.B1(n_339),
.B2(n_309),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_426),
.A2(n_436),
.B1(n_448),
.B2(n_450),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_412),
.A2(n_308),
.B(n_311),
.Y(n_427)
);

OAI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_428),
.A2(n_371),
.B1(n_376),
.B2(n_373),
.Y(n_463)
);

AO22x1_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_309),
.B1(n_308),
.B2(n_321),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_383),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_400),
.A2(n_311),
.B1(n_340),
.B2(n_318),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_344),
.C(n_324),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_400),
.A2(n_360),
.B1(n_356),
.B2(n_362),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_444),
.A2(n_393),
.B1(n_408),
.B2(n_383),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_395),
.A2(n_357),
.B(n_321),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_369),
.A2(n_395),
.B1(n_375),
.B2(n_371),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_363),
.C(n_337),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_451),
.C(n_441),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_369),
.A2(n_358),
.B1(n_353),
.B2(n_351),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_322),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_357),
.B(n_323),
.Y(n_454)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_414),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_455),
.Y(n_456)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_456),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_396),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_459),
.B(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_460),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_462),
.A2(n_463),
.B1(n_472),
.B2(n_479),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_416),
.B(n_378),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_464),
.Y(n_507)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_415),
.Y(n_465)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_465),
.Y(n_506)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

INVx13_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_467),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g468 ( 
.A(n_452),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_404),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_469),
.B(n_471),
.Y(n_495)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_470),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_407),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_425),
.A2(n_373),
.B1(n_379),
.B2(n_384),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_427),
.B(n_433),
.Y(n_494)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_475),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_476),
.A2(n_477),
.B1(n_436),
.B2(n_450),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_448),
.A2(n_389),
.B1(n_410),
.B2(n_380),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_418),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_424),
.A2(n_411),
.B1(n_394),
.B2(n_386),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_433),
.B1(n_443),
.B2(n_446),
.Y(n_500)
);

INVx13_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_490),
.Y(n_496)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_391),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_442),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_488),
.C(n_491),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_419),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_489),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_419),
.B(n_405),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_385),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_438),
.C(n_420),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_440),
.B(n_382),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_454),
.A2(n_402),
.B1(n_353),
.B2(n_332),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_492),
.A2(n_435),
.B1(n_367),
.B2(n_402),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_449),
.B(n_417),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_493),
.B(n_431),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_494),
.A2(n_478),
.B(n_462),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_500),
.A2(n_511),
.B1(n_519),
.B2(n_530),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_456),
.B(n_437),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_504),
.B(n_509),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_437),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_457),
.A2(n_424),
.B1(n_426),
.B2(n_444),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_458),
.B(n_446),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_524),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_479),
.B(n_332),
.Y(n_513)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_513),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_518),
.A2(n_489),
.B1(n_461),
.B2(n_477),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_457),
.A2(n_445),
.B1(n_431),
.B2(n_421),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_421),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_523),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_522),
.B(n_481),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_480),
.B(n_388),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_453),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_453),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_525),
.B(n_312),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_452),
.Y(n_526)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_526),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_485),
.B(n_435),
.Y(n_528)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_528),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_532),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_533),
.B(n_540),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_534),
.A2(n_536),
.B1(n_556),
.B2(n_557),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_480),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_535),
.B(n_563),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_518),
.A2(n_461),
.B1(n_478),
.B2(n_493),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_511),
.A2(n_476),
.B1(n_459),
.B2(n_473),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_539),
.A2(n_552),
.B1(n_530),
.B2(n_502),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_516),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_541),
.B(n_547),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_494),
.A2(n_473),
.B(n_491),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_543),
.Y(n_588)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_528),
.Y(n_544)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_544),
.Y(n_568)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_526),
.Y(n_545)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_545),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_521),
.B(n_484),
.C(n_475),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_529),
.C(n_527),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_516),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_495),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_548),
.B(n_551),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_460),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_558),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_505),
.A2(n_466),
.B(n_474),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_497),
.A2(n_470),
.B1(n_465),
.B2(n_468),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_505),
.B(n_468),
.Y(n_553)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_522),
.A2(n_482),
.B1(n_467),
.B2(n_310),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_554),
.A2(n_499),
.B1(n_514),
.B2(n_517),
.Y(n_575)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_503),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_498),
.A2(n_482),
.B(n_467),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_401),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_519),
.A2(n_310),
.B1(n_352),
.B2(n_306),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_559),
.A2(n_562),
.B1(n_506),
.B2(n_503),
.Y(n_586)
);

INVxp33_ASAP7_75t_SL g587 ( 
.A(n_561),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_507),
.A2(n_352),
.B1(n_306),
.B2(n_401),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_357),
.Y(n_563)
);

FAx1_ASAP7_75t_SL g564 ( 
.A(n_539),
.B(n_515),
.CI(n_498),
.CON(n_564),
.SN(n_564)
);

AOI31xp67_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_567),
.A3(n_568),
.B(n_542),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_531),
.B(n_515),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_565),
.B(n_576),
.Y(n_603)
);

FAx1_ASAP7_75t_SL g567 ( 
.A(n_532),
.B(n_500),
.CI(n_501),
.CON(n_567),
.SN(n_567)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_549),
.B(n_502),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_578),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_572),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_573),
.B(n_533),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_575),
.A2(n_581),
.B1(n_586),
.B2(n_589),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_531),
.B(n_529),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_535),
.B(n_527),
.C(n_517),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_510),
.C(n_508),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_579),
.B(n_590),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_538),
.A2(n_499),
.B1(n_510),
.B2(n_506),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_550),
.B(n_508),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_553),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_534),
.A2(n_557),
.B1(n_536),
.B2(n_563),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_560),
.B(n_312),
.Y(n_590)
);

AO221x1_ASAP7_75t_L g591 ( 
.A1(n_581),
.A2(n_559),
.B1(n_555),
.B2(n_541),
.C(n_552),
.Y(n_591)
);

AOI31xp33_ASAP7_75t_L g622 ( 
.A1(n_591),
.A2(n_594),
.A3(n_599),
.B(n_564),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_577),
.Y(n_593)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_593),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_SL g594 ( 
.A(n_588),
.B(n_544),
.C(n_542),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_546),
.C(n_543),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_596),
.B(n_607),
.C(n_610),
.Y(n_620)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_582),
.Y(n_598)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_598),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_585),
.A2(n_554),
.B(n_551),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_612),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_601),
.B(n_227),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_570),
.A2(n_545),
.B1(n_537),
.B2(n_556),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_602),
.B(n_604),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_574),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_573),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_255),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_387),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_537),
.C(n_401),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_585),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_609),
.B(n_580),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_579),
.B(n_246),
.C(n_365),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_611),
.B(n_583),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_225),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_569),
.B(n_269),
.C(n_232),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_565),
.C(n_567),
.Y(n_621)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_593),
.A2(n_566),
.B(n_588),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_615),
.A2(n_617),
.B(n_619),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_597),
.A2(n_566),
.B(n_584),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_618),
.A2(n_622),
.B1(n_626),
.B2(n_633),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_594),
.A2(n_567),
.B(n_564),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_623),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_329),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_624),
.B(n_632),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_595),
.B(n_403),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_625),
.B(n_630),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_611),
.A2(n_329),
.B1(n_260),
.B2(n_245),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_627),
.A2(n_272),
.B(n_289),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_596),
.B(n_290),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_592),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_628),
.B(n_600),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_634),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_628),
.B(n_603),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_636),
.B(n_642),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_610),
.C(n_603),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_637),
.B(n_638),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_620),
.B(n_613),
.C(n_293),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_617),
.A2(n_616),
.B1(n_619),
.B2(n_631),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_640),
.B(n_649),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_621),
.B(n_283),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_283),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_644),
.B(n_646),
.C(n_624),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_633),
.B(n_300),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_647),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_615),
.B(n_293),
.C(n_272),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_SL g650 ( 
.A(n_639),
.B(n_629),
.C(n_645),
.Y(n_650)
);

INVx11_ASAP7_75t_L g662 ( 
.A(n_650),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_635),
.B(n_630),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_651),
.B(n_656),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_653),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_643),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_654),
.B(n_655),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_629),
.C(n_626),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_646),
.B(n_623),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_636),
.C(n_642),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_659),
.B(n_660),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_SL g663 ( 
.A(n_661),
.B(n_648),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_663),
.B(n_669),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_658),
.B(n_647),
.C(n_649),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_666),
.B(n_667),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_657),
.B(n_644),
.C(n_294),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_657),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_670),
.B(n_15),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g671 ( 
.A1(n_669),
.A2(n_650),
.B(n_652),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_671),
.B(n_672),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_665),
.B(n_294),
.C(n_289),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_668),
.B(n_14),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_673),
.B(n_676),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_675),
.B(n_665),
.C(n_664),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_679),
.B(n_662),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_677),
.B(n_675),
.C(n_674),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_681),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_682),
.B(n_678),
.C(n_16),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_683),
.Y(n_684)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_16),
.Y(n_685)
);


endmodule