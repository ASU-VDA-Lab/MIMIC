module fake_jpeg_18884_n_379 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_8),
.B(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_14),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_1),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_21),
.C(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_29),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_25),
.B1(n_19),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_21),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_25),
.B1(n_19),
.B2(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_33),
.B1(n_22),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_26),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_33),
.B1(n_22),
.B2(n_24),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_38),
.A2(n_30),
.B(n_18),
.C(n_28),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_48),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_61),
.B1(n_44),
.B2(n_49),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_121),
.B1(n_92),
.B2(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_48),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_103),
.A2(n_83),
.B(n_64),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_79),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_119),
.Y(n_156)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_107),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_113),
.Y(n_150)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_34),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_122),
.Y(n_153)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_37),
.B1(n_56),
.B2(n_27),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_92),
.B1(n_73),
.B2(n_65),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_28),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_30),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_133),
.B1(n_88),
.B2(n_94),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_12),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

OR2x4_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_29),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_71),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_57),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_76),
.A2(n_29),
.B1(n_12),
.B2(n_11),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_139),
.B1(n_92),
.B2(n_88),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_76),
.A2(n_29),
.B1(n_12),
.B2(n_11),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_140),
.A2(n_152),
.B(n_164),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_136),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_145),
.B1(n_166),
.B2(n_168),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_173),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_161),
.A2(n_133),
.B1(n_104),
.B2(n_105),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_124),
.A2(n_94),
.B1(n_84),
.B2(n_35),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_84),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_113),
.B1(n_109),
.B2(n_114),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_189),
.B1(n_202),
.B2(n_130),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_137),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_181),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_100),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_182),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_197),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_101),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_107),
.B1(n_119),
.B2(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_103),
.B(n_128),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_201),
.B(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_100),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_192),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_121),
.C(n_134),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_157),
.C(n_127),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_141),
.B(n_123),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_143),
.B(n_146),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_208),
.B(n_159),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_147),
.B(n_102),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_110),
.B1(n_123),
.B2(n_118),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_156),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_103),
.B(n_162),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_145),
.B1(n_161),
.B2(n_156),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_212),
.B1(n_232),
.B2(n_202),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_140),
.B1(n_154),
.B2(n_173),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_162),
.C(n_146),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_192),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_214),
.A2(n_221),
.B(n_223),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_241),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_149),
.B(n_159),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_191),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_230),
.C(n_239),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_225),
.A2(n_210),
.B1(n_206),
.B2(n_196),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_157),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_115),
.B1(n_112),
.B2(n_172),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_149),
.B(n_170),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_170),
.B1(n_172),
.B2(n_163),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_179),
.B1(n_207),
.B2(n_184),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_127),
.C(n_163),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_68),
.C(n_132),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_177),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_177),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_197),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_250),
.A2(n_251),
.B(n_267),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_252),
.A2(n_263),
.B1(n_264),
.B2(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_260),
.B1(n_271),
.B2(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_185),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_201),
.Y(n_256)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_180),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_259),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_188),
.B1(n_194),
.B2(n_190),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_199),
.B1(n_195),
.B2(n_187),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_186),
.B1(n_204),
.B2(n_205),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_2),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_265),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_229),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_279),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_224),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_229),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_287),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_230),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_212),
.B1(n_215),
.B2(n_231),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_293),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_241),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_291),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_221),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_218),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_250),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_252),
.A2(n_233),
.B1(n_218),
.B2(n_231),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_249),
.C(n_260),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_295),
.C(n_270),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_214),
.C(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_247),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_237),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_310),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_307),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_305),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_266),
.B(n_240),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_273),
.C(n_272),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_309),
.C(n_289),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_284),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_315),
.B(n_317),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_266),
.B(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_319),
.B(n_263),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_294),
.B(n_276),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_324),
.B(n_331),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_275),
.B1(n_290),
.B2(n_287),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_319),
.B1(n_303),
.B2(n_318),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_334),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_280),
.B(n_292),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_285),
.C(n_274),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_314),
.C(n_316),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_274),
.B(n_275),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_305),
.A2(n_240),
.B(n_238),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_271),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_338),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_337),
.A2(n_341),
.B1(n_322),
.B2(n_340),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_307),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_309),
.B1(n_318),
.B2(n_245),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_316),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_345),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_347),
.Y(n_354)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_329),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_314),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_262),
.B(n_245),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_346),
.A2(n_325),
.B(n_321),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_226),
.B(n_238),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_6),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_348),
.B(n_330),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_334),
.B1(n_328),
.B2(n_331),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_351),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_348),
.B(n_326),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_353),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_6),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_L g359 ( 
.A1(n_350),
.A2(n_324),
.B1(n_320),
.B2(n_335),
.C(n_339),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_354),
.B(n_357),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_339),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_360),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_345),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_364),
.C(n_354),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_343),
.C(n_342),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_368),
.A2(n_6),
.B(n_7),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_371),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

NAND4xp25_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_365),
.C(n_361),
.D(n_363),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_372),
.A2(n_373),
.B(n_370),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_374),
.B1(n_8),
.B2(n_9),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_8),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_8),
.B1(n_9),
.B2(n_326),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_9),
.Y(n_379)
);


endmodule