module fake_jpeg_5443_n_152 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_47),
.Y(n_54)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_32),
.C(n_27),
.Y(n_61)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_2),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_41),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_55),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_27),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_14),
.Y(n_82)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_20),
.C(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_31),
.B1(n_8),
.B2(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_72),
.Y(n_94)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_22),
.B1(n_23),
.B2(n_18),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_15),
.B(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_61),
.B1(n_56),
.B2(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_109),
.B1(n_85),
.B2(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_108),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_55),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_51),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_57),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_91),
.C(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_58),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_114),
.C(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_101),
.C(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_118),
.C(n_109),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_93),
.C(n_96),
.Y(n_118)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_100),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_94),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_83),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_78),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_49),
.B1(n_63),
.B2(n_53),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_121),
.C(n_115),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_110),
.B(n_97),
.C(n_80),
.D(n_100),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_119),
.B(n_125),
.C(n_92),
.D(n_53),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.C(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_114),
.C(n_124),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_118),
.C(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_133),
.Y(n_140)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_139),
.A2(n_126),
.B(n_132),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_138),
.B(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_95),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.C(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_79),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.C(n_5),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_143),
.C(n_50),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_149),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_5),
.B(n_52),
.Y(n_152)
);


endmodule