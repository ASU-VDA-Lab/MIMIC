module fake_jpeg_11688_n_82 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_39),
.Y(n_42)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_13),
.B1(n_25),
.B2(n_24),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_32),
.B(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_45),
.B(n_6),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_38),
.C(n_14),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_17),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_7),
.B(n_8),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_53),
.B1(n_54),
.B2(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_68),
.B1(n_63),
.B2(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_76),
.B(n_74),
.Y(n_77)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_68),
.Y(n_79)
);

INVxp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_73),
.Y(n_82)
);


endmodule