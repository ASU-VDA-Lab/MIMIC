module fake_jpeg_24208_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_21),
.B1(n_31),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_54),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_29),
.B1(n_23),
.B2(n_32),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_67),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_36),
.B1(n_40),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_77),
.B1(n_81),
.B2(n_30),
.Y(n_107)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_65),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_32),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_78),
.B1(n_25),
.B2(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_82),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_1),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_37),
.B(n_34),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_28),
.B1(n_17),
.B2(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_30),
.B1(n_17),
.B2(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_88),
.B(n_3),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_37),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_101),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_106),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_84),
.B1(n_83),
.B2(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_52),
.C(n_41),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_59),
.C(n_52),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_117),
.B1(n_121),
.B2(n_94),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_57),
.B1(n_76),
.B2(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_77),
.B1(n_63),
.B2(n_76),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_127),
.B(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_63),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_59),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_92),
.B(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_101),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_146),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_97),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_127),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_87),
.B(n_97),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_144),
.B(n_145),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_115),
.B(n_136),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_108),
.B(n_106),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_104),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_103),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_161),
.B(n_116),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_107),
.A3(n_90),
.B1(n_95),
.B2(n_88),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_162),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_111),
.B(n_4),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_86),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_86),
.B(n_4),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_94),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_116),
.B1(n_118),
.B2(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_112),
.B1(n_121),
.B2(n_135),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_157),
.B1(n_142),
.B2(n_159),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_126),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_178),
.C(n_138),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_180),
.B1(n_149),
.B2(n_152),
.Y(n_189)
);

AOI21x1_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_126),
.B(n_127),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_171),
.B(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_133),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_137),
.C(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_186),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_144),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_99),
.B1(n_80),
.B2(n_66),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_99),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_99),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_80),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_156),
.A3(n_155),
.B1(n_145),
.B2(n_141),
.C(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_159),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_193),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_168),
.B1(n_176),
.B2(n_6),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_138),
.C(n_153),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_185),
.C(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_150),
.C(n_160),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_154),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_202),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_147),
.B1(n_161),
.B2(n_71),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_147),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_182),
.C(n_169),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_9),
.C(n_11),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_175),
.B(n_171),
.C(n_167),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_217),
.B1(n_195),
.B2(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_168),
.B(n_176),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_5),
.B(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_188),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_192),
.B1(n_203),
.B2(n_198),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_221),
.A2(n_227),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_190),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_225),
.B(n_227),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_7),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_228),
.B(n_11),
.Y(n_233)
);

OAI221xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_217),
.B1(n_204),
.B2(n_210),
.C(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_226),
.B1(n_15),
.B2(n_12),
.Y(n_239)
);

NAND4xp25_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_209),
.C(n_13),
.D(n_14),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_223),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_206),
.C(n_233),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_236),
.C(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_239),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_206),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_242),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_246),
.B(n_240),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_12),
.C(n_15),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_252),
.B(n_248),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_15),
.Y(n_254)
);


endmodule