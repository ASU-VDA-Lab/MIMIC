module real_aes_8270_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_1), .A2(n_151), .B(n_156), .C(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_2), .A2(n_146), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g462 ( .A(n_3), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_4), .B(n_170), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_5), .A2(n_16), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_5), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_6), .A2(n_146), .B(n_480), .Y(n_479) );
AND2x6_ASAP7_75t_L g151 ( .A(n_7), .B(n_152), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_8), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_8), .Y(n_724) );
INVx1_ASAP7_75t_L g180 ( .A(n_9), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_10), .B(n_45), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_11), .A2(n_258), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_12), .B(n_161), .Y(n_197) );
INVx1_ASAP7_75t_L g484 ( .A(n_13), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_14), .B(n_160), .Y(n_532) );
INVx1_ASAP7_75t_L g144 ( .A(n_15), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_16), .Y(n_729) );
INVx1_ASAP7_75t_L g544 ( .A(n_17), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_18), .A2(n_181), .B(n_206), .C(n_208), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_19), .B(n_170), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_473), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_21), .B(n_146), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_22), .B(n_266), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_23), .A2(n_160), .B(n_162), .C(n_166), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_24), .A2(n_49), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_24), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_24), .B(n_170), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_25), .B(n_161), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_26), .A2(n_164), .B(n_208), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_27), .B(n_161), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_28), .Y(n_226) );
INVx1_ASAP7_75t_L g240 ( .A(n_29), .Y(n_240) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_30), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_31), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_32), .B(n_161), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_33), .A2(n_448), .B1(n_722), .B2(n_723), .C1(n_732), .C2(n_733), .Y(n_447) );
INVx1_ASAP7_75t_L g263 ( .A(n_34), .Y(n_263) );
INVx1_ASAP7_75t_L g497 ( .A(n_35), .Y(n_497) );
INVx2_ASAP7_75t_L g149 ( .A(n_36), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_37), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_38), .A2(n_160), .B(n_219), .C(n_221), .Y(n_218) );
INVxp67_ASAP7_75t_L g264 ( .A(n_39), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_40), .A2(n_105), .B1(n_116), .B2(n_736), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g217 ( .A(n_41), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_42), .A2(n_156), .B(n_239), .C(n_245), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_43), .A2(n_151), .B(n_156), .C(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_44), .A2(n_93), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_44), .Y(n_130) );
INVx1_ASAP7_75t_L g496 ( .A(n_46), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_47), .A2(n_178), .B(n_179), .C(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_48), .B(n_161), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_49), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_50), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_51), .Y(n_260) );
INVx1_ASAP7_75t_L g154 ( .A(n_52), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_53), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_54), .B(n_146), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_55), .A2(n_156), .B1(n_166), .B2(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_56), .B(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_57), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_58), .Y(n_459) );
CKINVDCx14_ASAP7_75t_R g176 ( .A(n_59), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_60), .A2(n_178), .B(n_221), .C(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_61), .Y(n_525) );
INVx1_ASAP7_75t_L g481 ( .A(n_62), .Y(n_481) );
INVx1_ASAP7_75t_L g152 ( .A(n_63), .Y(n_152) );
INVx1_ASAP7_75t_L g143 ( .A(n_64), .Y(n_143) );
INVx1_ASAP7_75t_SL g220 ( .A(n_65), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_67), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g229 ( .A(n_68), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_SL g472 ( .A1(n_69), .A2(n_221), .B(n_473), .C(n_474), .Y(n_472) );
INVxp67_ASAP7_75t_L g475 ( .A(n_70), .Y(n_475) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_72), .A2(n_146), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_73), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_74), .A2(n_146), .B(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_75), .Y(n_500) );
INVx1_ASAP7_75t_L g519 ( .A(n_76), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_77), .A2(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g204 ( .A(n_78), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_79), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_80), .A2(n_151), .B(n_156), .C(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_81), .A2(n_146), .B(n_153), .Y(n_145) );
INVx1_ASAP7_75t_L g207 ( .A(n_82), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_83), .B(n_241), .Y(n_513) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx1_ASAP7_75t_L g194 ( .A(n_85), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_86), .B(n_473), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_87), .A2(n_151), .B(n_156), .C(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
OR2x2_ASAP7_75t_L g443 ( .A(n_88), .B(n_112), .Y(n_443) );
OR2x2_ASAP7_75t_L g721 ( .A(n_88), .B(n_113), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_89), .A2(n_156), .B(n_228), .C(n_231), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_90), .A2(n_727), .B1(n_728), .B2(n_731), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_90), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_91), .B(n_173), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_92), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_93), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_94), .A2(n_151), .B(n_156), .C(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_95), .Y(n_536) );
INVx1_ASAP7_75t_L g471 ( .A(n_96), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_97), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_98), .B(n_241), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_99), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_100), .B(n_139), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_101), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g163 ( .A(n_102), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_103), .A2(n_146), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g737 ( .A(n_106), .Y(n_737) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g734 ( .A(n_110), .Y(n_734) );
NOR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g449 ( .A(n_111), .B(n_113), .Y(n_449) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AO21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_446), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g735 ( .A(n_119), .Y(n_735) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_441), .B(n_444), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B1(n_439), .B2(n_440), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_124), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_127), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B1(n_437), .B2(n_438), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_128), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_131), .A2(n_449), .B1(n_450), .B2(n_719), .Y(n_448) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g438 ( .A(n_132), .Y(n_438) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_363), .Y(n_132) );
NOR4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_305), .C(n_335), .D(n_345), .Y(n_133) );
OAI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_210), .B(n_268), .C(n_295), .Y(n_134) );
OAI222xp33_ASAP7_75t_L g390 ( .A1(n_135), .A2(n_310), .B1(n_391), .B2(n_392), .C1(n_393), .C2(n_394), .Y(n_390) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_185), .Y(n_135) );
AOI33xp33_ASAP7_75t_L g316 ( .A1(n_136), .A2(n_303), .A3(n_304), .B1(n_317), .B2(n_322), .B3(n_324), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_136), .A2(n_374), .B(n_376), .C(n_378), .Y(n_373) );
OR2x2_ASAP7_75t_L g389 ( .A(n_136), .B(n_375), .Y(n_389) );
INVx1_ASAP7_75t_L g422 ( .A(n_136), .Y(n_422) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_172), .Y(n_136) );
INVx2_ASAP7_75t_L g299 ( .A(n_137), .Y(n_299) );
AND2x2_ASAP7_75t_L g315 ( .A(n_137), .B(n_201), .Y(n_315) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_137), .Y(n_350) );
AND2x2_ASAP7_75t_L g379 ( .A(n_137), .B(n_172), .Y(n_379) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_145), .B(n_169), .Y(n_137) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_138), .A2(n_202), .B(n_209), .Y(n_201) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_138), .A2(n_215), .B(n_223), .Y(n_214) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx4_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_139), .A2(n_469), .B(n_476), .Y(n_468) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g256 ( .A(n_140), .Y(n_256) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_141), .B(n_142), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx2_ASAP7_75t_L g258 ( .A(n_146), .Y(n_258) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_147), .B(n_151), .Y(n_191) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g244 ( .A(n_148), .Y(n_244) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx1_ASAP7_75t_L g167 ( .A(n_149), .Y(n_167) );
INVx1_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
INVx3_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_L g473 ( .A(n_150), .Y(n_473) );
INVx4_ASAP7_75t_SL g168 ( .A(n_151), .Y(n_168) );
BUFx3_ASAP7_75t_L g245 ( .A(n_151), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g153 ( .A1(n_154), .A2(n_155), .B(n_159), .C(n_168), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_155), .A2(n_168), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_155), .A2(n_168), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_155), .A2(n_168), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_155), .A2(n_168), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_155), .A2(n_168), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_155), .A2(n_168), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_155), .A2(n_168), .B(n_541), .C(n_542), .Y(n_540) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_157), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_160), .B(n_220), .Y(n_219) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_164), .B(n_207), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_164), .A2(n_241), .B1(n_263), .B2(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_164), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_165), .A2(n_196), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g464 ( .A(n_166), .Y(n_464) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_168), .A2(n_191), .B1(n_494), .B2(n_498), .Y(n_493) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_170), .A2(n_479), .B(n_485), .Y(n_478) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_171), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_171), .A2(n_225), .B(n_232), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_171), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g515 ( .A(n_171), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g279 ( .A(n_172), .Y(n_279) );
BUFx3_ASAP7_75t_L g287 ( .A(n_172), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_172), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_172), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_172), .B(n_186), .Y(n_327) );
AND2x2_ASAP7_75t_L g396 ( .A(n_172), .B(n_330), .Y(n_396) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_184), .Y(n_172) );
INVx1_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVx2_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_173), .A2(n_191), .B(n_237), .C(n_238), .Y(n_236) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_173), .A2(n_539), .B(n_545), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx5_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_181), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_181), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
INVx2_ASAP7_75t_SL g290 ( .A(n_185), .Y(n_290) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_201), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_186), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g332 ( .A(n_186), .Y(n_332) );
AND2x2_ASAP7_75t_L g343 ( .A(n_186), .B(n_299), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_186), .B(n_328), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_186), .B(n_330), .Y(n_375) );
AND2x2_ASAP7_75t_L g434 ( .A(n_186), .B(n_379), .Y(n_434) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g304 ( .A(n_187), .B(n_201), .Y(n_304) );
AND2x2_ASAP7_75t_L g314 ( .A(n_187), .B(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g336 ( .A(n_187), .Y(n_336) );
AND3x2_ASAP7_75t_L g395 ( .A(n_187), .B(n_396), .C(n_397), .Y(n_395) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_199), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_188), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_188), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_188), .B(n_536), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_191), .A2(n_226), .B(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_191), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_191), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_197), .C(n_198), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_198), .B(n_229), .C(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_198), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_198), .A2(n_522), .B(n_523), .Y(n_521) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_201), .Y(n_286) );
INVx1_ASAP7_75t_SL g330 ( .A(n_201), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_201), .B(n_279), .C(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_248), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_211), .A2(n_314), .B(n_366), .C(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_213), .B(n_235), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_213), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g382 ( .A(n_213), .Y(n_382) );
AND2x2_ASAP7_75t_L g403 ( .A(n_213), .B(n_250), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_213), .B(n_312), .Y(n_431) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AND2x2_ASAP7_75t_L g276 ( .A(n_214), .B(n_267), .Y(n_276) );
INVx2_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
AND2x2_ASAP7_75t_L g303 ( .A(n_214), .B(n_250), .Y(n_303) );
AND2x2_ASAP7_75t_L g353 ( .A(n_214), .B(n_235), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_214), .Y(n_357) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_222), .Y(n_533) );
INVx2_ASAP7_75t_SL g267 ( .A(n_224), .Y(n_267) );
BUFx2_ASAP7_75t_L g293 ( .A(n_224), .Y(n_293) );
AND2x2_ASAP7_75t_L g420 ( .A(n_224), .B(n_235), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_234), .A2(n_528), .B(n_535), .Y(n_527) );
INVx3_ASAP7_75t_SL g250 ( .A(n_235), .Y(n_250) );
AND2x2_ASAP7_75t_L g275 ( .A(n_235), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g282 ( .A(n_235), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g312 ( .A(n_235), .B(n_272), .Y(n_312) );
OR2x2_ASAP7_75t_L g321 ( .A(n_235), .B(n_267), .Y(n_321) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
AND2x2_ASAP7_75t_L g344 ( .A(n_235), .B(n_297), .Y(n_344) );
AND2x2_ASAP7_75t_L g372 ( .A(n_235), .B(n_252), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_235), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g410 ( .A(n_235), .B(n_251), .Y(n_410) );
OR2x6_ASAP7_75t_L g235 ( .A(n_236), .B(n_246), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_242), .C(n_243), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_241), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_244), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g334 ( .A(n_250), .B(n_283), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_250), .B(n_276), .Y(n_362) );
AND2x2_ASAP7_75t_L g380 ( .A(n_250), .B(n_297), .Y(n_380) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_267), .Y(n_251) );
AND2x2_ASAP7_75t_L g281 ( .A(n_252), .B(n_267), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_252), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
OR2x2_ASAP7_75t_L g367 ( .A(n_252), .B(n_287), .Y(n_367) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B(n_265), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_254), .A2(n_273), .B(n_274), .Y(n_272) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_254), .A2(n_518), .B(n_524), .Y(n_517) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_255), .A2(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_256), .A2(n_458), .B(n_465), .Y(n_457) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_256), .A2(n_493), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_256), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g273 ( .A(n_257), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_265), .Y(n_274) );
AND2x2_ASAP7_75t_L g302 ( .A(n_267), .B(n_272), .Y(n_302) );
INVx1_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
AND2x2_ASAP7_75t_L g405 ( .A(n_267), .B(n_283), .Y(n_405) );
AOI222xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_277), .B1(n_280), .B2(n_284), .C1(n_288), .C2(n_291), .Y(n_268) );
INVx1_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x2_ASAP7_75t_L g296 ( .A(n_270), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g307 ( .A(n_270), .B(n_276), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_270), .B(n_298), .Y(n_323) );
OAI222xp33_ASAP7_75t_L g345 ( .A1(n_270), .A2(n_346), .B1(n_351), .B2(n_352), .C1(n_360), .C2(n_362), .Y(n_345) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g333 ( .A(n_272), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_272), .B(n_353), .Y(n_393) );
AND2x2_ASAP7_75t_L g404 ( .A(n_272), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_275), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_277), .B(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_279), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g349 ( .A(n_279), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx3_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_282), .A2(n_385), .B(n_388), .C(n_390), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_282), .B(n_319), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_282), .B(n_302), .Y(n_424) );
AND2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_293), .Y(n_297) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_287), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g415 ( .A(n_287), .B(n_315), .Y(n_415) );
INVx1_ASAP7_75t_L g427 ( .A(n_287), .Y(n_427) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_290), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g408 ( .A(n_293), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .B(n_300), .C(n_304), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_296), .A2(n_326), .B1(n_341), .B2(n_344), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_297), .B(n_311), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_297), .B(n_319), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_298), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g361 ( .A(n_298), .Y(n_361) );
AND2x2_ASAP7_75t_L g368 ( .A(n_298), .B(n_348), .Y(n_368) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NOR4xp25_ASAP7_75t_L g306 ( .A(n_303), .B(n_307), .C(n_308), .D(n_311), .Y(n_306) );
INVx1_ASAP7_75t_SL g377 ( .A(n_304), .Y(n_377) );
AND2x2_ASAP7_75t_L g421 ( .A(n_304), .B(n_422), .Y(n_421) );
OAI211xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_313), .B(n_316), .C(n_325), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_312), .B(n_382), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_314), .A2(n_433), .B1(n_434), .B2(n_435), .Y(n_432) );
INVx1_ASAP7_75t_SL g387 ( .A(n_315), .Y(n_387) );
AND2x2_ASAP7_75t_L g426 ( .A(n_315), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_319), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_323), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_324), .B(n_349), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_331), .B(n_333), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g401 ( .A(n_328), .Y(n_401) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g429 ( .A(n_329), .Y(n_429) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B(n_340), .Y(n_335) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_336), .Y(n_348) );
OR2x2_ASAP7_75t_L g386 ( .A(n_336), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_339), .A2(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_343), .A2(n_370), .B1(n_373), .B2(n_380), .C(n_381), .Y(n_369) );
INVx1_ASAP7_75t_SL g413 ( .A(n_344), .Y(n_413) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g360 ( .A(n_348), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g397 ( .A(n_350), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_357), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_356), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_398), .C(n_411), .D(n_423), .Y(n_363) );
NAND3xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_369), .C(n_384), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_367), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_374), .B(n_379), .Y(n_383) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_386), .A2(n_412), .B1(n_413), .B2(n_414), .C(n_416), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_388), .A2(n_403), .B(n_404), .C(n_406), .Y(n_402) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_389), .A2(n_407), .B1(n_409), .B2(n_410), .Y(n_406) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_401), .C(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g417 ( .A(n_410), .Y(n_417) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI221xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .B1(n_428), .B2(n_430), .C(n_432), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_438), .A2(n_449), .B1(n_451), .B2(n_721), .Y(n_732) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_442), .Y(n_445) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_SL g446 ( .A1(n_444), .A2(n_447), .B(n_735), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_635), .Y(n_451) );
NOR5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_558), .C(n_590), .D(n_605), .E(n_622), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_486), .B(n_505), .C(n_546), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_467), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_455), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_455), .B(n_610), .Y(n_673) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_456), .B(n_502), .Y(n_559) );
AND2x2_ASAP7_75t_L g600 ( .A(n_456), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_456), .B(n_569), .Y(n_604) );
OR2x2_ASAP7_75t_L g641 ( .A(n_456), .B(n_492), .Y(n_641) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g491 ( .A(n_457), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
OR2x2_ASAP7_75t_L g712 ( .A(n_457), .B(n_552), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_467), .A2(n_615), .B1(n_616), .B2(n_619), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_467), .B(n_549), .Y(n_698) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
AND2x2_ASAP7_75t_L g504 ( .A(n_468), .B(n_492), .Y(n_504) );
AND2x2_ASAP7_75t_L g551 ( .A(n_468), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
INVx3_ASAP7_75t_L g569 ( .A(n_468), .Y(n_569) );
OR2x2_ASAP7_75t_L g589 ( .A(n_468), .B(n_552), .Y(n_589) );
AND2x2_ASAP7_75t_L g608 ( .A(n_468), .B(n_478), .Y(n_608) );
BUFx2_ASAP7_75t_L g640 ( .A(n_468), .Y(n_640) );
AND2x4_ASAP7_75t_L g555 ( .A(n_477), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g490 ( .A(n_478), .Y(n_490) );
INVx2_ASAP7_75t_L g503 ( .A(n_478), .Y(n_503) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_552), .Y(n_571) );
AND2x2_ASAP7_75t_L g601 ( .A(n_478), .B(n_492), .Y(n_601) );
AND2x2_ASAP7_75t_L g618 ( .A(n_478), .B(n_549), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_478), .B(n_569), .Y(n_658) );
AND2x2_ASAP7_75t_SL g694 ( .A(n_478), .B(n_504), .Y(n_694) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp33_ASAP7_75t_SL g487 ( .A(n_488), .B(n_501), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_489), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_490), .A2(n_504), .B(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_490), .B(n_492), .Y(n_688) );
AND2x2_ASAP7_75t_L g624 ( .A(n_491), .B(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_492), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_501), .B(n_549), .Y(n_717) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_502), .A2(n_660), .B1(n_661), .B2(n_666), .Y(n_659) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g550 ( .A(n_503), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g588 ( .A(n_503), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g625 ( .A(n_503), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_504), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g679 ( .A(n_504), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_526), .Y(n_506) );
INVx4_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
AND2x2_ASAP7_75t_L g643 ( .A(n_507), .B(n_610), .Y(n_643) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
INVx3_ASAP7_75t_L g562 ( .A(n_508), .Y(n_562) );
AND2x2_ASAP7_75t_L g576 ( .A(n_508), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
INVx2_ASAP7_75t_L g594 ( .A(n_508), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_508), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g651 ( .A(n_508), .B(n_646), .Y(n_651) );
AND2x2_ASAP7_75t_L g716 ( .A(n_508), .B(n_686), .Y(n_716) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
AND2x2_ASAP7_75t_L g557 ( .A(n_517), .B(n_538), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_517), .Y(n_577) );
INVx1_ASAP7_75t_L g582 ( .A(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g628 ( .A(n_526), .B(n_576), .Y(n_628) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
INVx2_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
INVx1_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_527), .B(n_577), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_567), .Y(n_610) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
AND2x2_ASAP7_75t_L g646 ( .A(n_538), .B(n_577), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_553), .B(n_557), .Y(n_546) );
INVx1_ASAP7_75t_SL g591 ( .A(n_547), .Y(n_591) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_548), .B(n_555), .Y(n_648) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g597 ( .A(n_549), .B(n_552), .Y(n_597) );
AND2x2_ASAP7_75t_L g626 ( .A(n_549), .B(n_570), .Y(n_626) );
OR2x2_ASAP7_75t_L g629 ( .A(n_549), .B(n_589), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g693 ( .A1(n_550), .A2(n_642), .B1(n_694), .B2(n_695), .C1(n_697), .C2(n_699), .Y(n_693) );
BUFx2_ASAP7_75t_L g607 ( .A(n_552), .Y(n_607) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_597), .Y(n_596) );
INVx3_ASAP7_75t_SL g613 ( .A(n_555), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_555), .B(n_607), .Y(n_667) );
AND2x2_ASAP7_75t_L g602 ( .A(n_557), .B(n_562), .Y(n_602) );
INVx1_ASAP7_75t_L g621 ( .A(n_557), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_560), .B1(n_564), .B2(n_568), .C(n_572), .Y(n_558) );
OR2x2_ASAP7_75t_L g630 ( .A(n_560), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g615 ( .A(n_562), .B(n_585), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_562), .B(n_575), .Y(n_655) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_610), .Y(n_660) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_562), .Y(n_670) );
NAND2x1_ASAP7_75t_SL g681 ( .A(n_562), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g566 ( .A(n_563), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g586 ( .A(n_563), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_563), .B(n_581), .Y(n_612) );
INVx1_ASAP7_75t_L g678 ( .A(n_563), .Y(n_678) );
INVx1_ASAP7_75t_L g653 ( .A(n_564), .Y(n_653) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g665 ( .A(n_565), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_565), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g682 ( .A(n_566), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_566), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g585 ( .A(n_567), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_567), .B(n_577), .Y(n_598) );
INVx1_ASAP7_75t_L g664 ( .A(n_567), .Y(n_664) );
INVx1_ASAP7_75t_L g685 ( .A(n_568), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_578), .B(n_587), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
AND2x2_ASAP7_75t_L g718 ( .A(n_574), .B(n_651), .Y(n_718) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g686 ( .A(n_575), .B(n_646), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g599 ( .A1(n_576), .A2(n_582), .A3(n_600), .B1(n_602), .B2(n_603), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g701 ( .A1(n_576), .A2(n_608), .A3(n_691), .B1(n_702), .B2(n_703), .C1(n_704), .C2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g581 ( .A(n_577), .Y(n_581) );
INVx1_ASAP7_75t_L g691 ( .A(n_577), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_579), .B(n_585), .Y(n_634) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_580), .B(n_646), .Y(n_696) );
INVx1_ASAP7_75t_L g583 ( .A(n_581), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_581), .B(n_610), .Y(n_700) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_589), .B(n_684), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B1(n_595), .B2(n_598), .C(n_599), .Y(n_590) );
OR2x2_ASAP7_75t_L g611 ( .A(n_592), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g620 ( .A(n_592), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g645 ( .A(n_593), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g649 ( .A(n_603), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_611), .B2(n_613), .C(n_614), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_607), .A2(n_638), .B1(n_642), .B2(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_608), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_608), .Y(n_713) );
INVx1_ASAP7_75t_L g707 ( .A(n_610), .Y(n_707) );
INVx1_ASAP7_75t_SL g642 ( .A(n_611), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_613), .B(n_641), .Y(n_703) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_618), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g684 ( .A(n_618), .Y(n_684) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_627), .B1(n_629), .B2(n_630), .C(n_632), .Y(n_622) );
NOR2xp33_ASAP7_75t_SL g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_624), .A2(n_642), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx14_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_629), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_668), .C(n_692), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_644), .C(n_652), .D(n_659), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g715 ( .A(n_640), .Y(n_715) );
INVx3_ASAP7_75t_SL g709 ( .A(n_641), .Y(n_709) );
OR2x2_ASAP7_75t_L g714 ( .A(n_641), .B(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_651), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_646), .B(n_664), .Y(n_705) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_656), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_671), .B(n_674), .C(n_687), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g702 ( .A(n_673), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B1(n_680), .B2(n_683), .C1(n_685), .C2(n_686), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND4xp25_ASAP7_75t_SL g711 ( .A(n_684), .B(n_712), .C(n_713), .D(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_701), .C(n_710), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_710) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
endmodule