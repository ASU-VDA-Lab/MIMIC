module fake_jpeg_24709_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_53),
.B1(n_38),
.B2(n_18),
.Y(n_75)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_76),
.Y(n_98)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_58),
.B1(n_60),
.B2(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_97),
.B1(n_109),
.B2(n_71),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_61),
.B(n_58),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_19),
.B(n_24),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_77),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_48),
.B1(n_49),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_104),
.B1(n_106),
.B2(n_112),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_26),
.B1(n_65),
.B2(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_107),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_19),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_43),
.B1(n_34),
.B2(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_34),
.B1(n_32),
.B2(n_39),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_114),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_19),
.B1(n_57),
.B2(n_24),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_28),
.B1(n_34),
.B2(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_39),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_23),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_111),
.B1(n_99),
.B2(n_103),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_133),
.B(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_23),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_132),
.B1(n_136),
.B2(n_139),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_36),
.C(n_19),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_99),
.C(n_103),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_76),
.B1(n_84),
.B2(n_67),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_107),
.B(n_101),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_28),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_67),
.B1(n_90),
.B2(n_24),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_36),
.Y(n_137)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_110),
.B1(n_113),
.B2(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_110),
.B(n_74),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_148),
.B(n_164),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_25),
.B(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_157),
.B(n_165),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_74),
.B(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_36),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_130),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_160),
.B1(n_118),
.B2(n_136),
.Y(n_168)
);

OAI31xp33_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_25),
.A3(n_27),
.B(n_20),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_116),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_115),
.B1(n_105),
.B2(n_25),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_92),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_132),
.B1(n_116),
.B2(n_121),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_31),
.B1(n_21),
.B2(n_17),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_0),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_20),
.B(n_3),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_176),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_120),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_116),
.A3(n_135),
.B1(n_139),
.B2(n_124),
.C1(n_125),
.C2(n_126),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_184),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_92),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_105),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_116),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_54),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_115),
.B1(n_31),
.B2(n_21),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_31),
.B1(n_21),
.B2(n_17),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_155),
.B1(n_145),
.B2(n_159),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_144),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_212),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_157),
.C(n_148),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_204),
.B(n_207),
.Y(n_225)
);

XOR2x1_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_146),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_197),
.B(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_143),
.C(n_165),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_201),
.C(n_31),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_179),
.C(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_143),
.B1(n_158),
.B2(n_164),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_186),
.C(n_171),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_173),
.B1(n_169),
.B2(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_223),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_169),
.B1(n_189),
.B2(n_171),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.C(n_227),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_141),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_200),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_9),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_201),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_211),
.C(n_193),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_243),
.C(n_248),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_203),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_211),
.C(n_212),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_203),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_249),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_197),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_195),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_226),
.B1(n_218),
.B2(n_195),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_202),
.B1(n_219),
.B2(n_220),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_214),
.B(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_9),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_260),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_238),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_239),
.B1(n_235),
.B2(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_2),
.C(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_17),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_274),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_8),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_282),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_255),
.B(n_253),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_273),
.B(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_7),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_267),
.B1(n_271),
.B2(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_288),
.B(n_289),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_279),
.A2(n_10),
.B(n_12),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_10),
.B(n_12),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_11),
.B(n_13),
.Y(n_291)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_284),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_2),
.B(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_296),
.C(n_292),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_297),
.B(n_4),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_5),
.B(n_2),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_147),
.Y(n_303)
);


endmodule