module real_aes_1673_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g578 ( .A(n_0), .B(n_192), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_1), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g150 ( .A(n_2), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_3), .B(n_540), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g621 ( .A(n_4), .B(n_179), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_5), .B(n_159), .Y(n_183) );
INVx1_ASAP7_75t_L g614 ( .A(n_6), .Y(n_614) );
INVx1_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_9), .Y(n_221) );
AND2x2_ASAP7_75t_L g537 ( .A(n_10), .B(n_236), .Y(n_537) );
INVx2_ASAP7_75t_L g158 ( .A(n_11), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g193 ( .A(n_13), .Y(n_193) );
AOI221x1_ASAP7_75t_L g617 ( .A1(n_14), .A2(n_210), .B1(n_542), .B2(n_618), .C(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_15), .B(n_540), .Y(n_601) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g190 ( .A(n_17), .Y(n_190) );
INVx1_ASAP7_75t_SL g265 ( .A(n_18), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_19), .B(n_170), .Y(n_169) );
AOI33xp33_ASAP7_75t_L g242 ( .A1(n_20), .A2(n_49), .A3(n_147), .B1(n_165), .B2(n_243), .B3(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_21), .A2(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_22), .B(n_192), .Y(n_544) );
AOI221xp5_ASAP7_75t_SL g588 ( .A1(n_23), .A2(n_39), .B1(n_540), .B2(n_542), .C(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g214 ( .A(n_24), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_25), .A2(n_104), .B1(n_120), .B2(n_511), .C(n_514), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_25), .A2(n_126), .B1(n_127), .B2(n_507), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_25), .Y(n_126) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_26), .A2(n_91), .B(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g160 ( .A(n_26), .B(n_91), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_27), .B(n_195), .Y(n_605) );
INVxp67_ASAP7_75t_L g616 ( .A(n_28), .Y(n_616) );
AND2x2_ASAP7_75t_L g563 ( .A(n_29), .B(n_235), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_30), .B(n_203), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_31), .A2(n_542), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_32), .B(n_195), .Y(n_590) );
AND2x2_ASAP7_75t_L g153 ( .A(n_33), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g164 ( .A(n_33), .Y(n_164) );
AND2x2_ASAP7_75t_L g179 ( .A(n_33), .B(n_150), .Y(n_179) );
OR2x6_ASAP7_75t_L g114 ( .A(n_34), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_35), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_36), .B(n_203), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_37), .A2(n_144), .B1(n_156), .B2(n_159), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_38), .B(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_40), .A2(n_81), .B1(n_162), .B2(n_542), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_41), .B(n_170), .Y(n_266) );
AOI22xp5_ASAP7_75t_SL g815 ( .A1(n_42), .A2(n_72), .B1(n_816), .B2(n_817), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_42), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_43), .B(n_192), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_44), .B(n_181), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_45), .B(n_170), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_46), .Y(n_155) );
AND2x2_ASAP7_75t_L g581 ( .A(n_47), .B(n_235), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_48), .B(n_235), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_50), .B(n_170), .Y(n_233) );
INVx1_ASAP7_75t_L g148 ( .A(n_51), .Y(n_148) );
INVx1_ASAP7_75t_L g172 ( .A(n_51), .Y(n_172) );
XOR2x2_ASAP7_75t_L g814 ( .A(n_52), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g234 ( .A(n_53), .B(n_235), .Y(n_234) );
AOI221xp5_ASAP7_75t_L g202 ( .A1(n_54), .A2(n_74), .B1(n_162), .B2(n_203), .C(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_55), .B(n_203), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_56), .B(n_540), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_57), .B(n_156), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g253 ( .A1(n_58), .A2(n_162), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g554 ( .A(n_59), .B(n_235), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_60), .B(n_195), .Y(n_579) );
INVx1_ASAP7_75t_L g186 ( .A(n_61), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_62), .B(n_192), .Y(n_552) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_63), .B(n_236), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_64), .A2(n_542), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g232 ( .A(n_65), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_66), .B(n_195), .Y(n_545) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_67), .B(n_181), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_68), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_69), .A2(n_162), .B(n_231), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_70), .A2(n_89), .B1(n_132), .B2(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_70), .Y(n_133) );
INVx1_ASAP7_75t_L g154 ( .A(n_71), .Y(n_154) );
INVx1_ASAP7_75t_L g174 ( .A(n_71), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_72), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_73), .B(n_203), .Y(n_245) );
AND2x2_ASAP7_75t_L g267 ( .A(n_75), .B(n_210), .Y(n_267) );
INVx1_ASAP7_75t_L g187 ( .A(n_76), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_77), .A2(n_162), .B(n_264), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_78), .A2(n_162), .B(n_168), .C(n_180), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_79), .B(n_540), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_80), .A2(n_84), .B1(n_203), .B2(n_540), .Y(n_568) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_83), .B(n_210), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_85), .A2(n_162), .B1(n_240), .B2(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_86), .B(n_192), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_87), .B(n_192), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_88), .A2(n_130), .B1(n_131), .B2(n_134), .Y(n_129) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_89), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_89), .B(n_137), .C(n_478), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_90), .A2(n_542), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g255 ( .A(n_92), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_93), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_94), .B(n_195), .Y(n_551) );
AND2x2_ASAP7_75t_L g246 ( .A(n_95), .B(n_210), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_96), .A2(n_212), .B(n_213), .C(n_215), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_97), .B(n_540), .Y(n_580) );
INVxp67_ASAP7_75t_L g619 ( .A(n_98), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_99), .B(n_195), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_100), .A2(n_542), .B(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_SL g108 ( .A(n_101), .Y(n_108) );
BUFx2_ASAP7_75t_L g513 ( .A(n_101), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_102), .B(n_170), .Y(n_256) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B(n_118), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx8_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_110), .B(n_510), .Y(n_509) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g124 ( .A(n_111), .Y(n_124) );
BUFx2_ASAP7_75t_L g831 ( .A(n_111), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x6_ASAP7_75t_SL g529 ( .A(n_112), .B(n_114), .Y(n_529) );
OR2x6_ASAP7_75t_SL g813 ( .A(n_112), .B(n_113), .Y(n_813) );
OR2x2_ASAP7_75t_L g825 ( .A(n_112), .B(n_114), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OR2x2_ASAP7_75t_SL g512 ( .A(n_118), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g830 ( .A(n_118), .Y(n_830) );
OAI21xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_508), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
CKINVDCx11_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g507 ( .A(n_127), .Y(n_507) );
XNOR2x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_135), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_132), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_SL g523 ( .A1(n_132), .A2(n_524), .B(n_525), .Y(n_523) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_441), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_364), .Y(n_136) );
INVxp67_ASAP7_75t_L g522 ( .A(n_137), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_311), .C(n_344), .Y(n_137) );
AOI211xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_268), .B(n_277), .C(n_301), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_197), .B(n_247), .Y(n_139) );
OR2x2_ASAP7_75t_L g321 ( .A(n_140), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g476 ( .A(n_140), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_141), .A2(n_367), .B1(n_371), .B2(n_373), .Y(n_366) );
AND2x2_ASAP7_75t_L g403 ( .A(n_141), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_182), .Y(n_141) );
INVx1_ASAP7_75t_L g300 ( .A(n_142), .Y(n_300) );
AND2x4_ASAP7_75t_L g317 ( .A(n_142), .B(n_298), .Y(n_317) );
INVx2_ASAP7_75t_L g339 ( .A(n_142), .Y(n_339) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_142), .Y(n_422) );
AND2x2_ASAP7_75t_L g493 ( .A(n_142), .B(n_250), .Y(n_493) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_161), .Y(n_142) );
NOR3xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_151), .C(n_155), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g203 ( .A(n_146), .B(n_152), .Y(n_203) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
OR2x6_ASAP7_75t_L g177 ( .A(n_147), .B(n_166), .Y(n_177) );
INVxp33_ASAP7_75t_L g243 ( .A(n_147), .Y(n_243) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g167 ( .A(n_148), .B(n_150), .Y(n_167) );
AND2x4_ASAP7_75t_L g195 ( .A(n_148), .B(n_173), .Y(n_195) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g542 ( .A(n_153), .B(n_167), .Y(n_542) );
INVx2_ASAP7_75t_L g166 ( .A(n_154), .Y(n_166) );
AND2x6_ASAP7_75t_L g192 ( .A(n_154), .B(n_171), .Y(n_192) );
INVx4_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_156), .B(n_220), .Y(n_219) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_156), .A2(n_575), .B(n_581), .Y(n_574) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_157), .Y(n_181) );
AND2x4_ASAP7_75t_L g159 ( .A(n_158), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_158), .B(n_160), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_159), .B(n_178), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_159), .A2(n_253), .B(n_257), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_159), .A2(n_539), .B(n_541), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_159), .B(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_159), .B(n_616), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_159), .B(n_619), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_159), .B(n_188), .C(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g222 ( .A(n_162), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_162), .A2(n_203), .B1(n_613), .B2(n_615), .Y(n_612) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
NOR2x1p5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx1_ASAP7_75t_L g244 ( .A(n_165), .Y(n_244) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_175), .B(n_178), .Y(n_168) );
INVx1_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
AND2x4_ASAP7_75t_L g540 ( .A(n_170), .B(n_179), .Y(n_540) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_177), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_SL g204 ( .A1(n_177), .A2(n_178), .B(n_205), .C(n_206), .Y(n_204) );
INVxp67_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_177), .A2(n_178), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_177), .A2(n_178), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_177), .A2(n_178), .B(n_265), .C(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_178), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_178), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_178), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_178), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_178), .A2(n_590), .B(n_591), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_178), .A2(n_604), .B(n_605), .Y(n_603) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_179), .Y(n_215) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_180), .A2(n_238), .B(n_246), .Y(n_237) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_180), .A2(n_238), .B(n_246), .Y(n_282) );
AOI21x1_ASAP7_75t_L g566 ( .A1(n_180), .A2(n_567), .B(n_570), .Y(n_566) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_181), .A2(n_202), .B(n_207), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_181), .A2(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g258 ( .A(n_182), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g287 ( .A(n_182), .Y(n_287) );
INVx3_ASAP7_75t_L g298 ( .A(n_182), .Y(n_298) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_189), .B(n_196), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_188), .B(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_193), .B2(n_194), .Y(n_189) );
INVxp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_197), .A2(n_488), .B1(n_490), .B2(n_492), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_197), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_225), .Y(n_198) );
INVx3_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_199), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_199), .Y(n_309) );
NAND2x1_ASAP7_75t_SL g503 ( .A(n_199), .B(n_270), .Y(n_503) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_208), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g276 ( .A(n_201), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_201), .B(n_282), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_201), .B(n_208), .Y(n_307) );
AND2x4_ASAP7_75t_L g314 ( .A(n_201), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_201), .Y(n_363) );
INVxp67_ASAP7_75t_L g370 ( .A(n_201), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_201), .Y(n_375) );
INVx1_ASAP7_75t_L g224 ( .A(n_203), .Y(n_224) );
INVx1_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_208), .B(n_284), .Y(n_293) );
INVx2_ASAP7_75t_L g361 ( .A(n_208), .Y(n_361) );
INVx1_ASAP7_75t_L g400 ( .A(n_208), .Y(n_400) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_218), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B1(n_216), .B2(n_217), .Y(n_209) );
INVx3_ASAP7_75t_L g217 ( .A(n_210), .Y(n_217) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_228), .B(n_234), .Y(n_227) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_217), .A2(n_228), .B(n_234), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B1(n_223), .B2(n_224), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g330 ( .A(n_225), .B(n_307), .Y(n_330) );
AND2x2_ASAP7_75t_L g398 ( .A(n_225), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g412 ( .A(n_225), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_225), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_237), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_227), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g368 ( .A(n_227), .B(n_361), .Y(n_368) );
AND2x2_ASAP7_75t_L g459 ( .A(n_227), .B(n_281), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_235), .Y(n_260) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_235), .A2(n_588), .B(n_592), .Y(n_587) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g270 ( .A(n_237), .Y(n_270) );
INVx2_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
AND2x2_ASAP7_75t_L g360 ( .A(n_237), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_239), .B(n_245), .Y(n_238) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_258), .Y(n_248) );
AND2x2_ASAP7_75t_L g402 ( .A(n_249), .B(n_403), .Y(n_402) );
OR2x6_ASAP7_75t_L g461 ( .A(n_249), .B(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g291 ( .A(n_250), .Y(n_291) );
AND2x4_ASAP7_75t_L g299 ( .A(n_250), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g334 ( .A(n_250), .B(n_259), .Y(n_334) );
INVx2_ASAP7_75t_L g383 ( .A(n_250), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_250), .B(n_357), .Y(n_432) );
AND2x2_ASAP7_75t_L g469 ( .A(n_250), .B(n_287), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_250), .B(n_352), .Y(n_477) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g310 ( .A(n_258), .B(n_299), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_258), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_258), .B(n_337), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_258), .B(n_350), .Y(n_471) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_259), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
INVx2_ASAP7_75t_L g323 ( .A(n_259), .Y(n_323) );
INVx1_ASAP7_75t_L g356 ( .A(n_259), .Y(n_356) );
INVx1_ASAP7_75t_L g404 ( .A(n_259), .Y(n_404) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_267), .Y(n_259) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_260), .A2(n_548), .B(n_554), .Y(n_547) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_260), .A2(n_557), .B(n_563), .Y(n_556) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_260), .A2(n_557), .B(n_563), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_270), .B(n_273), .Y(n_346) );
OR2x2_ASAP7_75t_L g418 ( .A(n_270), .B(n_419), .Y(n_418) );
AND4x1_ASAP7_75t_SL g464 ( .A(n_270), .B(n_446), .C(n_465), .D(n_466), .Y(n_464) );
OR2x2_ASAP7_75t_L g488 ( .A(n_271), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g325 ( .A(n_274), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_274), .B(n_283), .Y(n_475) );
AND2x2_ASAP7_75t_L g500 ( .A(n_275), .B(n_360), .Y(n_500) );
OAI32xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_285), .A3(n_290), .B1(n_292), .B2(n_295), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g373 ( .A(n_280), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g473 ( .A(n_280), .B(n_427), .Y(n_473) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AND2x2_ASAP7_75t_L g369 ( .A(n_281), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g455 ( .A(n_281), .Y(n_455) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_282), .B(n_284), .Y(n_489) );
INVx3_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_283), .B(n_411), .Y(n_484) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_284), .Y(n_343) );
AND2x2_ASAP7_75t_L g362 ( .A(n_284), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g496 ( .A(n_286), .Y(n_496) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g336 ( .A(n_287), .Y(n_336) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_287), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_290), .B(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g328 ( .A(n_291), .B(n_296), .Y(n_328) );
AND2x4_ASAP7_75t_L g350 ( .A(n_291), .B(n_300), .Y(n_350) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_291), .B(n_422), .Y(n_421) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_291), .B(n_372), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_292), .A2(n_415), .B1(n_418), .B2(n_420), .Y(n_414) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_SL g434 ( .A(n_293), .Y(n_434) );
INVx2_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_297), .B(n_303), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_297), .A2(n_433), .B1(n_436), .B2(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g357 ( .A(n_298), .Y(n_357) );
AND2x2_ASAP7_75t_L g380 ( .A(n_298), .B(n_339), .Y(n_380) );
INVx2_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
OAI21xp5_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_304), .B(n_308), .Y(n_301) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_305), .A2(n_377), .B1(n_381), .B2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_306), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_306), .B(n_374), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_306), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_327), .C(n_331), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B1(n_321), .B2(n_324), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g341 ( .A(n_314), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g381 ( .A(n_314), .B(n_368), .Y(n_381) );
AND2x2_ASAP7_75t_L g433 ( .A(n_314), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g450 ( .A(n_314), .B(n_400), .Y(n_450) );
AND2x2_ASAP7_75t_L g505 ( .A(n_314), .B(n_399), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx4_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g382 ( .A(n_317), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
AND2x2_ASAP7_75t_L g396 ( .A(n_320), .B(n_380), .Y(n_396) );
INVx1_ASAP7_75t_L g431 ( .A(n_322), .Y(n_431) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_325), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_326), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_340), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_333), .B(n_372), .Y(n_481) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AOI21xp33_ASAP7_75t_SL g344 ( .A1(n_336), .A2(n_345), .B(n_347), .Y(n_344) );
AND2x2_ASAP7_75t_L g491 ( .A(n_336), .B(n_350), .Y(n_491) );
AND2x4_ASAP7_75t_L g354 ( .A(n_337), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g388 ( .A(n_337), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_337), .B(n_404), .Y(n_470) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_353), .B(n_358), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_350), .B(n_355), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_351), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g413 ( .A(n_351), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_351), .Y(n_417) );
AND2x2_ASAP7_75t_L g501 ( .A(n_351), .B(n_469), .Y(n_501) );
AND2x2_ASAP7_75t_L g504 ( .A(n_351), .B(n_421), .Y(n_504) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_SL g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_356), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g483 ( .A(n_360), .Y(n_483) );
AND2x2_ASAP7_75t_L g374 ( .A(n_361), .B(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_364), .B(n_442), .Y(n_519) );
INVxp67_ASAP7_75t_L g521 ( .A(n_364), .Y(n_521) );
NAND4xp75_ASAP7_75t_L g364 ( .A(n_365), .B(n_384), .C(n_405), .D(n_423), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_376), .Y(n_365) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_368), .B(n_455), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_369), .B(n_434), .Y(n_440) );
NAND2xp5_ASAP7_75t_R g456 ( .A(n_372), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g506 ( .A(n_372), .Y(n_506) );
INVx2_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
BUFx3_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g462 ( .A(n_380), .Y(n_462) );
AND2x2_ASAP7_75t_L g416 ( .A(n_382), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g438 ( .A(n_383), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B(n_391), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_387), .B(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_388), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_390), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B1(n_397), .B2(n_401), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_399), .A2(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g458 ( .A(n_400), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_401), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g436 ( .A(n_404), .B(n_437), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .B(n_414), .Y(n_405) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g453 ( .A(n_410), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
INVx2_ASAP7_75t_SL g457 ( .A(n_421), .Y(n_457) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_435), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_428), .B1(n_430), .B2(n_433), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_478), .Y(n_441) );
INVxp67_ASAP7_75t_L g525 ( .A(n_442), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .C(n_463), .Y(n_442) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_448), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_456), .B1(n_458), .B2(n_460), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .C(n_474), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B(n_472), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_497), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_487), .C(n_494), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_485), .B2(n_486), .Y(n_480) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_488), .B(n_493), .C(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B1(n_502), .B2(n_504), .C1(n_505), .C2(n_506), .Y(n_497) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g829 ( .A(n_513), .B(n_830), .Y(n_829) );
AOI31xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_818), .A3(n_821), .B(n_826), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_814), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_526), .B1(n_530), .B2(n_811), .Y(n_516) );
AO22x2_ASAP7_75t_L g820 ( .A1(n_517), .A2(n_527), .B1(n_530), .B2(n_812), .Y(n_820) );
AOI211x1_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .C(n_523), .Y(n_517) );
INVx4_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_741), .Y(n_531) );
NOR4xp25_ASAP7_75t_SL g532 ( .A(n_533), .B(n_634), .C(n_678), .D(n_705), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_597), .B1(n_607), .B2(n_622), .C(n_624), .Y(n_533) );
AOI32xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_564), .A3(n_571), .B1(n_582), .B2(n_593), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_535), .B(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_535), .A2(n_747), .B1(n_805), .B2(n_808), .Y(n_804) );
AND2x4_ASAP7_75t_SL g535 ( .A(n_536), .B(n_546), .Y(n_535) );
INVx5_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
OR2x2_ASAP7_75t_L g623 ( .A(n_536), .B(n_595), .Y(n_623) );
AND2x4_ASAP7_75t_L g625 ( .A(n_536), .B(n_556), .Y(n_625) );
INVx2_ASAP7_75t_L g640 ( .A(n_536), .Y(n_640) );
OR2x2_ASAP7_75t_L g652 ( .A(n_536), .B(n_565), .Y(n_652) );
AND2x2_ASAP7_75t_L g659 ( .A(n_536), .B(n_555), .Y(n_659) );
AND2x2_ASAP7_75t_SL g701 ( .A(n_536), .B(n_584), .Y(n_701) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_536), .Y(n_758) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx3_ASAP7_75t_SL g653 ( .A(n_546), .Y(n_653) );
AND2x2_ASAP7_75t_L g672 ( .A(n_546), .B(n_596), .Y(n_672) );
AOI32xp33_ASAP7_75t_L g787 ( .A1(n_546), .A2(n_658), .A3(n_688), .B1(n_718), .B2(n_753), .Y(n_787) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_555), .Y(n_546) );
AND2x2_ASAP7_75t_L g627 ( .A(n_547), .B(n_565), .Y(n_627) );
OR2x2_ASAP7_75t_L g643 ( .A(n_547), .B(n_556), .Y(n_643) );
INVx1_ASAP7_75t_L g666 ( .A(n_547), .Y(n_666) );
INVx2_ASAP7_75t_L g682 ( .A(n_547), .Y(n_682) );
AND2x2_ASAP7_75t_L g719 ( .A(n_547), .B(n_584), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_547), .B(n_556), .Y(n_738) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_547), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g774 ( .A(n_556), .B(n_565), .Y(n_774) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_556), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
OR2x2_ASAP7_75t_L g622 ( .A(n_564), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g628 ( .A(n_564), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g641 ( .A(n_564), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g803 ( .A(n_564), .B(n_672), .Y(n_803) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g732 ( .A(n_565), .B(n_682), .Y(n_732) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_566), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_571), .B(n_699), .Y(n_801) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_572), .B(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g586 ( .A(n_573), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
AND2x2_ASAP7_75t_L g632 ( .A(n_573), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_573), .B(n_610), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_573), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g690 ( .A(n_573), .Y(n_690) );
OR2x2_ASAP7_75t_L g709 ( .A(n_573), .B(n_636), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_573), .Y(n_716) );
NOR2xp33_ASAP7_75t_R g768 ( .A(n_573), .B(n_599), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_573), .B(n_611), .Y(n_772) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
AOI32xp33_ASAP7_75t_L g795 ( .A1(n_582), .A2(n_631), .A3(n_796), .B1(n_797), .B2(n_798), .Y(n_795) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
AND2x4_ASAP7_75t_L g681 ( .A(n_584), .B(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_584), .B(n_653), .Y(n_710) );
OR2x2_ASAP7_75t_L g764 ( .A(n_584), .B(n_765), .Y(n_764) );
OR2x2_ASAP7_75t_L g722 ( .A(n_585), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g780 ( .A(n_585), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_586), .B(n_599), .Y(n_746) );
AND2x2_ASAP7_75t_L g783 ( .A(n_586), .B(n_749), .Y(n_783) );
INVx2_ASAP7_75t_L g633 ( .A(n_587), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_587), .B(n_599), .Y(n_656) );
INVx1_ASAP7_75t_L g687 ( .A(n_587), .Y(n_687) );
OR2x2_ASAP7_75t_L g713 ( .A(n_587), .B(n_599), .Y(n_713) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_587), .Y(n_765) );
BUFx3_ASAP7_75t_L g794 ( .A(n_587), .Y(n_794) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g663 ( .A(n_594), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_594), .B(n_681), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_594), .B(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_595), .B(n_666), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_595), .A2(n_662), .B(n_680), .Y(n_695) );
OAI32xp33_ASAP7_75t_L g717 ( .A1(n_596), .A2(n_718), .A3(n_720), .B1(n_722), .B2(n_724), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_596), .B(n_681), .Y(n_790) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g723 ( .A(n_598), .Y(n_723) );
NOR2x1p5_ASAP7_75t_L g793 ( .A(n_598), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g609 ( .A(n_599), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_SL g631 ( .A(n_599), .B(n_611), .Y(n_631) );
OR2x2_ASAP7_75t_L g635 ( .A(n_599), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g670 ( .A(n_599), .Y(n_670) );
AND2x2_ASAP7_75t_L g688 ( .A(n_599), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g699 ( .A(n_599), .B(n_611), .Y(n_699) );
OR2x2_ASAP7_75t_L g761 ( .A(n_599), .B(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g778 ( .A(n_599), .B(n_709), .Y(n_778) );
INVx1_ASAP7_75t_L g810 ( .A(n_599), .Y(n_810) );
OR2x6_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_608), .B(n_687), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_609), .B(n_721), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g725 ( .A1(n_609), .A2(n_726), .B1(n_731), .B2(n_733), .C1(n_736), .C2(n_739), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_609), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g753 ( .A(n_609), .B(n_632), .Y(n_753) );
AND2x2_ASAP7_75t_L g715 ( .A(n_610), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g730 ( .A(n_610), .B(n_635), .Y(n_730) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_611), .B(n_636), .Y(n_668) );
AND2x4_ASAP7_75t_L g689 ( .A(n_611), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g749 ( .A(n_611), .B(n_670), .Y(n_749) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
INVx1_ASAP7_75t_SL g629 ( .A(n_623), .Y(n_629) );
NAND2xp33_ASAP7_75t_SL g798 ( .A(n_623), .B(n_653), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_628), .C(n_630), .Y(n_624) );
INVx2_ASAP7_75t_SL g675 ( .A(n_625), .Y(n_675) );
AND2x2_ASAP7_75t_L g679 ( .A(n_626), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_627), .B(n_675), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_627), .A2(n_665), .B(n_701), .C(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g777 ( .A(n_627), .B(n_758), .Y(n_777) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x4_ASAP7_75t_L g676 ( .A(n_631), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g781 ( .A(n_631), .Y(n_781) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B(n_644), .C(n_671), .Y(n_634) );
INVx2_ASAP7_75t_L g646 ( .A(n_635), .Y(n_646) );
OR2x2_ASAP7_75t_L g693 ( .A(n_635), .B(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_636), .Y(n_677) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_639), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g731 ( .A(n_639), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_639), .B(n_719), .Y(n_785) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_641), .A2(n_744), .B1(n_745), .B2(n_747), .C1(n_750), .C2(n_753), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_642), .A2(n_707), .B1(n_710), .B2(n_711), .C(n_717), .Y(n_706) );
AND2x2_ASAP7_75t_L g744 ( .A(n_642), .B(n_701), .Y(n_744) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_643), .B(n_658), .Y(n_657) );
AOI221x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_654), .B2(n_657), .C(n_660), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g797 ( .A(n_647), .B(n_735), .Y(n_797) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g655 ( .A(n_648), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g763 ( .A1(n_653), .A2(n_694), .A3(n_764), .B1(n_766), .B2(n_770), .Y(n_763) );
OAI21xp33_ASAP7_75t_SL g782 ( .A1(n_654), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_667), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
OR2x2_ASAP7_75t_L g664 ( .A(n_662), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g737 ( .A(n_662), .B(n_738), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_666), .A2(n_692), .B1(n_695), .B2(n_696), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g767 ( .A(n_666), .Y(n_767) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_666), .Y(n_773) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_675), .B(n_740), .Y(n_739) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_683), .B(n_691), .Y(n_678) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_682), .Y(n_752) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_685), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g704 ( .A(n_687), .Y(n_704) );
INVx1_ASAP7_75t_L g694 ( .A(n_689), .Y(n_694) );
AND2x2_ASAP7_75t_SL g703 ( .A(n_689), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_689), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_689), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g708 ( .A(n_699), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_704), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_725), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g721 ( .A(n_709), .Y(n_721) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_SL g735 ( .A(n_713), .Y(n_735) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_715), .B(n_793), .Y(n_792) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_716), .Y(n_729) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_727), .B(n_730), .Y(n_726) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g740 ( .A(n_732), .Y(n_740) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g759 ( .A(n_738), .Y(n_759) );
NOR4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_775), .C(n_786), .D(n_799), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_754), .Y(n_742) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_744), .A2(n_755), .B(n_760), .C(n_763), .Y(n_754) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_759), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g766 ( .A1(n_757), .A2(n_767), .B(n_768), .C(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_773), .B(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_774), .B(n_806), .Y(n_805) );
OAI221xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_778), .B1(n_779), .B2(n_780), .C(n_782), .Y(n_775) );
INVx1_ASAP7_75t_SL g779 ( .A(n_777), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND3xp33_ASAP7_75t_SL g786 ( .A(n_787), .B(n_788), .C(n_795), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI21xp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B(n_804), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVxp33_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
CKINVDCx11_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_814), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_831), .Y(n_827) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
endmodule