module real_aes_2575_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_0), .B(n_177), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_1), .A2(n_67), .B1(n_127), .B2(n_128), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_2), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_2), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_2), .A2(n_185), .B(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_3), .A2(n_82), .B1(n_83), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_3), .Y(n_503) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_4), .A2(n_57), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_5), .B(n_192), .Y(n_255) );
INVx1_ASAP7_75t_L g161 ( .A(n_6), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g145 ( .A1(n_7), .A2(n_41), .B1(n_146), .B2(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_7), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_8), .B(n_192), .Y(n_230) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_9), .A2(n_27), .B1(n_90), .B2(n_91), .Y(n_89) );
NAND2xp33_ASAP7_75t_L g193 ( .A(n_10), .B(n_194), .Y(n_193) );
AO222x2_ASAP7_75t_SL g86 ( .A1(n_11), .A2(n_22), .B1(n_50), .B2(n_87), .C1(n_103), .C2(n_106), .Y(n_86) );
INVx2_ASAP7_75t_L g174 ( .A(n_12), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_13), .A2(n_52), .B1(n_139), .B2(n_140), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_14), .A2(n_48), .B1(n_112), .B2(n_115), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_15), .A2(n_142), .B1(n_148), .B2(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g148 ( .A(n_15), .Y(n_148) );
AOI221x1_ASAP7_75t_L g271 ( .A1(n_16), .A2(n_23), .B1(n_177), .B2(n_185), .C(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_17), .B(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_18), .A2(n_172), .B(n_175), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_19), .B(n_210), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_20), .B(n_192), .Y(n_219) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_21), .A2(n_177), .B(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_24), .A2(n_36), .B1(n_118), .B2(n_121), .Y(n_117) );
NAND2x1_ASAP7_75t_L g241 ( .A(n_25), .B(n_192), .Y(n_241) );
NAND2x1_ASAP7_75t_L g229 ( .A(n_26), .B(n_194), .Y(n_229) );
OAI221xp5_ASAP7_75t_L g153 ( .A1(n_27), .A2(n_57), .B1(n_62), .B2(n_154), .C(n_156), .Y(n_153) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_28), .A2(n_68), .B(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g197 ( .A(n_28), .B(n_68), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_29), .B(n_194), .Y(n_209) );
INVx3_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_31), .B(n_192), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_32), .A2(n_46), .B1(n_131), .B2(n_132), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_33), .B(n_194), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_34), .A2(n_185), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_SL g98 ( .A(n_35), .Y(n_98) );
INVx1_ASAP7_75t_L g163 ( .A(n_37), .Y(n_163) );
AND2x2_ASAP7_75t_L g183 ( .A(n_37), .B(n_161), .Y(n_183) );
AND2x2_ASAP7_75t_L g186 ( .A(n_37), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_38), .B(n_177), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_39), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_40), .B(n_194), .Y(n_262) );
INVx1_ASAP7_75t_L g146 ( .A(n_41), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_42), .A2(n_185), .B(n_228), .Y(n_227) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_43), .A2(n_62), .B1(n_90), .B2(n_102), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_44), .A2(n_63), .B1(n_136), .B2(n_137), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_45), .B(n_194), .Y(n_242) );
INVx1_ASAP7_75t_L g180 ( .A(n_47), .Y(n_180) );
INVx1_ASAP7_75t_L g189 ( .A(n_47), .Y(n_189) );
INVx1_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_51), .B(n_192), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_53), .A2(n_185), .B(n_240), .Y(n_239) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_54), .A2(n_185), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_55), .B(n_177), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_56), .B(n_177), .Y(n_231) );
INVxp33_ASAP7_75t_L g158 ( .A(n_57), .Y(n_158) );
INVx1_ASAP7_75t_L g81 ( .A(n_58), .Y(n_81) );
AND2x2_ASAP7_75t_L g265 ( .A(n_59), .B(n_211), .Y(n_265) );
INVx1_ASAP7_75t_L g182 ( .A(n_60), .Y(n_182) );
INVx1_ASAP7_75t_L g187 ( .A(n_60), .Y(n_187) );
AND2x2_ASAP7_75t_L g233 ( .A(n_61), .B(n_202), .Y(n_233) );
INVxp67_ASAP7_75t_L g157 ( .A(n_62), .Y(n_157) );
AND2x2_ASAP7_75t_L g201 ( .A(n_64), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_65), .B(n_177), .Y(n_221) );
AND2x2_ASAP7_75t_L g251 ( .A(n_66), .B(n_196), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_69), .B(n_194), .Y(n_220) );
INVx1_ASAP7_75t_L g512 ( .A(n_69), .Y(n_512) );
AND2x2_ASAP7_75t_L g245 ( .A(n_70), .B(n_202), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_71), .B(n_192), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_72), .A2(n_185), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g496 ( .A(n_72), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_73), .B(n_194), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_74), .B(n_192), .Y(n_208) );
BUFx2_ASAP7_75t_SL g155 ( .A(n_75), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_76), .A2(n_185), .B(n_190), .Y(n_184) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_150), .B1(n_164), .B2(n_486), .C(n_493), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_141), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_82), .A2(n_83), .B1(n_495), .B2(n_496), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2x1_ASAP7_75t_L g84 ( .A(n_85), .B(n_124), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_110), .Y(n_85) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g140 ( .A(n_88), .B(n_133), .Y(n_140) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_93), .Y(n_105) );
INVx1_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
INVx1_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
INVx2_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
OAI22x1_ASAP7_75t_L g96 ( .A1(n_90), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_90), .Y(n_97) );
INVx1_ASAP7_75t_L g102 ( .A(n_90), .Y(n_102) );
AND2x4_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g119 ( .A(n_93), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g118 ( .A(n_95), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g131 ( .A(n_95), .B(n_108), .Y(n_131) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_100), .Y(n_95) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_96), .Y(n_104) );
AND2x2_ASAP7_75t_L g107 ( .A(n_96), .B(n_101), .Y(n_107) );
INVx2_ASAP7_75t_L g114 ( .A(n_96), .Y(n_114) );
AND2x4_ASAP7_75t_L g133 ( .A(n_100), .B(n_114), .Y(n_133) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g113 ( .A(n_101), .B(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g129 ( .A(n_101), .Y(n_129) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x4_ASAP7_75t_L g128 ( .A(n_105), .B(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g132 ( .A(n_105), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g115 ( .A(n_107), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g121 ( .A(n_107), .B(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_L g136 ( .A(n_108), .B(n_113), .Y(n_136) );
AND2x2_ASAP7_75t_L g139 ( .A(n_108), .B(n_133), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_117), .Y(n_110) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_113), .B(n_119), .Y(n_127) );
AND2x6_ASAP7_75t_L g137 ( .A(n_119), .B(n_133), .Y(n_137) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_120), .Y(n_123) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_134), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_138), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_142), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
AND3x1_ASAP7_75t_SL g152 ( .A(n_153), .B(n_159), .C(n_162), .Y(n_152) );
INVxp67_ASAP7_75t_L g501 ( .A(n_153), .Y(n_501) );
CKINVDCx8_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_159), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g508 ( .A1(n_159), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g490 ( .A(n_160), .B(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_SL g506 ( .A(n_160), .B(n_162), .Y(n_506) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g188 ( .A(n_161), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_162), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_407), .Y(n_165) );
NOR3xp33_ASAP7_75t_SL g166 ( .A(n_167), .B(n_319), .C(n_359), .Y(n_166) );
OAI221xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_234), .B1(n_283), .B2(n_298), .C(n_301), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_198), .Y(n_169) );
INVx2_ASAP7_75t_L g316 ( .A(n_170), .Y(n_316) );
AND2x2_ASAP7_75t_L g346 ( .A(n_170), .B(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g284 ( .A(n_171), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g291 ( .A(n_171), .B(n_224), .Y(n_291) );
INVx2_ASAP7_75t_L g297 ( .A(n_171), .Y(n_297) );
AND2x2_ASAP7_75t_L g306 ( .A(n_171), .B(n_200), .Y(n_306) );
INVx1_ASAP7_75t_L g322 ( .A(n_171), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_171), .B(n_368), .Y(n_367) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g203 ( .A(n_173), .Y(n_203) );
AND2x4_ASAP7_75t_L g196 ( .A(n_174), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_174), .B(n_197), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_184), .B(n_196), .Y(n_175) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_183), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
AND2x6_ASAP7_75t_L g194 ( .A(n_179), .B(n_187), .Y(n_194) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x4_ASAP7_75t_L g192 ( .A(n_181), .B(n_189), .Y(n_192) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx5_ASAP7_75t_L g195 ( .A(n_183), .Y(n_195) );
AND2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
BUFx3_ASAP7_75t_L g492 ( .A(n_186), .Y(n_492) );
INVx2_ASAP7_75t_L g491 ( .A(n_189), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_195), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_195), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_195), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_195), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_195), .A2(n_254), .B(n_255), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_195), .A2(n_262), .B(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_195), .A2(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g215 ( .A(n_196), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_196), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_199), .B(n_212), .Y(n_198) );
INVx4_ASAP7_75t_L g287 ( .A(n_199), .Y(n_287) );
AND2x2_ASAP7_75t_L g318 ( .A(n_199), .B(n_225), .Y(n_318) );
AND2x2_ASAP7_75t_L g394 ( .A(n_199), .B(n_368), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_199), .B(n_224), .Y(n_436) );
INVx5_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_200), .B(n_224), .Y(n_323) );
AND2x2_ASAP7_75t_L g347 ( .A(n_200), .B(n_225), .Y(n_347) );
BUFx2_ASAP7_75t_L g363 ( .A(n_200), .Y(n_363) );
NOR2x1_ASAP7_75t_SL g466 ( .A(n_200), .B(n_368), .Y(n_466) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_204), .Y(n_200) );
INVx3_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_210), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_210), .Y(n_232) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_210), .A2(n_271), .B(n_275), .Y(n_270) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_210), .A2(n_271), .B(n_275), .Y(n_333) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g343 ( .A(n_212), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_212), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_419), .Y(n_409) );
AND2x2_ASAP7_75t_L g429 ( .A(n_212), .B(n_322), .Y(n_429) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_224), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
INVx1_ASAP7_75t_L g338 ( .A(n_214), .Y(n_338) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_215), .B(n_223), .Y(n_222) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_215), .A2(n_216), .B(n_222), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_224), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_224), .B(n_295), .Y(n_307) );
INVx2_ASAP7_75t_L g349 ( .A(n_224), .Y(n_349) );
AND2x2_ASAP7_75t_L g482 ( .A(n_224), .B(n_297), .Y(n_482) );
INVx4_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_225), .Y(n_339) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_233), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
NOR3xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_266), .C(n_281), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_246), .Y(n_235) );
INVx2_ASAP7_75t_L g396 ( .A(n_236), .Y(n_396) );
AND2x2_ASAP7_75t_L g441 ( .A(n_236), .B(n_318), .Y(n_441) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g386 ( .A(n_237), .Y(n_386) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_237), .B(n_313), .Y(n_401) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B(n_245), .Y(n_237) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_238), .A2(n_244), .B(n_245), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_244), .A2(n_259), .B(n_265), .Y(n_258) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_244), .A2(n_259), .B(n_265), .Y(n_278) );
INVx2_ASAP7_75t_L g355 ( .A(n_246), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_246), .B(n_385), .Y(n_411) );
AND2x4_ASAP7_75t_L g444 ( .A(n_246), .B(n_391), .Y(n_444) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_258), .Y(n_246) );
AND2x2_ASAP7_75t_L g282 ( .A(n_247), .B(n_277), .Y(n_282) );
OR2x2_ASAP7_75t_L g312 ( .A(n_247), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_247), .B(n_333), .Y(n_381) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
OAI21x1_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_252), .B(n_256), .Y(n_249) );
INVx1_ASAP7_75t_L g257 ( .A(n_251), .Y(n_257) );
INVx2_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_260), .B(n_264), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_266), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_276), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_268), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g354 ( .A(n_268), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g439 ( .A(n_268), .Y(n_439) );
BUFx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g418 ( .A(n_269), .B(n_278), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_269), .B(n_288), .Y(n_422) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g391 ( .A(n_270), .Y(n_391) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_270), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_276), .B(n_299), .Y(n_375) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_277), .B(n_300), .Y(n_485) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_280), .Y(n_289) );
AND2x2_ASAP7_75t_L g371 ( .A(n_278), .B(n_333), .Y(n_371) );
AND2x2_ASAP7_75t_L g390 ( .A(n_278), .B(n_279), .Y(n_390) );
BUFx2_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_279), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g288 ( .A(n_280), .Y(n_288) );
INVxp67_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
INVx1_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
AND2x2_ASAP7_75t_L g340 ( .A(n_282), .B(n_311), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_282), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g458 ( .A(n_282), .B(n_459), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B1(n_289), .B2(n_290), .C(n_292), .Y(n_283) );
AND2x2_ASAP7_75t_L g387 ( .A(n_284), .B(n_287), .Y(n_387) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_284), .B(n_347), .Y(n_406) );
AND2x2_ASAP7_75t_L g424 ( .A(n_284), .B(n_349), .Y(n_424) );
AND2x2_ASAP7_75t_L g479 ( .A(n_284), .B(n_318), .Y(n_479) );
INVx1_ASAP7_75t_L g295 ( .A(n_285), .Y(n_295) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_285), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_286), .Y(n_431) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_287), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_287), .B(n_338), .Y(n_413) );
AND2x2_ASAP7_75t_L g380 ( .A(n_288), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g416 ( .A(n_288), .Y(n_416) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_289), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g467 ( .A(n_289), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_289), .B(n_391), .Y(n_477) );
AND2x4_ASAP7_75t_L g393 ( .A(n_290), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g464 ( .A(n_291), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
OR2x2_ASAP7_75t_L g335 ( .A(n_296), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g342 ( .A(n_297), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g373 ( .A(n_297), .B(n_347), .Y(n_373) );
AND2x2_ASAP7_75t_L g447 ( .A(n_297), .B(n_368), .Y(n_447) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g395 ( .A(n_299), .B(n_396), .Y(n_395) );
OAI32xp33_ASAP7_75t_L g460 ( .A1(n_299), .A2(n_461), .A3(n_463), .B1(n_464), .B2(n_467), .Y(n_460) );
AND2x4_ASAP7_75t_L g332 ( .A(n_300), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g430 ( .A(n_300), .B(n_333), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_308), .B2(n_314), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_SL g419 ( .A1(n_303), .A2(n_317), .B(n_420), .C(n_421), .Y(n_419) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g403 ( .A(n_304), .B(n_331), .Y(n_403) );
INVx1_ASAP7_75t_SL g474 ( .A(n_305), .Y(n_474) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x4_ASAP7_75t_L g377 ( .A(n_307), .B(n_316), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_307), .A2(n_456), .B1(n_457), .B2(n_458), .C(n_460), .Y(n_455) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_312), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_315), .A2(n_345), .B1(n_398), .B2(n_399), .Y(n_397) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_316), .A2(n_434), .B(n_442), .C(n_455), .Y(n_433) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g353 ( .A(n_318), .B(n_322), .Y(n_353) );
OAI211xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_324), .B(n_327), .C(n_356), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g350 ( .A(n_322), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g470 ( .A(n_322), .B(n_466), .Y(n_470) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_323), .A2(n_428), .A3(n_430), .B1(n_431), .B2(n_432), .Y(n_427) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_326), .B(n_418), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_334), .B1(n_340), .B2(n_341), .C(n_344), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g484 ( .A(n_331), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_332), .B(n_396), .Y(n_398) );
A2O1A1O1Ixp25_ASAP7_75t_L g469 ( .A1(n_332), .A2(n_401), .B(n_417), .C(n_463), .D(n_470), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g471 ( .A1(n_332), .A2(n_353), .A3(n_463), .B(n_470), .Y(n_471) );
AND2x2_ASAP7_75t_L g385 ( .A(n_333), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_335), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx2_ASAP7_75t_L g462 ( .A(n_337), .Y(n_462) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g457 ( .A(n_338), .B(n_349), .Y(n_457) );
INVx1_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
AND2x2_ASAP7_75t_L g357 ( .A(n_341), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AOI31xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .A3(n_352), .B(n_354), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_347), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g480 ( .A(n_347), .B(n_426), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g425 ( .A(n_349), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g451 ( .A(n_349), .Y(n_451) );
INVxp67_ASAP7_75t_L g420 ( .A(n_350), .Y(n_420) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g358 ( .A(n_354), .Y(n_358) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_376), .C(n_392), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_369), .B1(n_373), .B2(n_374), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g446 ( .A(n_363), .Y(n_446) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_367), .Y(n_426) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_367), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_367), .B(n_436), .Y(n_453) );
NAND2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_387), .B2(n_388), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_390), .B1(n_424), .B2(n_425), .C(n_427), .Y(n_423) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g463 ( .A(n_390), .Y(n_463) );
AND2x2_ASAP7_75t_L g400 ( .A(n_391), .B(n_401), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_SL g448 ( .A1(n_391), .A2(n_449), .B(n_453), .C(n_454), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_397), .C(n_402), .Y(n_392) );
AND2x2_ASAP7_75t_L g443 ( .A(n_396), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
AOI21xp33_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B(n_405), .Y(n_402) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_433), .C(n_468), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_423), .Y(n_408) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
INVxp67_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g440 ( .A(n_430), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_440), .B2(n_441), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_445), .B(n_448), .Y(n_442) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g481 ( .A(n_466), .B(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_472), .B2(n_475), .C(n_478), .Y(n_468) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI31xp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .A3(n_481), .B(n_483), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_491), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_492), .Y(n_511) );
OAI222xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B1(n_502), .B2(n_504), .C1(n_507), .C2(n_512), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
endmodule