module real_jpeg_30347_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_685, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_685;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_666;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_578;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_372;
wire n_219;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_0),
.Y(n_290)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_0),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_60),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_1),
.A2(n_181),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_1),
.A2(n_181),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_1),
.A2(n_181),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_2),
.A2(n_125),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_2),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_2),
.A2(n_329),
.B1(n_470),
.B2(n_474),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_2),
.A2(n_329),
.B1(n_516),
.B2(n_520),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_2),
.A2(n_35),
.B1(n_329),
.B2(n_593),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_3),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_4),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_33),
.B1(n_125),
.B2(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_33),
.B1(n_167),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_5),
.A2(n_33),
.B1(n_416),
.B2(n_420),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_6),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_124),
.B1(n_164),
.B2(n_167),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g249 ( 
.A1(n_6),
.A2(n_124),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_6),
.A2(n_124),
.B1(n_670),
.B2(n_673),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_9),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_10),
.A2(n_59),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_10),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_10),
.A2(n_88),
.B1(n_226),
.B2(n_259),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_10),
.A2(n_259),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_10),
.A2(n_259),
.B1(n_395),
.B2(n_399),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_11),
.A2(n_313),
.B1(n_314),
.B2(n_317),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_11),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_11),
.A2(n_313),
.B1(n_355),
.B2(n_360),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_11),
.A2(n_313),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_11),
.A2(n_313),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_13),
.B(n_40),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_13),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_13),
.B(n_424),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_13),
.A2(n_372),
.B1(n_479),
.B2(n_482),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_13),
.A2(n_287),
.B(n_504),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_14),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_14),
.A2(n_57),
.B1(n_222),
.B2(n_226),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_14),
.A2(n_57),
.B1(n_293),
.B2(n_297),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_14),
.A2(n_57),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_15),
.B(n_661),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_15),
.B(n_660),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_16),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_16),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_17),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_17),
.A2(n_86),
.B1(n_193),
.B2(n_198),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_17),
.A2(n_86),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_18),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_658),
.B(n_680),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_204),
.B(n_656),
.Y(n_20)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_21),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_185),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_22),
.B(n_185),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_171),
.C(n_184),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_24),
.A2(n_179),
.B1(n_184),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_24),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_78),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_25),
.B(n_170),
.C(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_38),
.B1(n_52),
.B2(n_62),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_26),
.Y(n_191)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_32),
.Y(n_183)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g318 ( 
.A(n_37),
.Y(n_318)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_39),
.A2(n_53),
.B1(n_63),
.B2(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_39),
.A2(n_63),
.B1(n_192),
.B2(n_669),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_40),
.B(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_40),
.B(n_258),
.Y(n_310)
);

AO22x1_ASAP7_75t_SL g591 ( 
.A1(n_40),
.A2(n_64),
.B1(n_312),
.B2(n_592),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_40),
.B(n_592),
.Y(n_622)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_46),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_46),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g485 ( 
.A(n_47),
.Y(n_485)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_49),
.Y(n_428)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_61),
.Y(n_595)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_63),
.A2(n_191),
.B1(n_192),
.B2(n_201),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_64),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_64),
.B(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_64),
.A2(n_443),
.B(n_446),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_76),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_135),
.B2(n_170),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B1(n_123),
.B2(n_132),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_81),
.A2(n_92),
.B1(n_132),
.B2(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_84),
.Y(n_304)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_84),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_85),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_86),
.A2(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_86),
.B(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_91),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_92),
.A2(n_123),
.B(n_132),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_92),
.A2(n_132),
.B1(n_176),
.B2(n_221),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g300 ( 
.A1(n_92),
.A2(n_134),
.B1(n_221),
.B2(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_92),
.B(n_333),
.Y(n_332)
);

AOI22x1_ASAP7_75t_L g454 ( 
.A1(n_92),
.A2(n_132),
.B1(n_328),
.B2(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_92),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B1(n_101),
.B2(n_104),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_97),
.Y(n_388)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_100),
.Y(n_376)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_106),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_111),
.Y(n_459)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_112),
.Y(n_481)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_126),
.Y(n_457)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_128),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_128),
.Y(n_436)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_133),
.A2(n_327),
.B(n_332),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_133),
.B(n_372),
.Y(n_507)
);

OAI22x1_ASAP7_75t_L g597 ( 
.A1(n_133),
.A2(n_477),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_134),
.B(n_333),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_135),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_175),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_151),
.B(n_163),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_136),
.A2(n_151),
.B1(n_163),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_136),
.B(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_136),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_136),
.B(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_136),
.A2(n_151),
.B1(n_364),
.B2(n_449),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_153),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B1(n_145),
.B2(n_147),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_142),
.Y(n_286)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g342 ( 
.A(n_143),
.Y(n_342)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_144),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_144),
.Y(n_503)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_144),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_146),
.Y(n_348)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_148),
.Y(n_536)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_151),
.B(n_364),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_151),
.B(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_152),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_152),
.A2(n_234),
.B1(n_292),
.B2(n_298),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_152),
.Y(n_353)
);

OA22x2_ASAP7_75t_L g585 ( 
.A1(n_152),
.A2(n_292),
.B1(n_298),
.B2(n_450),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_155),
.Y(n_362)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_162),
.Y(n_367)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_162),
.Y(n_473)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_168),
.B(n_372),
.Y(n_538)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_172),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.C(n_179),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_183),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_186),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_202),
.B2(n_203),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_189),
.B(n_203),
.C(n_666),
.Y(n_665)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_197),
.Y(n_425)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_SL g680 ( 
.A1(n_205),
.A2(n_681),
.B(n_682),
.C(n_683),
.Y(n_680)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_319),
.B(n_652),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_267),
.Y(n_207)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_208),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_264),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_209),
.B(n_264),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_229),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_212),
.A2(n_229),
.B1(n_230),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_213),
.A2(n_214),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_240),
.B(n_256),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B(n_240),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_232),
.B(n_233),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_240),
.A2(n_241),
.B1(n_256),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_240),
.A2(n_241),
.B1(n_602),
.B2(n_603),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_244),
.B(n_249),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_243),
.Y(n_414)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_244),
.B(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_244),
.A2(n_412),
.B1(n_413),
.B2(n_415),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_244),
.A2(n_514),
.B1(n_523),
.B2(n_525),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_244),
.B(n_415),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_245),
.Y(n_524)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_SL g506 ( 
.A(n_246),
.Y(n_506)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_248),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_253),
.Y(n_532)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_255),
.Y(n_350)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_255),
.Y(n_519)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_257),
.B(n_622),
.Y(n_621)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_262),
.Y(n_672)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_262),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_268),
.B(n_271),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.C(n_276),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_272),
.B(n_277),
.Y(n_609)
);

XNOR2x1_ASAP7_75t_L g608 ( 
.A(n_273),
.B(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_299),
.C(n_308),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_279),
.B(n_606),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

XOR2x2_ASAP7_75t_L g615 ( 
.A(n_280),
.B(n_616),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_287),
.B(n_288),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_281),
.A2(n_587),
.B(n_590),
.Y(n_586)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_282),
.Y(n_498)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_287),
.A2(n_337),
.B1(n_343),
.B2(n_346),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_287),
.A2(n_497),
.B(n_504),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_291),
.Y(n_616)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_298),
.A2(n_353),
.B1(n_354),
.B2(n_469),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_298),
.A2(n_469),
.B(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_298),
.B(n_372),
.Y(n_554)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_300),
.B(n_309),
.Y(n_606)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_301),
.Y(n_599)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_310),
.Y(n_446)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2x1p5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_643),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_578),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_460),
.B(n_576),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_402),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_324),
.B(n_577),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_351),
.C(n_369),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_325),
.B(n_463),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_334),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_326),
.A2(n_406),
.B(n_408),
.Y(n_405)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_333),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_335),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_407),
.Y(n_408)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_337),
.A2(n_390),
.B(n_393),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_344),
.Y(n_562)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_351),
.A2(n_352),
.B1(n_369),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_354),
.B(n_363),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_SL g551 ( 
.A1(n_356),
.A2(n_372),
.B(n_538),
.Y(n_551)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_359),
.Y(n_548)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_363),
.B(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_367),
.Y(n_451)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_389),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_370),
.B(n_389),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_375),
.B1(n_377),
.B2(n_381),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_372),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_372),
.B(n_560),
.Y(n_559)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_376),
.Y(n_380)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

INVx3_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_392),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_393),
.A2(n_515),
.B(n_524),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_397),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_441),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_409),
.B2(n_410),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_404),
.B(n_410),
.C(n_441),
.Y(n_642)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_422),
.Y(n_410)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_411),
.Y(n_624)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_422),
.B(n_624),
.Y(n_623)
);

AO32x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_426),
.A3(n_429),
.B1(n_432),
.B2(n_433),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_447),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g638 ( 
.A(n_442),
.B(n_448),
.C(n_454),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_454),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_456),
.A2(n_477),
.B(n_486),
.Y(n_619)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_487),
.B(n_575),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g575 ( 
.A(n_462),
.B(n_465),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.C(n_476),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_466),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_466),
.A2(n_490),
.B1(n_491),
.B2(n_493),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_476),
.Y(n_491)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_477),
.A2(n_478),
.B(n_486),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

OAI321xp33_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_511),
.A3(n_568),
.B1(n_572),
.B2(n_573),
.C(n_685),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_492),
.B(n_494),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_494),
.B(n_574),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_507),
.C(n_508),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_496),
.B(n_571),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_507),
.B(n_509),
.Y(n_571)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_512),
.A2(n_552),
.B(n_567),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_526),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_513),
.B(n_526),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_524),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_549),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_527),
.B(n_549),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_537),
.B1(n_539),
.B2(n_544),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_533),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_545),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_553),
.A2(n_556),
.B(n_566),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_554),
.B(n_555),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_557),
.B(n_558),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_559),
.B(n_563),
.Y(n_558)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_570),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_569),
.B(n_570),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_579),
.B(n_628),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_579),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_580),
.A2(n_607),
.B(n_610),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_580),
.B(n_607),
.Y(n_651)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_581),
.B(n_608),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_600),
.C(n_604),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_582),
.B(n_626),
.Y(n_625)
);

MAJx2_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_591),
.C(n_596),
.Y(n_582)
);

XOR2x1_ASAP7_75t_SL g613 ( 
.A(n_583),
.B(n_614),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_586),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_585),
.B(n_586),
.Y(n_636)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

XNOR2x1_ASAP7_75t_SL g614 ( 
.A(n_591),
.B(n_597),
.Y(n_614)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_595),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_601),
.Y(n_627)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_605),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_627),
.Y(n_626)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_625),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_611),
.B(n_625),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_615),
.C(n_617),
.Y(n_611)
);

INVxp33_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

XOR2x1_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_615),
.Y(n_630)
);

XNOR2x1_ASAP7_75t_L g629 ( 
.A(n_617),
.B(n_630),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_620),
.C(n_623),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_618),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.Y(n_634)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_623),
.B(n_634),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_629),
.A2(n_631),
.B(n_639),
.Y(n_628)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_629),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_632),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_645),
.C(n_646),
.Y(n_644)
);

MAJx2_ASAP7_75t_L g632 ( 
.A(n_633),
.B(n_635),
.C(n_637),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_633),
.B(n_641),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_638),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_640),
.B(n_642),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_640),
.B(n_642),
.Y(n_646)
);

AOI21x1_ASAP7_75t_L g643 ( 
.A1(n_644),
.A2(n_647),
.B(n_648),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_649),
.A2(n_650),
.B(n_651),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_653),
.A2(n_654),
.B(n_655),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_656),
.B(n_660),
.C(n_662),
.Y(n_682)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_659),
.B(n_662),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_660),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_663),
.B(n_677),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_665),
.B(n_667),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_665),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_668),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_668),
.B(n_679),
.Y(n_678)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_671),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_674),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_675),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g677 ( 
.A(n_678),
.Y(n_677)
);


endmodule