module fake_jpeg_1391_n_663 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_663);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_663;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_455;
wire n_544;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_19),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_13),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_5),
.B(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_58),
.Y(n_183)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_63),
.B(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_64),
.Y(n_186)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_72),
.Y(n_215)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_31),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_92),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_89),
.Y(n_210)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_44),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_95),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_0),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_97),
.B(n_98),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_99),
.B(n_102),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_103),
.Y(n_227)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_29),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_108),
.B(n_113),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_47),
.Y(n_110)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_2),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_49),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_3),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_47),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_120),
.B(n_32),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_21),
.Y(n_121)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_20),
.Y(n_122)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_129),
.Y(n_209)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_32),
.Y(n_130)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_149),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

BUFx24_ASAP7_75t_L g292 ( 
.A(n_159),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_166),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_69),
.A2(n_40),
.B1(n_32),
.B2(n_51),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_170),
.A2(n_84),
.B1(n_83),
.B2(n_77),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_172),
.B(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_214),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_82),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_212),
.Y(n_252)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_127),
.B(n_56),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_189),
.B(n_155),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_86),
.B(n_40),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_205),
.Y(n_247)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

INVx2_ASAP7_75t_R g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx9p33_ASAP7_75t_R g239 ( 
.A(n_204),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_112),
.B(n_40),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_66),
.Y(n_213)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_101),
.B(n_33),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_220),
.B(n_226),
.Y(n_268)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_67),
.Y(n_222)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_100),
.Y(n_224)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_71),
.B(n_25),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_74),
.B(n_33),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_25),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_56),
.B1(n_35),
.B2(n_51),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_232),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_236),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_132),
.Y(n_238)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_80),
.B1(n_115),
.B2(n_103),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_240),
.A2(n_267),
.B1(n_269),
.B2(n_273),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_241),
.B(n_251),
.C(n_261),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_40),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_243),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_188),
.A2(n_35),
.B(n_41),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_246),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_248),
.B(n_249),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_41),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_40),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_250),
.B(n_310),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_164),
.B(n_37),
.Y(n_251)
);

CKINVDCx12_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_253),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_154),
.B(n_55),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_256),
.B(n_258),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_117),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_142),
.Y(n_260)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_154),
.B(n_55),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_265),
.B(n_280),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_206),
.A2(n_94),
.B1(n_89),
.B2(n_88),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_173),
.A2(n_46),
.B1(n_37),
.B2(n_79),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_270),
.A2(n_290),
.B1(n_307),
.B2(n_146),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_271),
.B(n_289),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_195),
.A2(n_161),
.B1(n_135),
.B2(n_138),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_148),
.A2(n_46),
.B1(n_45),
.B2(n_6),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_134),
.Y(n_277)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_195),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_305),
.Y(n_328)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g342 ( 
.A(n_279),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_5),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_281),
.B(n_249),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_155),
.B(n_147),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_283),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_186),
.B(n_6),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_205),
.B(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_285),
.B(n_151),
.C(n_139),
.Y(n_352)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_201),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_190),
.B(n_7),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_288),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_196),
.B(n_7),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_211),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_131),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g293 ( 
.A1(n_170),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_139),
.B1(n_221),
.B2(n_227),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_149),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_294),
.B(n_297),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_153),
.B(n_10),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_165),
.B(n_13),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_180),
.B(n_13),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_143),
.B(n_14),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_298),
.B(n_301),
.Y(n_349)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_145),
.B(n_14),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_156),
.Y(n_303)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_142),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_162),
.B(n_15),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_183),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_150),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_308)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_187),
.B1(n_221),
.B2(n_152),
.Y(n_372)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_141),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

AO22x1_ASAP7_75t_L g310 ( 
.A1(n_183),
.A2(n_16),
.B1(n_19),
.B2(n_215),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_215),
.B(n_16),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_185),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_177),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_133),
.Y(n_313)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_344),
.B1(n_250),
.B2(n_243),
.Y(n_376)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_331),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_178),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_369),
.C(n_250),
.Y(n_385)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_240),
.A2(n_267),
.B1(n_273),
.B2(n_233),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_308),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_230),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_352),
.C(n_356),
.Y(n_408)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_254),
.Y(n_353)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_239),
.A2(n_268),
.B(n_310),
.C(n_293),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_355),
.A2(n_231),
.B(n_235),
.Y(n_418)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_255),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_259),
.Y(n_361)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_247),
.B(n_157),
.C(n_224),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_239),
.B(n_246),
.CI(n_247),
.CON(n_370),
.SN(n_370)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_187),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_252),
.A2(n_185),
.B1(n_210),
.B2(n_152),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_306),
.B1(n_284),
.B2(n_304),
.Y(n_403)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_242),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_374),
.B(n_375),
.Y(n_382)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_245),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_376),
.A2(n_384),
.B1(n_387),
.B2(n_404),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_332),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_377),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_302),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_379),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_275),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_334),
.A2(n_363),
.B1(n_356),
.B2(n_333),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_388),
.C(n_392),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_262),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_394),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_334),
.A2(n_278),
.B1(n_285),
.B2(n_243),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_285),
.C(n_313),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_317),
.B(n_245),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_391),
.B(n_395),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_262),
.C(n_279),
.Y(n_392)
);

OR2x4_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_244),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_393),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_364),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_263),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_397),
.C(n_352),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_286),
.C(n_309),
.Y(n_397)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_399),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_316),
.B(n_312),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_400),
.B(n_401),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_324),
.B(n_340),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_300),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_412),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_403),
.A2(n_329),
.B1(n_404),
.B2(n_421),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_334),
.A2(n_192),
.B1(n_210),
.B2(n_227),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_263),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_405),
.B(n_411),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_413),
.B(n_328),
.Y(n_434)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_244),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_359),
.B(n_349),
.Y(n_412)
);

OR2x4_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_292),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_347),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_422),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_318),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_345),
.B(n_235),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_420),
.B(n_423),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_372),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_335),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_330),
.B(n_276),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_382),
.Y(n_428)
);

INVx13_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_439),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_344),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_435),
.B(n_446),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_376),
.A2(n_413),
.B1(n_418),
.B2(n_408),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_437),
.A2(n_416),
.B1(n_415),
.B2(n_389),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_328),
.B(n_336),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_406),
.A2(n_372),
.B1(n_336),
.B2(n_325),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_450),
.B1(n_453),
.B2(n_458),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_427),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_377),
.B(n_365),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_444),
.B(n_462),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_419),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_409),
.A2(n_372),
.B1(n_171),
.B2(n_167),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_346),
.C(n_335),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_397),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_409),
.A2(n_163),
.B1(n_171),
.B2(n_167),
.Y(n_453)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_454),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_384),
.A2(n_342),
.B1(n_347),
.B2(n_323),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_455),
.A2(n_456),
.B1(n_460),
.B2(n_464),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_387),
.A2(n_342),
.B1(n_323),
.B2(n_350),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_457),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_393),
.A2(n_163),
.B1(n_238),
.B2(n_236),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_422),
.Y(n_459)
);

INVx13_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_392),
.A2(n_326),
.B1(n_350),
.B2(n_327),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_410),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_405),
.A2(n_318),
.B(n_315),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_395),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_388),
.A2(n_327),
.B1(n_319),
.B2(n_322),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_466),
.B(n_483),
.C(n_484),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_449),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_473),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_428),
.B(n_383),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_468),
.B(n_474),
.C(n_477),
.Y(n_531)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_403),
.B(n_419),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_454),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_447),
.B(n_443),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_449),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_501),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_315),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_338),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_479),
.B(n_489),
.Y(n_510)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_427),
.B(n_411),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_440),
.A2(n_416),
.B1(n_417),
.B2(n_399),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g503 ( 
.A(n_487),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_389),
.Y(n_488)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_338),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_490),
.B(n_498),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_426),
.A2(n_415),
.B1(n_390),
.B2(n_414),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_492),
.A2(n_448),
.B1(n_444),
.B2(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_494),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_390),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_495),
.B(n_496),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_424),
.B(n_407),
.Y(n_496)
);

OA22x2_ASAP7_75t_L g498 ( 
.A1(n_426),
.A2(n_455),
.B1(n_445),
.B2(n_456),
.Y(n_498)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_451),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_451),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_407),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_SL g502 ( 
.A(n_445),
.B(n_331),
.C(n_292),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_472),
.C(n_490),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_434),
.B(n_446),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_504),
.A2(n_517),
.B(n_530),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_441),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_512),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_491),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_506),
.B(n_516),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_507),
.A2(n_538),
.B1(n_471),
.B2(n_470),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_488),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_509),
.B(n_524),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_452),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_454),
.Y(n_514)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_430),
.Y(n_515)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_515),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_491),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_499),
.A2(n_446),
.B(n_436),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_465),
.A2(n_448),
.B1(n_436),
.B2(n_435),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_521),
.A2(n_525),
.B1(n_431),
.B2(n_425),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_430),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_523),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_473),
.B(n_460),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_501),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_465),
.A2(n_450),
.B1(n_458),
.B2(n_439),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_442),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_526),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_532),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_499),
.A2(n_463),
.B(n_442),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_462),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_466),
.B(n_464),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_486),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_425),
.Y(n_563)
);

AO22x1_ASAP7_75t_L g538 ( 
.A1(n_472),
.A2(n_453),
.B1(n_461),
.B2(n_431),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_498),
.C(n_492),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_539),
.B(n_541),
.C(n_565),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_498),
.C(n_485),
.Y(n_541)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_542),
.A2(n_519),
.B(n_523),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_515),
.A2(n_481),
.B1(n_478),
.B2(n_471),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_546),
.A2(n_549),
.B1(n_552),
.B2(n_560),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_480),
.C(n_481),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_551),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_529),
.B(n_480),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_548),
.B(n_536),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_521),
.A2(n_478),
.B1(n_471),
.B2(n_498),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_520),
.B(n_534),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_553),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_502),
.C(n_470),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_522),
.A2(n_471),
.B1(n_493),
.B2(n_494),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_504),
.B(n_469),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_562),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_508),
.A2(n_475),
.B1(n_469),
.B2(n_497),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_556),
.A2(n_558),
.B1(n_535),
.B2(n_528),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_508),
.A2(n_475),
.B1(n_497),
.B2(n_500),
.Y(n_558)
);

XOR2x2_ASAP7_75t_L g562 ( 
.A(n_517),
.B(n_425),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_563),
.B(n_511),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_398),
.C(n_380),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_537),
.B(n_380),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_514),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_533),
.A2(n_451),
.B1(n_366),
.B2(n_398),
.Y(n_567)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_567),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_506),
.A2(n_366),
.B1(n_319),
.B2(n_260),
.Y(n_568)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_568),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_555),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_583),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_564),
.A2(n_516),
.B1(n_519),
.B2(n_525),
.Y(n_572)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_572),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_576),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_577),
.A2(n_549),
.B(n_552),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_581),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_555),
.A2(n_530),
.B(n_510),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_580),
.B(n_559),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_582),
.B(n_339),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_511),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_545),
.B(n_518),
.C(n_519),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_565),
.C(n_539),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_513),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_588),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_543),
.B(n_526),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_586),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_554),
.B(n_513),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_589),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_566),
.B(n_550),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_590),
.B(n_592),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_546),
.A2(n_507),
.B1(n_518),
.B2(n_538),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_591),
.A2(n_542),
.B1(n_561),
.B2(n_544),
.Y(n_596)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_SL g628 ( 
.A(n_594),
.B(n_272),
.Y(n_628)
);

OAI31xp33_ASAP7_75t_SL g595 ( 
.A1(n_572),
.A2(n_562),
.A3(n_557),
.B(n_553),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_595),
.B(n_601),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_596),
.A2(n_604),
.B1(n_571),
.B2(n_587),
.Y(n_613)
);

AO221x1_ASAP7_75t_L g599 ( 
.A1(n_591),
.A2(n_556),
.B1(n_558),
.B2(n_536),
.C(n_538),
.Y(n_599)
);

INVxp33_ASAP7_75t_SL g619 ( 
.A(n_599),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_545),
.C(n_557),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_600),
.B(n_603),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_602),
.A2(n_231),
.B(n_136),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_559),
.C(n_532),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_571),
.A2(n_535),
.B1(n_503),
.B2(n_528),
.Y(n_604)
);

AOI322xp5_ASAP7_75t_L g605 ( 
.A1(n_569),
.A2(n_503),
.A3(n_272),
.B1(n_299),
.B2(n_216),
.C1(n_197),
.C2(n_200),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_605),
.B(n_299),
.Y(n_627)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_609),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_588),
.B(n_360),
.Y(n_610)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_610),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_613),
.B(n_615),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_583),
.C(n_584),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_618),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_603),
.B(n_574),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_575),
.B1(n_574),
.B2(n_578),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_617),
.A2(n_625),
.B1(n_627),
.B2(n_606),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_581),
.C(n_585),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_597),
.B(n_590),
.C(n_573),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_607),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_602),
.A2(n_573),
.B(n_257),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_622),
.A2(n_628),
.B(n_595),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_606),
.A2(n_596),
.B1(n_601),
.B2(n_593),
.Y(n_625)
);

MAJx2_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_609),
.C(n_599),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_623),
.B(n_608),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_632),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_631),
.A2(n_638),
.B1(n_626),
.B2(n_625),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_617),
.A2(n_612),
.B(n_598),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_633),
.B(n_634),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_618),
.B(n_612),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_611),
.C(n_597),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_635),
.B(n_636),
.C(n_637),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_619),
.A2(n_611),
.B1(n_610),
.B2(n_229),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_SL g640 ( 
.A(n_621),
.B(n_272),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_R g647 ( 
.A1(n_640),
.A2(n_229),
.B1(n_264),
.B2(n_158),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_630),
.A2(n_624),
.B1(n_616),
.B2(n_615),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_642),
.B(n_264),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_644),
.B(n_647),
.Y(n_650)
);

OAI221xp5_ASAP7_75t_L g645 ( 
.A1(n_638),
.A2(n_613),
.B1(n_621),
.B2(n_620),
.C(n_272),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_645),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_639),
.A2(n_299),
.B(n_264),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_648),
.B(n_237),
.C(n_158),
.Y(n_653)
);

AOI322xp5_ASAP7_75t_L g649 ( 
.A1(n_641),
.A2(n_639),
.A3(n_640),
.B1(n_636),
.B2(n_216),
.C1(n_257),
.C2(n_209),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_649),
.B(n_651),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_653),
.B(n_229),
.Y(n_655)
);

FAx1_ASAP7_75t_SL g654 ( 
.A(n_652),
.B(n_643),
.CI(n_646),
.CON(n_654),
.SN(n_654)
);

OAI331xp33_ASAP7_75t_L g658 ( 
.A1(n_654),
.A2(n_650),
.A3(n_653),
.B1(n_217),
.B2(n_166),
.B3(n_237),
.C1(n_175),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_655),
.B(n_647),
.C(n_648),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_657),
.B(n_658),
.Y(n_659)
);

AO21x1_ASAP7_75t_L g660 ( 
.A1(n_659),
.A2(n_654),
.B(n_656),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_650),
.Y(n_661)
);

BUFx24_ASAP7_75t_SL g662 ( 
.A(n_661),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_662),
.B(n_137),
.Y(n_663)
);


endmodule