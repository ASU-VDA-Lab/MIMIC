module real_jpeg_28799_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_0),
.A2(n_61),
.B1(n_62),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_0),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_140),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_140),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_140),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_1),
.B(n_57),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_44),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_44),
.B(n_227),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_186),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_30),
.B(n_33),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_136),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_1),
.A2(n_85),
.B1(n_132),
.B2(n_275),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_7),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_188),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_188),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_188),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_8),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_167),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_167),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_167),
.Y(n_267)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_11),
.A2(n_33),
.B1(n_35),
.B2(n_54),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_48)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_13),
.Y(n_226)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_64),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_15),
.A2(n_33),
.B1(n_35),
.B2(n_64),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_98),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_82),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_21),
.A2(n_22),
.B1(n_72),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_22)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_24),
.A2(n_25),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_40),
.C(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_26),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_26),
.A2(n_32),
.B1(n_93),
.B2(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_26),
.A2(n_36),
.B(n_94),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_26),
.A2(n_32),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_26),
.A2(n_77),
.B(n_235),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_26),
.A2(n_32),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_26),
.A2(n_32),
.B1(n_234),
.B2(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_28),
.A2(n_45),
.A3(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_29),
.B(n_225),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_29),
.A2(n_31),
.B(n_186),
.C(n_254),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_32),
.A2(n_79),
.B(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_32),
.B(n_186),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_35),
.B(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_37),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B(n_52),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_41),
.A2(n_52),
.B(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_41),
.A2(n_108),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_53),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_42),
.A2(n_48),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_42),
.A2(n_48),
.B1(n_182),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_42),
.A2(n_48),
.B1(n_210),
.B2(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_44),
.B(n_58),
.Y(n_199)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_45),
.A2(n_67),
.B1(n_185),
.B2(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_71),
.B1(n_100),
.B2(n_112),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_65),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_60),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_56),
.A2(n_102),
.B1(n_139),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_56),
.A2(n_102),
.B1(n_166),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_58),
.B(n_62),
.C(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_57),
.B(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_57),
.A2(n_66),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_62),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_62),
.B(n_186),
.CON(n_185),
.SN(n_185)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_110),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_83),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B(n_95),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_95),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_92),
.B1(n_121),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_85),
.A2(n_132),
.B1(n_158),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_85),
.A2(n_130),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_85),
.A2(n_214),
.B1(n_267),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_86),
.A2(n_90),
.B(n_160),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_86),
.A2(n_131),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_92),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_111),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_146),
.B(n_319),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_142),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_117),
.B(n_142),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_123),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_122),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_124),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.C(n_137),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_126),
.B(n_133),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_201),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_171),
.B(n_318),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_168),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_148),
.B(n_168),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_155),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_153),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_155),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.C(n_164),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_156),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_162),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_312),
.B(n_317),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_215),
.B(n_298),
.C(n_311),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_202),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_174),
.B(n_202),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_189),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_176),
.B(n_177),
.C(n_189),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_186),
.B(n_214),
.Y(n_279)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_197),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_191),
.B(n_195),
.C(n_197),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_200),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.C(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_203),
.A2(n_204),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.C(n_213),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_297),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_290),
.B(n_296),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_245),
.B(n_289),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_236),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_219),
.B(n_236),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_229),
.C(n_232),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_220),
.A2(n_221),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_223),
.Y(n_243)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_243),
.C(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_283),
.B(n_288),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_263),
.B(n_282),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_262),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_271),
.B(n_281),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_269),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_276),
.B(n_280),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_309),
.B2(n_310),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_306),
.C(n_310),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);


endmodule