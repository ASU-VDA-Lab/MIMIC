module fake_ariane_571_n_1771 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1771);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1771;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_89),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_47),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_24),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_156),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_40),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_106),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_6),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_40),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_59),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_23),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_56),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_33),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_71),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_23),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_83),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_55),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_65),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_143),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_123),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_137),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_60),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_16),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_51),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_100),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_35),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_91),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_74),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_30),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_113),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_80),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_78),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_62),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_155),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_87),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_101),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_13),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_52),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_129),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_109),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_110),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_145),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_130),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_31),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_29),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_81),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_41),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_34),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_118),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_8),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_20),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_4),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_63),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_116),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_48),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_98),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_93),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_2),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_117),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_50),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_128),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_121),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_49),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_105),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_124),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_34),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_133),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_73),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_66),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_102),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_122),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_28),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_57),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_115),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_30),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_72),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_46),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_45),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_138),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_12),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_27),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_24),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_205),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_236),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_177),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_161),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_168),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_202),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_180),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_297),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_207),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_220),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_224),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_168),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_191),
.B(n_1),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_224),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_194),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_194),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_293),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_295),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_266),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_167),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_178),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_314),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_285),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_204),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_179),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_200),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_179),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_214),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_240),
.B(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_185),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_223),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_228),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_240),
.B(n_3),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_226),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_170),
.B(n_3),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_226),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_241),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_226),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_240),
.B(n_267),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_285),
.B(n_4),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_285),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_164),
.B(n_169),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_258),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_248),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_214),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_170),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_286),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_248),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_171),
.B(n_7),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_271),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_248),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_300),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_287),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_296),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_217),
.B(n_10),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_270),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_246),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

AND3x2_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_165),
.C(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_359),
.B(n_270),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_246),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_270),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_371),
.B(n_359),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_272),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_333),
.B(n_187),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_176),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_326),
.B(n_283),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_318),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_333),
.B(n_210),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_332),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_352),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_374),
.B(n_376),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_272),
.Y(n_438)
);

AND3x1_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_300),
.C(n_221),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_213),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_343),
.B(n_229),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_338),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_383),
.B(n_167),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_389),
.A2(n_255),
.B(n_235),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_390),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_391),
.B(n_265),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_391),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_346),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_392),
.A2(n_278),
.B(n_274),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_325),
.B(n_281),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_345),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_349),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_360),
.B(n_284),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_361),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_321),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_362),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_421),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_365),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_422),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_412),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_394),
.B(n_393),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_365),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_395),
.A2(n_354),
.B1(n_344),
.B2(n_382),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_421),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_395),
.A2(n_355),
.B1(n_353),
.B2(n_369),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_329),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_172),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

CKINVDCx6p67_ASAP7_75t_R g491 ( 
.A(n_453),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_410),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_406),
.B(n_367),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_399),
.B(n_395),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_399),
.B(n_367),
.Y(n_496)
);

OA22x2_ASAP7_75t_L g497 ( 
.A1(n_397),
.A2(n_366),
.B1(n_387),
.B2(n_373),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_446),
.Y(n_498)
);

AOI22x1_ASAP7_75t_L g499 ( 
.A1(n_395),
.A2(n_176),
.B1(n_181),
.B2(n_183),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_398),
.B(n_329),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_433),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_406),
.B(n_386),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_395),
.B(n_377),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_428),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_395),
.B(n_437),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_445),
.B(n_172),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_377),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_398),
.A2(n_319),
.B1(n_375),
.B2(n_303),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_452),
.B(n_351),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_424),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_422),
.B(n_386),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_439),
.A2(n_348),
.B1(n_366),
.B2(n_198),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_445),
.B(n_172),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_446),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_394),
.B(n_372),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_438),
.A2(n_456),
.B1(n_455),
.B2(n_440),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_410),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_396),
.B(n_378),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_283),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_410),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_394),
.B(n_320),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_405),
.B(n_350),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_449),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_405),
.B(n_283),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_405),
.B(n_324),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_439),
.B(n_160),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_462),
.B(n_160),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_438),
.B(n_250),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_438),
.B(n_441),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_464),
.B(n_290),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_438),
.B(n_167),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_459),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_416),
.B(n_183),
.C(n_181),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_455),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_445),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_458),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_416),
.A2(n_243),
.B1(n_233),
.B2(n_237),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_449),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_438),
.B(n_167),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_414),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_430),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_438),
.B(n_327),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_408),
.B(n_273),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_408),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_430),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_462),
.A2(n_282),
.B1(n_184),
.B2(n_189),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_408),
.B(n_162),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_462),
.B(n_330),
.Y(n_584)
);

AND3x2_ASAP7_75t_L g585 ( 
.A(n_396),
.B(n_342),
.C(n_341),
.Y(n_585)
);

AOI22x1_ASAP7_75t_L g586 ( 
.A1(n_447),
.A2(n_454),
.B1(n_418),
.B2(n_417),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_456),
.A2(n_290),
.B1(n_215),
.B2(n_263),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_408),
.B(n_423),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_449),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_423),
.A2(n_216),
.B1(n_230),
.B2(n_231),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_408),
.B(n_331),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_408),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_449),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_433),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_460),
.A2(n_317),
.B1(n_315),
.B2(n_313),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_440),
.B(n_162),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_460),
.A2(n_315),
.B1(n_313),
.B2(n_311),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_430),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_449),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_430),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_449),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_440),
.B(n_166),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_456),
.B(n_167),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_414),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_434),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_418),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_434),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_434),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_418),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_434),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_440),
.B(n_166),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_440),
.B(n_173),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_397),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_434),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_455),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_490),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_559),
.B(n_576),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_559),
.B(n_440),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_494),
.A2(n_304),
.B1(n_189),
.B2(n_184),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_451),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_566),
.B(n_451),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_555),
.B(n_451),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_537),
.A2(n_455),
.B1(n_445),
.B2(n_451),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_470),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_510),
.B(n_445),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_492),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_486),
.B(n_451),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_515),
.B(n_456),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_468),
.A2(n_311),
.B1(n_310),
.B2(n_304),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_474),
.B(n_458),
.Y(n_632)
);

XOR2x2_ASAP7_75t_L g633 ( 
.A(n_485),
.B(n_455),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_496),
.B(n_451),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_513),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_504),
.B(n_456),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

BUFx4_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_513),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_501),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_456),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_587),
.A2(n_301),
.B1(n_282),
.B2(n_291),
.C(n_298),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_L g645 ( 
.A(n_491),
.B(n_291),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_538),
.B(n_299),
.C(n_298),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_550),
.A2(n_463),
.B1(n_461),
.B2(n_458),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_564),
.A2(n_310),
.B1(n_301),
.B2(n_299),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_607),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_568),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_541),
.B(n_417),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_566),
.A2(n_448),
.B(n_447),
.C(n_454),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_541),
.B(n_418),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_568),
.A2(n_219),
.B1(n_193),
.B2(n_209),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_464),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_550),
.B(n_418),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_469),
.B(n_458),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_469),
.B(n_458),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_566),
.B(n_458),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_614),
.B(n_464),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_522),
.B(n_458),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_554),
.B(n_458),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_481),
.B(n_461),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_490),
.B(n_461),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_481),
.B(n_461),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_523),
.A2(n_464),
.B1(n_447),
.B2(n_454),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_466),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_447),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_536),
.B(n_461),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_481),
.B(n_461),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_475),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_500),
.B(n_461),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_493),
.B(n_461),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_490),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_475),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_480),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_547),
.B(n_463),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_479),
.B(n_463),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_503),
.B(n_473),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_516),
.A2(n_454),
.B(n_417),
.C(n_419),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_463),
.Y(n_682)
);

BUFx6f_ASAP7_75t_SL g683 ( 
.A(n_473),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_610),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_473),
.B(n_463),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_517),
.A2(n_455),
.B1(n_419),
.B2(n_420),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_482),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_539),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_482),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_562),
.B(n_463),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_594),
.B(n_290),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_473),
.B(n_588),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_565),
.B(n_463),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_584),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_488),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_560),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_553),
.B(n_463),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_479),
.B(n_448),
.Y(n_698)
);

CKINVDCx11_ASAP7_75t_R g699 ( 
.A(n_582),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_525),
.B(n_429),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_479),
.B(n_448),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_539),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_552),
.B(n_429),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_490),
.B(n_173),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_580),
.B(n_419),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_580),
.B(n_420),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_592),
.B(n_420),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_490),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_499),
.B(n_174),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_592),
.A2(n_402),
.B1(n_403),
.B2(n_409),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_488),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_505),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_551),
.B(n_436),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_579),
.B(n_402),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_603),
.B(n_403),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_505),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_596),
.B(n_409),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_531),
.A2(n_415),
.B(n_407),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_518),
.B(n_415),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_436),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_518),
.B(n_427),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_563),
.B(n_279),
.C(n_212),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_501),
.B(n_238),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_526),
.B(n_427),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_509),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_526),
.Y(n_726)
);

NOR2x1p5_ASAP7_75t_SL g727 ( 
.A(n_467),
.B(n_172),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_613),
.B(n_443),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_548),
.B(n_443),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_509),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_499),
.A2(n_276),
.B1(n_239),
.B2(n_247),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_614),
.B(n_444),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_517),
.A2(n_425),
.B1(n_442),
.B2(n_435),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_512),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_507),
.B(n_174),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_512),
.B(n_427),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_514),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_514),
.B(n_431),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_520),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_495),
.B(n_434),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_546),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_520),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_483),
.B(n_444),
.Y(n_744)
);

AO221x1_ASAP7_75t_L g745 ( 
.A1(n_517),
.A2(n_434),
.B1(n_431),
.B2(n_432),
.C(n_435),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_517),
.A2(n_435),
.B1(n_432),
.B2(n_425),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_527),
.A2(n_431),
.B(n_435),
.C(n_432),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_583),
.B(n_434),
.Y(n_748)
);

NOR2x1_ASAP7_75t_L g749 ( 
.A(n_591),
.B(n_425),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_616),
.A2(n_442),
.B1(n_432),
.B2(n_425),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_560),
.A2(n_182),
.B1(n_307),
.B2(n_305),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_527),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_590),
.B(n_595),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_530),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_530),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_560),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_560),
.B(n_442),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_467),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_597),
.B(n_175),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_471),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_575),
.B(n_442),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_571),
.B(n_175),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_575),
.B(n_182),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_575),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_471),
.Y(n_765)
);

AND2x2_ASAP7_75t_SL g766 ( 
.A(n_487),
.B(n_401),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_575),
.B(n_188),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_616),
.B(n_188),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_604),
.B(n_251),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_604),
.A2(n_495),
.B1(n_528),
.B2(n_511),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_604),
.B(n_190),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_604),
.B(n_190),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_495),
.B(n_252),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_507),
.B(n_192),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_586),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_497),
.B(n_256),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_585),
.B(n_269),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_608),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_608),
.B(n_192),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_507),
.B(n_280),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_497),
.A2(n_280),
.B1(n_289),
.B2(n_292),
.C(n_294),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_608),
.B(n_289),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_476),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_497),
.A2(n_292),
.B1(n_294),
.B2(n_305),
.C(n_307),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_476),
.B(n_11),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_753),
.A2(n_544),
.B(n_531),
.C(n_535),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_660),
.A2(n_544),
.B(n_569),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_656),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_655),
.B(n_472),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_472),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_669),
.B(n_472),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_660),
.A2(n_572),
.B(n_589),
.Y(n_793)
);

AOI21xp33_ASAP7_75t_L g794 ( 
.A1(n_742),
.A2(n_487),
.B(n_511),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_502),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_698),
.A2(n_572),
.B(n_535),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_641),
.B(n_508),
.Y(n_797)
);

AOI21xp33_ASAP7_75t_L g798 ( 
.A1(n_736),
.A2(n_528),
.B(n_570),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_696),
.B(n_508),
.Y(n_799)
);

AOI21xp33_ASAP7_75t_L g800 ( 
.A1(n_732),
.A2(n_570),
.B(n_569),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_628),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_723),
.B(n_498),
.Y(n_802)
);

O2A1O1Ixp5_ASAP7_75t_L g803 ( 
.A1(n_709),
.A2(n_502),
.B(n_529),
.C(n_540),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_661),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_729),
.B(n_502),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_652),
.A2(n_549),
.B(n_589),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_624),
.A2(n_549),
.B(n_593),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_688),
.B(n_702),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_692),
.B(n_529),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_632),
.A2(n_593),
.B(n_598),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_684),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_642),
.B(n_615),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_626),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_627),
.A2(n_598),
.B(n_529),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_649),
.B(n_507),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_662),
.A2(n_540),
.B(n_600),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_622),
.A2(n_540),
.B(n_600),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_712),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_649),
.B(n_507),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_630),
.A2(n_615),
.B(n_611),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_732),
.B(n_602),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_630),
.A2(n_498),
.B(n_609),
.C(n_477),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_623),
.A2(n_602),
.B(n_609),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_664),
.A2(n_611),
.B(n_477),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_629),
.B(n_478),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_626),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_651),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_664),
.A2(n_478),
.B(n_484),
.Y(n_829)
);

NOR2x1p5_ASAP7_75t_L g830 ( 
.A(n_770),
.B(n_484),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_649),
.B(n_524),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_649),
.B(n_524),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_651),
.B(n_489),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_640),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_651),
.B(n_489),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_633),
.A2(n_745),
.B1(n_686),
.B2(n_625),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_666),
.A2(n_542),
.B(n_506),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_666),
.A2(n_542),
.B(n_506),
.Y(n_838)
);

INVx11_ASAP7_75t_L g839 ( 
.A(n_651),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_741),
.A2(n_556),
.B(n_599),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_670),
.A2(n_543),
.B(n_521),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_651),
.B(n_521),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_634),
.A2(n_543),
.B(n_534),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_725),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_668),
.B(n_534),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_649),
.B(n_524),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_649),
.B(n_524),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_781),
.A2(n_556),
.B(n_573),
.C(n_599),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_744),
.B(n_573),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_661),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_692),
.A2(n_574),
.B1(n_577),
.B2(n_581),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_620),
.A2(n_574),
.B1(n_577),
.B2(n_581),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_657),
.B(n_524),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_770),
.B(n_532),
.Y(n_854)
);

O2A1O1Ixp5_ASAP7_75t_L g855 ( 
.A1(n_781),
.A2(n_400),
.B(n_401),
.C(n_407),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_661),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_637),
.A2(n_606),
.B1(n_601),
.B2(n_532),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_696),
.B(n_508),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_740),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_653),
.B(n_532),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_694),
.B(n_778),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_637),
.A2(n_606),
.B1(n_601),
.B2(n_532),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_644),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_679),
.A2(n_606),
.B(n_601),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_700),
.B(n_532),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_703),
.A2(n_606),
.B(n_601),
.C(n_533),
.Y(n_866)
);

NOR2x1p5_ASAP7_75t_L g867 ( 
.A(n_639),
.B(n_533),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_679),
.A2(n_533),
.B(n_558),
.Y(n_868)
);

AOI21xp33_ASAP7_75t_L g869 ( 
.A1(n_621),
.A2(n_533),
.B(n_558),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_703),
.B(n_533),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_671),
.A2(n_567),
.B(n_558),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_631),
.A2(n_225),
.B(n_222),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_715),
.A2(n_567),
.B(n_558),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_756),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_766),
.B(n_508),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_714),
.B(n_508),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_625),
.A2(n_567),
.B1(n_558),
.B2(n_400),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_766),
.B(n_567),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_748),
.A2(n_567),
.B(n_411),
.Y(n_879)
);

INVx6_ASAP7_75t_L g880 ( 
.A(n_640),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_748),
.A2(n_411),
.B(n_407),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_764),
.B(n_400),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_737),
.A2(n_411),
.B(n_407),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_739),
.A2(n_411),
.B(n_401),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_721),
.A2(n_724),
.B(n_701),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_680),
.B(n_11),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_698),
.A2(n_401),
.B(n_400),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_618),
.B(n_172),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_701),
.A2(n_400),
.B(n_404),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_672),
.A2(n_232),
.B(n_277),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_672),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_747),
.A2(n_227),
.B(n_275),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_676),
.A2(n_218),
.B(n_268),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_680),
.B(n_617),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_726),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_643),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_743),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_769),
.A2(n_195),
.B(n_260),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_645),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_R g900 ( 
.A(n_691),
.B(n_196),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_676),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_717),
.B(n_199),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_636),
.B(n_14),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_717),
.A2(n_242),
.B(n_259),
.C(n_257),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_720),
.B(n_201),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_L g907 ( 
.A1(n_731),
.A2(n_203),
.B(n_206),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_677),
.A2(n_234),
.B(n_253),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_720),
.B(n_249),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_677),
.A2(n_244),
.B(n_208),
.Y(n_910)
);

CKINVDCx8_ASAP7_75t_R g911 ( 
.A(n_774),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_638),
.B(n_15),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_SL g913 ( 
.A1(n_776),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_913)
);

OAI22xp33_ASAP7_75t_L g914 ( 
.A1(n_782),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_687),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_650),
.B(n_19),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_774),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_768),
.A2(n_404),
.B(n_211),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_728),
.B(n_25),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_750),
.A2(n_211),
.B(n_172),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_689),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_728),
.B(n_26),
.Y(n_922)
);

AOI221x1_ASAP7_75t_L g923 ( 
.A1(n_674),
.A2(n_685),
.B1(n_722),
.B2(n_697),
.C(n_663),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_685),
.A2(n_404),
.B(n_32),
.C(n_36),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_695),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_647),
.B(n_667),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_750),
.A2(n_211),
.B(n_172),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_695),
.A2(n_404),
.B(n_211),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_749),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_711),
.A2(n_211),
.B(n_172),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_711),
.A2(n_64),
.B(n_150),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_730),
.A2(n_159),
.B(n_146),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_763),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_730),
.A2(n_132),
.B(n_131),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_734),
.A2(n_126),
.B(n_114),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_734),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_618),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_710),
.B(n_31),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_738),
.A2(n_104),
.B(n_97),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_738),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_762),
.B(n_785),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_779),
.B(n_32),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_686),
.B(n_36),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_752),
.A2(n_94),
.B(n_90),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_SL g945 ( 
.A(n_618),
.B(n_37),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_752),
.A2(n_85),
.B(n_76),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_673),
.A2(n_68),
.B(n_67),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_754),
.B(n_38),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_754),
.A2(n_38),
.B(n_39),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_755),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_618),
.B(n_42),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_755),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_678),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_682),
.A2(n_58),
.B(n_45),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_758),
.A2(n_44),
.B(n_47),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_733),
.B(n_44),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_733),
.B(n_746),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_690),
.A2(n_50),
.B(n_53),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_693),
.A2(n_53),
.B(n_54),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_719),
.A2(n_54),
.B(n_55),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_658),
.A2(n_57),
.B(n_58),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_659),
.A2(n_765),
.B(n_784),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_746),
.B(n_705),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_759),
.A2(n_697),
.B1(n_683),
.B2(n_646),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_681),
.A2(n_707),
.B(n_706),
.C(n_771),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_758),
.A2(n_760),
.B(n_784),
.Y(n_966)
);

INVx11_ASAP7_75t_L g967 ( 
.A(n_683),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_635),
.B(n_783),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_699),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_635),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_757),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_918),
.A2(n_786),
.B(n_718),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_789),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_808),
.Y(n_974)
);

NOR2x1_ASAP7_75t_L g975 ( 
.A(n_895),
.B(n_767),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_811),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_971),
.B(n_779),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_SL g978 ( 
.A(n_914),
.B(n_648),
.C(n_654),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_911),
.B(n_751),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_854),
.B(n_675),
.Y(n_981)
);

CKINVDCx8_ASAP7_75t_R g982 ( 
.A(n_856),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_809),
.B(n_760),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_919),
.A2(n_783),
.B(n_674),
.C(n_780),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_809),
.B(n_765),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_SL g986 ( 
.A1(n_951),
.A2(n_772),
.B(n_773),
.C(n_761),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_885),
.A2(n_665),
.B(n_675),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_801),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_917),
.B(n_777),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_867),
.B(n_675),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_967),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_828),
.B(n_675),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_933),
.B(n_708),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_836),
.A2(n_957),
.B1(n_886),
.B2(n_941),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_937),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_886),
.A2(n_727),
.B(n_704),
.C(n_735),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_894),
.B(n_708),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_849),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_818),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_804),
.B(n_718),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_941),
.A2(n_775),
.B(n_708),
.C(n_718),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_900),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_830),
.B(n_708),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_922),
.A2(n_896),
.B(n_904),
.C(n_924),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_895),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_836),
.A2(n_804),
.B1(n_850),
.B2(n_956),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_969),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_812),
.B(n_825),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_844),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_859),
.B(n_897),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_904),
.A2(n_924),
.B(n_914),
.C(n_938),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_900),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_845),
.B(n_874),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_L g1014 ( 
.A1(n_964),
.A2(n_899),
.B1(n_874),
.B2(n_943),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_968),
.A2(n_826),
.B(n_870),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_965),
.A2(n_951),
.B(n_902),
.C(n_909),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_795),
.B(n_805),
.Y(n_1017)
);

OAI21xp33_ASAP7_75t_SL g1018 ( 
.A1(n_955),
.A2(n_839),
.B(n_942),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_929),
.B(n_906),
.Y(n_1019)
);

BUFx2_ASAP7_75t_SL g1020 ( 
.A(n_861),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_828),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_880),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_SL g1023 ( 
.A1(n_903),
.A2(n_912),
.B1(n_916),
.B2(n_898),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_915),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_865),
.A2(n_862),
.B(n_857),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_858),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_797),
.B(n_794),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_815),
.A2(n_819),
.B(n_846),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_937),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_858),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_815),
.A2(n_819),
.B(n_846),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_903),
.A2(n_916),
.B1(n_912),
.B2(n_872),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_925),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_880),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_963),
.A2(n_921),
.B1(n_936),
.B2(n_863),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_880),
.B(n_834),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_813),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_965),
.A2(n_926),
.B(n_942),
.C(n_853),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_891),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_831),
.A2(n_832),
.B(n_847),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_834),
.B(n_905),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_940),
.B(n_950),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_940),
.B(n_950),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_799),
.B(n_802),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_882),
.B(n_905),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_831),
.A2(n_832),
.B(n_847),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_827),
.B(n_901),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_866),
.A2(n_803),
.B(n_888),
.C(n_848),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_843),
.A2(n_816),
.B(n_814),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_882),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_821),
.A2(n_792),
.B1(n_790),
.B2(n_948),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_953),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_851),
.B(n_960),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_907),
.B(n_970),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_791),
.A2(n_822),
.B1(n_853),
.B2(n_860),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_913),
.A2(n_822),
.B(n_866),
.C(n_954),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_860),
.B(n_876),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_920),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_961),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_875),
.A2(n_878),
.B1(n_842),
.B2(n_833),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_913),
.A2(n_958),
.B(n_949),
.C(n_798),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_937),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_923),
.B(n_807),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_799),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_835),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_889),
.A2(n_796),
.B(n_887),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_852),
.A2(n_787),
.B(n_892),
.C(n_800),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_820),
.A2(n_910),
.B(n_890),
.C(n_908),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_888),
.B(n_893),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_945),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_875),
.B(n_878),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_877),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_869),
.B(n_934),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_927),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_966),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_962),
.B(n_817),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_841),
.B(n_930),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_947),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_806),
.A2(n_823),
.B(n_855),
.C(n_840),
.Y(n_1081)
);

AOI32xp33_ASAP7_75t_L g1082 ( 
.A1(n_931),
.A2(n_946),
.A3(n_944),
.B1(n_939),
.B2(n_935),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_864),
.B(n_873),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_824),
.A2(n_837),
.B(n_838),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_829),
.A2(n_788),
.B(n_793),
.Y(n_1085)
);

CKINVDCx14_ASAP7_75t_R g1086 ( 
.A(n_932),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_883),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_884),
.B(n_881),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_810),
.A2(n_879),
.B(n_868),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_871),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_928),
.B(n_624),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_919),
.A2(n_753),
.B(n_496),
.C(n_736),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_839),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_889),
.A2(n_796),
.B(n_918),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_971),
.B(n_624),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_937),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_858),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_886),
.A2(n_742),
.B1(n_492),
.B2(n_545),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_854),
.B(n_661),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_836),
.A2(n_633),
.B1(n_578),
.B2(n_497),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_789),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_828),
.B(n_797),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_885),
.A2(n_968),
.B(n_826),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_828),
.B(n_628),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_885),
.A2(n_968),
.B(n_826),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_911),
.B(n_742),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_914),
.B(n_742),
.C(n_753),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_867),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_867),
.B(n_661),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_789),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_919),
.A2(n_494),
.B1(n_922),
.B2(n_624),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_808),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_789),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_894),
.B(n_736),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_919),
.A2(n_494),
.B1(n_922),
.B2(n_624),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_911),
.B(n_742),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_808),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_919),
.A2(n_922),
.B(n_898),
.C(n_709),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_886),
.A2(n_742),
.B1(n_492),
.B2(n_545),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_894),
.B(n_736),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_789),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1050),
.A2(n_1084),
.B(n_1085),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1111),
.A2(n_1115),
.B(n_1038),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_987),
.A2(n_1105),
.B(n_1103),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1117),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_972),
.A2(n_1078),
.B(n_1088),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_R g1129 ( 
.A(n_1002),
.B(n_1034),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_974),
.B(n_1112),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1106),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1060),
.B(n_1080),
.Y(n_1132)
);

AOI221x1_ASAP7_75t_L g1133 ( 
.A1(n_1107),
.A2(n_1023),
.B1(n_1014),
.B2(n_1065),
.C(n_1111),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1025),
.A2(n_1016),
.B(n_1015),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1114),
.B(n_1120),
.Y(n_1135)
);

BUFx2_ASAP7_75t_SL g1136 ( 
.A(n_991),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_998),
.B(n_974),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1013),
.B(n_1100),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1116),
.B(n_994),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1007),
.B(n_980),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_973),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_1012),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1032),
.B(n_997),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1052),
.A2(n_1056),
.A3(n_1001),
.B(n_1115),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1074),
.A2(n_1095),
.B1(n_1008),
.B2(n_1109),
.Y(n_1145)
);

BUFx8_ASAP7_75t_L g1146 ( 
.A(n_1022),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1078),
.A2(n_1058),
.B(n_1052),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_982),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1095),
.A2(n_978),
.B1(n_1010),
.B2(n_1011),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1058),
.A2(n_1056),
.B(n_1018),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1092),
.A2(n_1004),
.B(n_1019),
.C(n_1069),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1079),
.A2(n_1091),
.B(n_1088),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1091),
.A2(n_985),
.B(n_983),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1059),
.A2(n_1076),
.A3(n_1071),
.B(n_1077),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1020),
.Y(n_1155)
);

AOI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_976),
.A2(n_1121),
.B1(n_1101),
.B2(n_999),
.C(n_1110),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_983),
.A2(n_985),
.B(n_1017),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1118),
.A2(n_1062),
.B(n_1057),
.C(n_996),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_990),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_988),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1070),
.A2(n_984),
.B(n_1113),
.C(n_1009),
.Y(n_1161)
);

OAI211xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1041),
.A2(n_1053),
.B(n_1046),
.C(n_1031),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1036),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1081),
.A2(n_1040),
.B(n_1028),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_993),
.B(n_989),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1087),
.A2(n_1073),
.A3(n_1042),
.B(n_1043),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1006),
.A2(n_1099),
.B1(n_1102),
.B2(n_1027),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1045),
.B(n_1099),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1024),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1102),
.A2(n_1027),
.B1(n_1086),
.B2(n_1054),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_977),
.A2(n_1104),
.B(n_1048),
.C(n_1055),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1033),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_L g1173 ( 
.A(n_992),
.B(n_979),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1082),
.A2(n_1061),
.B(n_977),
.C(n_975),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1109),
.A2(n_1090),
.B(n_1026),
.C(n_1097),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1000),
.A2(n_1047),
.B(n_1037),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_979),
.A2(n_1072),
.B(n_992),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1044),
.A2(n_1047),
.B(n_1003),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1066),
.A2(n_1049),
.B(n_1030),
.C(n_1026),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1039),
.Y(n_1180)
);

AO32x2_ASAP7_75t_L g1181 ( 
.A1(n_1064),
.A2(n_986),
.A3(n_1021),
.B1(n_1035),
.B2(n_1093),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1093),
.B(n_1109),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_1030),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1066),
.A2(n_1097),
.B(n_1044),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1051),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_990),
.B(n_981),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1067),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1005),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_995),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1067),
.A2(n_979),
.B(n_995),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_995),
.A2(n_1029),
.B(n_1096),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1108),
.A2(n_1005),
.B1(n_1029),
.B2(n_1096),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1029),
.B(n_1096),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1108),
.A2(n_1038),
.B(n_1075),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1107),
.A2(n_742),
.B1(n_483),
.B2(n_1023),
.C(n_416),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1107),
.A2(n_1023),
.B1(n_994),
.B2(n_1098),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_974),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1107),
.A2(n_1023),
.B1(n_994),
.B2(n_1098),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_973),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1060),
.B(n_1080),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1034),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_973),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_1102),
.B(n_828),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1038),
.A2(n_1016),
.B(n_822),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1107),
.A2(n_496),
.B(n_736),
.C(n_753),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_1023),
.A2(n_1056),
.A3(n_1052),
.B1(n_1115),
.B2(n_1111),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1098),
.A2(n_1119),
.B1(n_584),
.B2(n_406),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1065),
.A2(n_1050),
.B(n_1078),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_973),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_994),
.A2(n_1011),
.B(n_1023),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1038),
.A2(n_1016),
.B(n_822),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_973),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1107),
.A2(n_1023),
.B1(n_994),
.B2(n_1098),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1107),
.B(n_1032),
.C(n_978),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1034),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_973),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1021),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_994),
.A2(n_1032),
.B1(n_1023),
.B2(n_1038),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1021),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1034),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1034),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1060),
.B(n_1080),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1114),
.B(n_1120),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_994),
.A2(n_1032),
.B1(n_1023),
.B2(n_1038),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1032),
.A2(n_1011),
.B(n_1092),
.C(n_1107),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_973),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1075),
.A2(n_1065),
.B(n_1060),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1098),
.B(n_742),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1107),
.A2(n_496),
.B(n_736),
.C(n_753),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1107),
.B(n_1032),
.C(n_978),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1034),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1093),
.B(n_1099),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1060),
.B(n_1080),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_973),
.Y(n_1251)
);

BUFx2_ASAP7_75t_R g1252 ( 
.A(n_1002),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1021),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1098),
.B(n_742),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1060),
.B(n_1080),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1107),
.A2(n_496),
.B(n_736),
.C(n_753),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1260)
);

AO32x2_ASAP7_75t_L g1261 ( 
.A1(n_1023),
.A2(n_1056),
.A3(n_1052),
.B1(n_1115),
.B2(n_1111),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1089),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1021),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1264)
);

OAI22x1_ASAP7_75t_L g1265 ( 
.A1(n_1098),
.A2(n_1119),
.B1(n_742),
.B2(n_1032),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_973),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1038),
.A2(n_965),
.B(n_1120),
.C(n_1114),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1098),
.B(n_1119),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1038),
.A2(n_1075),
.B(n_1025),
.Y(n_1269)
);

AOI31xp67_ASAP7_75t_L g1270 ( 
.A1(n_1075),
.A2(n_1063),
.A3(n_1083),
.B(n_1080),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1141),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1142),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1198),
.A2(n_1202),
.B1(n_1223),
.B2(n_1195),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1203),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1207),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1209),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1230),
.B(n_1237),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1230),
.A2(n_1237),
.B1(n_1226),
.B2(n_1205),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1232),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1233),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1146),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1217),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1198),
.A2(n_1202),
.B1(n_1223),
.B2(n_1215),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1219),
.A2(n_1246),
.B1(n_1224),
.B2(n_1139),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1129),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1155),
.Y(n_1286)
);

INVx6_ASAP7_75t_SL g1287 ( 
.A(n_1248),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1222),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1146),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1219),
.A2(n_1246),
.B1(n_1224),
.B2(n_1265),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1247),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1123),
.A2(n_1268),
.B1(n_1256),
.B2(n_1259),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1140),
.B(n_1130),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1227),
.Y(n_1294)
);

BUFx8_ASAP7_75t_SL g1295 ( 
.A(n_1225),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1204),
.A2(n_1250),
.B1(n_1243),
.B2(n_1255),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1163),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1145),
.A2(n_1167),
.B1(n_1165),
.B2(n_1170),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1240),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1138),
.A2(n_1143),
.B1(n_1167),
.B2(n_1149),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1125),
.A2(n_1239),
.B1(n_1236),
.B2(n_1151),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1150),
.A2(n_1149),
.B(n_1213),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1252),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_1170),
.B1(n_1137),
.B2(n_1180),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1251),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_1135),
.B1(n_1176),
.B2(n_1187),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1176),
.A2(n_1194),
.B1(n_1211),
.B2(n_1172),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1266),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1131),
.A2(n_1211),
.B1(n_1182),
.B2(n_1127),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1148),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1193),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1212),
.A2(n_1221),
.B1(n_1261),
.B2(n_1214),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1188),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1212),
.A2(n_1221),
.B1(n_1214),
.B2(n_1261),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1169),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1185),
.A2(n_1156),
.B1(n_1186),
.B2(n_1157),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1136),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1160),
.B(n_1168),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1147),
.A2(n_1258),
.B1(n_1244),
.B2(n_1214),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1186),
.B(n_1184),
.Y(n_1320)
);

CKINVDCx6p67_ASAP7_75t_R g1321 ( 
.A(n_1192),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1229),
.A2(n_1253),
.B1(n_1231),
.B2(n_1263),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1133),
.A2(n_1183),
.B1(n_1261),
.B2(n_1220),
.Y(n_1323)
);

BUFx5_ASAP7_75t_L g1324 ( 
.A(n_1270),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1181),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1200),
.A2(n_1241),
.B1(n_1228),
.B2(n_1264),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1210),
.A2(n_1269),
.B1(n_1234),
.B2(n_1238),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1191),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1144),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1190),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1153),
.A2(n_1162),
.B1(n_1242),
.B2(n_1263),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1173),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1174),
.A2(n_1134),
.B1(n_1158),
.B2(n_1152),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1181),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1161),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1144),
.A2(n_1267),
.B1(n_1242),
.B2(n_1216),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1144),
.B(n_1166),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1216),
.A2(n_1177),
.B1(n_1164),
.B2(n_1128),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1178),
.A2(n_1126),
.B1(n_1175),
.B2(n_1171),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1179),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1124),
.A2(n_1166),
.B1(n_1154),
.B2(n_1132),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1154),
.A2(n_1257),
.B1(n_1132),
.B2(n_1249),
.Y(n_1343)
);

INVx4_ASAP7_75t_SL g1344 ( 
.A(n_1206),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1122),
.A2(n_1262),
.B1(n_1196),
.B2(n_1197),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1235),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1201),
.A2(n_1208),
.B1(n_1218),
.B2(n_1245),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1254),
.A2(n_1260),
.B1(n_1249),
.B2(n_1257),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1257),
.Y(n_1349)
);

OAI22x1_ASAP7_75t_L g1350 ( 
.A1(n_1198),
.A2(n_1202),
.B1(n_1223),
.B2(n_1170),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1142),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1230),
.B(n_994),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1159),
.B(n_979),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1129),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1141),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1232),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1146),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1098),
.Y(n_1359)
);

BUFx4_ASAP7_75t_R g1360 ( 
.A(n_1148),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1141),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1098),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1232),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1198),
.A2(n_742),
.B1(n_1223),
.B2(n_1202),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1142),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_1223),
.B(n_1202),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1230),
.A2(n_1237),
.B(n_1224),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1230),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1230),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1141),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1141),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1141),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1129),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1230),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1379)
);

AOI21xp33_ASAP7_75t_L g1380 ( 
.A1(n_1230),
.A2(n_1237),
.B(n_1011),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1129),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1230),
.B(n_994),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1230),
.A2(n_1100),
.B1(n_633),
.B2(n_1107),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1098),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1198),
.A2(n_1223),
.B1(n_1202),
.B2(n_1230),
.Y(n_1385)
);

CKINVDCx6p67_ASAP7_75t_R g1386 ( 
.A(n_1207),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1146),
.Y(n_1387)
);

NOR2x1_ASAP7_75t_SL g1388 ( 
.A(n_1230),
.B(n_1237),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1329),
.Y(n_1389)
);

AO21x1_ASAP7_75t_L g1390 ( 
.A1(n_1368),
.A2(n_1378),
.B(n_1370),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1346),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1318),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1338),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1330),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1367),
.A2(n_1370),
.B(n_1368),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1323),
.A2(n_1367),
.B(n_1378),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1349),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1312),
.B(n_1314),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1297),
.B(n_1296),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1324),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1325),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1331),
.B(n_1344),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1271),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1274),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1276),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1312),
.B(n_1314),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1282),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1288),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1324),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1294),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1348),
.A2(n_1302),
.B(n_1339),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1345),
.A2(n_1347),
.B(n_1334),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1331),
.B(n_1388),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1278),
.B(n_1299),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1305),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1351),
.A2(n_1371),
.B1(n_1377),
.B2(n_1379),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1308),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1385),
.A2(n_1277),
.B(n_1380),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1326),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1278),
.B(n_1315),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1385),
.B(n_1293),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1292),
.B(n_1366),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1273),
.A2(n_1364),
.B1(n_1283),
.B2(n_1372),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1311),
.B(n_1353),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1356),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1290),
.B(n_1284),
.C(n_1301),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1361),
.B(n_1373),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1324),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1324),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1374),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1375),
.B(n_1350),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1343),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1333),
.B(n_1298),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1320),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1334),
.A2(n_1332),
.B(n_1340),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1319),
.A2(n_1307),
.B(n_1336),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1343),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1313),
.B(n_1310),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1337),
.B(n_1380),
.Y(n_1440)
);

NAND2x1_ASAP7_75t_L g1441 ( 
.A(n_1341),
.B(n_1319),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1306),
.A2(n_1382),
.B(n_1300),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1342),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1337),
.B(n_1301),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1328),
.Y(n_1445)
);

CKINVDCx6p67_ASAP7_75t_R g1446 ( 
.A(n_1352),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1382),
.B(n_1362),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1335),
.Y(n_1448)
);

CKINVDCx10_ASAP7_75t_R g1449 ( 
.A(n_1360),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1359),
.A2(n_1384),
.B(n_1309),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1327),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1316),
.A2(n_1304),
.B(n_1354),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1341),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1322),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1369),
.A2(n_1383),
.B(n_1333),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1321),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1326),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1287),
.A2(n_1387),
.B1(n_1358),
.B2(n_1289),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1357),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1291),
.A2(n_1272),
.B(n_1381),
.C(n_1376),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1279),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1279),
.B(n_1387),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1317),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1405),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1423),
.A2(n_1285),
.B(n_1358),
.C(n_1281),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1444),
.B(n_1281),
.Y(n_1467)
);

INVx11_ASAP7_75t_L g1468 ( 
.A(n_1449),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1435),
.B(n_1355),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1460),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1392),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1426),
.A2(n_1303),
.B(n_1295),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1412),
.A2(n_1363),
.B(n_1289),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1437),
.A2(n_1365),
.B(n_1289),
.Y(n_1474)
);

AO32x2_ASAP7_75t_L g1475 ( 
.A1(n_1389),
.A2(n_1281),
.A3(n_1358),
.B1(n_1275),
.B2(n_1386),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1280),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1421),
.B(n_1286),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1399),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1414),
.B(n_1286),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1444),
.B(n_1427),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1407),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1395),
.A2(n_1426),
.B1(n_1416),
.B2(n_1423),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1395),
.A2(n_1418),
.B(n_1447),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_1447),
.B(n_1440),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1427),
.B(n_1403),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1410),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1440),
.A2(n_1451),
.B(n_1453),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1390),
.A2(n_1450),
.B1(n_1456),
.B2(n_1396),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1390),
.A2(n_1422),
.B(n_1456),
.C(n_1450),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1408),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1428),
.A2(n_1429),
.B(n_1430),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1441),
.A2(n_1422),
.B(n_1398),
.C(n_1406),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1451),
.A2(n_1453),
.B(n_1441),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1439),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1436),
.A2(n_1414),
.B(n_1420),
.C(n_1452),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1415),
.B(n_1417),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1446),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1402),
.B(n_1413),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1450),
.A2(n_1396),
.B1(n_1420),
.B2(n_1432),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1432),
.B(n_1396),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1396),
.B(n_1425),
.Y(n_1503)
);

INVx5_ASAP7_75t_L g1504 ( 
.A(n_1454),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1431),
.B(n_1411),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1436),
.A2(n_1452),
.B(n_1401),
.C(n_1455),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1434),
.A2(n_1445),
.B(n_1459),
.C(n_1458),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1452),
.A2(n_1401),
.B(n_1443),
.C(n_1438),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1433),
.A2(n_1438),
.B(n_1445),
.C(n_1448),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1411),
.B(n_1433),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1446),
.B(n_1461),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1391),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1485),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1503),
.B(n_1394),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1481),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1513),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1505),
.B(n_1400),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1491),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1505),
.B(n_1394),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1492),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1502),
.B(n_1412),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1511),
.B(n_1409),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1511),
.B(n_1409),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1483),
.B(n_1397),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1489),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1498),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1504),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1397),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1526),
.B(n_1516),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1518),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1515),
.B(n_1524),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1527),
.A2(n_1482),
.B1(n_1488),
.B2(n_1501),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1515),
.B(n_1510),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1526),
.B(n_1465),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1518),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1518),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1522),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1515),
.B(n_1497),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1515),
.B(n_1497),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1523),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1473),
.Y(n_1548)
);

OAI211xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1526),
.A2(n_1472),
.B(n_1490),
.C(n_1470),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1486),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1471),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1522),
.A2(n_1508),
.B(n_1506),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1527),
.A2(n_1442),
.B1(n_1487),
.B2(n_1478),
.Y(n_1553)
);

NAND4xp75_ASAP7_75t_L g1554 ( 
.A(n_1532),
.B(n_1457),
.C(n_1495),
.D(n_1476),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1517),
.B(n_1479),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1530),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1500),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1519),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1530),
.Y(n_1559)
);

AOI211xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1523),
.A2(n_1512),
.B(n_1499),
.C(n_1494),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.B(n_1473),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1534),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1543),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1534),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1543),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1534),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1557),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1517),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1544),
.B(n_1527),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1521),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1546),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1540),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1519),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1543),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1556),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1547),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1546),
.B(n_1519),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1519),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1499),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1535),
.B(n_1528),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1529),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1529),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.B(n_1529),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1537),
.B(n_1529),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1539),
.B(n_1529),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1549),
.A2(n_1536),
.B1(n_1532),
.B2(n_1553),
.C(n_1494),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1542),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1545),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1590),
.A2(n_1536),
.B1(n_1554),
.B2(n_1553),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1590),
.A2(n_1554),
.B1(n_1552),
.B2(n_1474),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_SL g1596 ( 
.A(n_1582),
.B(n_1572),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1562),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1572),
.B(n_1565),
.Y(n_1598)
);

NAND4xp25_ASAP7_75t_L g1599 ( 
.A(n_1582),
.B(n_1560),
.C(n_1555),
.D(n_1556),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.B(n_1556),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1565),
.B(n_1559),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1559),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1578),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1570),
.B(n_1559),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1564),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1559),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1570),
.B(n_1558),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1576),
.A2(n_1554),
.B1(n_1552),
.B2(n_1474),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1558),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1576),
.B(n_1580),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1551),
.Y(n_1617)
);

NAND4xp25_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1560),
.C(n_1555),
.D(n_1466),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.B(n_1584),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1567),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1558),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1580),
.B(n_1557),
.Y(n_1623)
);

OAI321xp33_ASAP7_75t_L g1624 ( 
.A1(n_1579),
.A2(n_1508),
.A3(n_1523),
.B1(n_1509),
.B2(n_1506),
.C(n_1532),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1591),
.B(n_1557),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1573),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1573),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1557),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1591),
.B(n_1557),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1571),
.B(n_1551),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1632)
);

NAND2x1_ASAP7_75t_L g1633 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1574),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1598),
.B(n_1584),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1616),
.B(n_1578),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1616),
.B(n_1600),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1631),
.B(n_1584),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1597),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1594),
.B(n_1587),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1587),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1581),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1589),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1620),
.B(n_1589),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1468),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1583),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1604),
.B(n_1583),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1607),
.B(n_1531),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1619),
.B(n_1569),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1602),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1596),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1595),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1585),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

NAND2x1_ASAP7_75t_SL g1664 ( 
.A(n_1613),
.B(n_1568),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1619),
.B(n_1603),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1599),
.B(n_1568),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1610),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1614),
.B(n_1568),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1614),
.B(n_1568),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1660),
.A2(n_1552),
.B1(n_1523),
.B2(n_1548),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1644),
.A2(n_1552),
.B1(n_1548),
.B2(n_1561),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1650),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1669),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1639),
.B(n_1632),
.Y(n_1680)
);

AND3x2_ASAP7_75t_L g1681 ( 
.A(n_1638),
.B(n_1467),
.C(n_1607),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1641),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1643),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1665),
.B(n_1638),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1646),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1638),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1637),
.A2(n_1624),
.B1(n_1596),
.B2(n_1601),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1655),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1656),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1663),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1670),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1601),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1636),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1653),
.B(n_1623),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1664),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1673),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1687),
.A2(n_1668),
.B1(n_1552),
.B2(n_1651),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1654),
.Y(n_1700)
);

AOI32xp33_ASAP7_75t_L g1701 ( 
.A1(n_1697),
.A2(n_1642),
.A3(n_1640),
.B1(n_1648),
.B2(n_1649),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1684),
.Y(n_1702)
);

OAI32xp33_ASAP7_75t_L g1703 ( 
.A1(n_1695),
.A2(n_1653),
.A3(n_1637),
.B1(n_1642),
.B2(n_1648),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1686),
.B(n_1647),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1688),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1688),
.Y(n_1706)
);

O2A1O1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1677),
.A2(n_1649),
.B(n_1569),
.C(n_1640),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1686),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1694),
.B(n_1684),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1678),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1677),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1675),
.A2(n_1461),
.B(n_1603),
.C(n_1645),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1682),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1679),
.A2(n_1652),
.B1(n_1662),
.B2(n_1657),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1683),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1689),
.B(n_1615),
.C(n_1610),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_R g1717 ( 
.A(n_1710),
.B(n_1672),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1716),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1709),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1712),
.A2(n_1690),
.B(n_1685),
.C(n_1672),
.Y(n_1720)
);

XNOR2x2_ASAP7_75t_SL g1721 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1698),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1704),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1704),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1700),
.B(n_1691),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1711),
.B(n_1692),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1705),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1718),
.B(n_1706),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1724),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1718),
.A2(n_1701),
.B(n_1708),
.C(n_1707),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1719),
.A2(n_1721),
.B1(n_1726),
.B2(n_1725),
.Y(n_1731)
);

NOR3x1_ASAP7_75t_L g1732 ( 
.A(n_1726),
.B(n_1715),
.C(n_1713),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1720),
.A2(n_1703),
.B1(n_1702),
.B2(n_1693),
.C(n_1714),
.Y(n_1733)
);

AOI211x1_ASAP7_75t_L g1734 ( 
.A1(n_1722),
.A2(n_1696),
.B(n_1716),
.C(n_1680),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1735)
);

XNOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1727),
.B(n_1681),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1717),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1734),
.A2(n_1731),
.B1(n_1728),
.B2(n_1735),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1730),
.A2(n_1696),
.B1(n_1577),
.B2(n_1566),
.C(n_1563),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1737),
.B(n_1647),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1733),
.A2(n_1671),
.B1(n_1670),
.B2(n_1627),
.C(n_1635),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1729),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1736),
.A2(n_1566),
.B1(n_1563),
.B2(n_1577),
.C(n_1615),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1738),
.A2(n_1732),
.B(n_1633),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1740),
.A2(n_1633),
.B(n_1626),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1743),
.A2(n_1627),
.B(n_1635),
.C(n_1605),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1741),
.A2(n_1671),
.B(n_1659),
.C(n_1667),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1659),
.B1(n_1605),
.B2(n_1623),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_SL g1749 ( 
.A1(n_1739),
.A2(n_1496),
.B(n_1634),
.C(n_1628),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1738),
.A2(n_1634),
.B(n_1621),
.C(n_1626),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1748),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1750),
.B(n_1621),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1749),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1747),
.B(n_1625),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1746),
.Y(n_1755)
);

AOI221x1_ASAP7_75t_L g1756 ( 
.A1(n_1751),
.A2(n_1744),
.B1(n_1745),
.B2(n_1628),
.C(n_1574),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1755),
.B(n_1566),
.C(n_1563),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1753),
.B(n_1577),
.C(n_1507),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1754),
.Y(n_1759)
);

OAI22x1_ASAP7_75t_L g1760 ( 
.A1(n_1759),
.A2(n_1752),
.B1(n_1757),
.B2(n_1756),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1760),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1760),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1761),
.B(n_1752),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1762),
.A2(n_1419),
.B1(n_1477),
.B2(n_1469),
.Y(n_1764)
);

AOI21xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1763),
.A2(n_1469),
.B(n_1625),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1630),
.B(n_1629),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1765),
.A2(n_1630),
.B(n_1629),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1767),
.B(n_1766),
.Y(n_1768)
);

AO22x2_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1458),
.B1(n_1593),
.B2(n_1592),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1463),
.B1(n_1593),
.B2(n_1592),
.C(n_1575),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1469),
.B(n_1467),
.C(n_1462),
.Y(n_1771)
);


endmodule