module fake_jpeg_27150_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_21),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_17),
.B1(n_29),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_56),
.B1(n_26),
.B2(n_19),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_20),
.B2(n_30),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_54),
.B(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_17),
.B1(n_30),
.B2(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_31),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_19),
.B1(n_23),
.B2(n_32),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_32),
.B1(n_33),
.B2(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_80),
.B1(n_81),
.B2(n_12),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_35),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_84),
.B(n_4),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_73),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_11),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_32),
.B1(n_23),
.B2(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_94),
.B1(n_98),
.B2(n_11),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_34),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_33),
.B(n_18),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_6),
.B(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_16),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_27),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_2),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_33),
.B1(n_18),
.B2(n_4),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_33),
.B1(n_18),
.B2(n_4),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_2),
.B(n_3),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_9),
.C(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_5),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_94),
.B(n_84),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_5),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_120),
.C(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_108),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_13),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_9),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_10),
.C(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_10),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_129),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_126),
.B1(n_78),
.B2(n_77),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_136),
.B1(n_156),
.B2(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_146),
.B(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_119),
.B(n_98),
.Y(n_187)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_84),
.C(n_79),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_87),
.C(n_89),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_69),
.B1(n_81),
.B2(n_71),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_81),
.B1(n_72),
.B2(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_72),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_87),
.Y(n_161)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_176),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_110),
.B(n_107),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_168),
.B(n_190),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_110),
.B(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_108),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_154),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_123),
.B1(n_126),
.B2(n_115),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_178),
.B1(n_169),
.B2(n_133),
.Y(n_191)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_126),
.B1(n_115),
.B2(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_120),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_184),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_128),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_104),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_182),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_130),
.B(n_119),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_212),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_196),
.Y(n_219)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_145),
.B1(n_156),
.B2(n_158),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_202),
.B1(n_210),
.B2(n_190),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_185),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_154),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_138),
.B1(n_157),
.B2(n_150),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_104),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_134),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_171),
.B(n_101),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_124),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_170),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_189),
.C(n_163),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_218),
.C(n_225),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_224),
.B1(n_231),
.B2(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_179),
.C(n_166),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_167),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_228),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_174),
.B1(n_178),
.B2(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_166),
.C(n_168),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_194),
.C(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_208),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_196),
.A2(n_181),
.B1(n_186),
.B2(n_124),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_181),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_238),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_201),
.B1(n_204),
.B2(n_211),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_220),
.B1(n_197),
.B2(n_223),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_241),
.B1(n_242),
.B2(n_250),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_246),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_245),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_230),
.B1(n_203),
.B2(n_201),
.Y(n_241)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_225),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_250),
.B(n_221),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_206),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_216),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

BUFx12f_ASAP7_75t_SL g250 ( 
.A(n_229),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_261),
.B1(n_239),
.B2(n_198),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_262),
.B(n_175),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_164),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_218),
.C(n_197),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_205),
.B(n_176),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_246),
.B(n_241),
.C(n_244),
.D(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_193),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_272),
.B1(n_87),
.B2(n_82),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_175),
.B1(n_87),
.B2(n_90),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_255),
.B1(n_259),
.B2(n_96),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_14),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_13),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_256),
.B(n_101),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_273),
.B(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_268),
.C(n_265),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_279),
.A3(n_276),
.B1(n_280),
.B2(n_275),
.C1(n_96),
.C2(n_15),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_286),
.B(n_15),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_289),
.B(n_282),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_287),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_291),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_15),
.Y(n_294)
);


endmodule