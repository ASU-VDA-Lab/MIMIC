module fake_netlist_1_1385_n_883 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_883);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_883;
wire n_117;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_704;
wire n_611;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_703;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_649;
wire n_526;
wire n_276;
wire n_527;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_822;
wire n_823;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_695;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g104 ( .A(n_17), .Y(n_104) );
BUFx10_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_60), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_75), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_28), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_87), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_45), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_26), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_15), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_22), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_6), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_41), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_91), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_16), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_14), .Y(n_131) );
INVxp33_ASAP7_75t_L g132 ( .A(n_50), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_19), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_30), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_37), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_12), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_58), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_21), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_32), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_111), .B(n_0), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_125), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_125), .B(n_1), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_111), .B(n_3), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_113), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_110), .A2(n_51), .B(n_101), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_110), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_107), .B(n_4), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_123), .B(n_5), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_112), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_116), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_105), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_105), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_116), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_132), .B(n_5), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_120), .B(n_24), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_129), .B(n_6), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_127), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_155), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_161), .B(n_138), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
XNOR2xp5_ASAP7_75t_L g173 ( .A(n_145), .B(n_135), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
BUFx10_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_161), .B(n_142), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_161), .B(n_140), .Y(n_180) );
INVxp33_ASAP7_75t_SL g181 ( .A(n_159), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_160), .B(n_105), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_146), .B(n_107), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_161), .B(n_109), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_146), .A2(n_118), .B1(n_124), .B2(n_104), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_160), .B(n_127), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_145), .A2(n_108), .B1(n_117), .B2(n_128), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_160), .B(n_105), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_160), .B(n_108), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_147), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_158), .B(n_117), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_154), .A2(n_141), .B(n_133), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_146), .A2(n_128), .B1(n_130), .B2(n_122), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_148), .A2(n_130), .B1(n_133), .B2(n_134), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_166), .B(n_114), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_159), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_158), .B(n_134), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_144), .B(n_136), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_171), .B(n_148), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_183), .A2(n_148), .B1(n_143), .B2(n_166), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_180), .B(n_164), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_201), .B(n_164), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_192), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_198), .B(n_165), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_198), .B(n_164), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_211), .B(n_143), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_183), .B(n_166), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_183), .A2(n_167), .B1(n_157), .B2(n_156), .Y(n_228) );
INVx5_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_201), .B(n_144), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_191), .B(n_154), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_201), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_200), .B(n_150), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_192), .Y(n_235) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_198), .B(n_151), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g237 ( .A(n_212), .B(n_139), .C(n_119), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_214), .B(n_150), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_198), .B(n_152), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_194), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_213), .B(n_152), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_214), .B(n_153), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_183), .B(n_153), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_183), .A2(n_167), .B1(n_157), .B2(n_156), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_195), .B(n_115), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_209), .A2(n_141), .B1(n_136), .B2(n_137), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_195), .B(n_121), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_206), .B(n_126), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_196), .A2(n_151), .B1(n_8), .B2(n_9), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_194), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_206), .B(n_7), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_181), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_199), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_186), .B(n_7), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_215), .B(n_213), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_54), .B(n_100), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_186), .B(n_9), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_202), .Y(n_259) );
BUFx8_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_168), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_191), .B(n_10), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_196), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_213), .B(n_59), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_215), .A2(n_213), .B1(n_208), .B2(n_168), .Y(n_265) );
INVxp33_ASAP7_75t_L g266 ( .A(n_173), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_188), .B(n_57), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_168), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_186), .B(n_11), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_178), .A2(n_65), .B(n_98), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_170), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_223), .A2(n_175), .B(n_177), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_238), .B(n_215), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_260), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_223), .A2(n_175), .B(n_177), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_229), .Y(n_277) );
INVx6_ASAP7_75t_L g278 ( .A(n_260), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_267), .A2(n_215), .B(n_170), .C(n_175), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_242), .B(n_210), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_227), .B(n_173), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_243), .B(n_208), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_217), .B(n_208), .Y(n_284) );
AOI22x1_ASAP7_75t_L g285 ( .A1(n_270), .A2(n_185), .B1(n_193), .B2(n_197), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_234), .A2(n_175), .B(n_177), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_229), .B(n_176), .Y(n_287) );
OAI321xp33_ASAP7_75t_L g288 ( .A1(n_249), .A2(n_216), .A3(n_204), .B1(n_207), .B2(n_205), .C(n_190), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_227), .B(n_229), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_225), .A2(n_170), .B(n_177), .C(n_204), .Y(n_290) );
OR2x6_ASAP7_75t_SL g291 ( .A(n_252), .B(n_190), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_233), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_256), .B(n_176), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_231), .B(n_208), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_262), .A2(n_170), .B1(n_176), .B2(n_203), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_241), .A2(n_189), .B(n_169), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_225), .B(n_185), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_239), .A2(n_185), .B(n_197), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_228), .A2(n_185), .B1(n_193), .B2(n_197), .Y(n_299) );
OA22x2_ASAP7_75t_L g300 ( .A1(n_227), .A2(n_207), .B1(n_205), .B2(n_203), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_239), .A2(n_185), .B(n_197), .Y(n_301) );
NAND2xp33_ASAP7_75t_L g302 ( .A(n_265), .B(n_193), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_230), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_241), .A2(n_197), .B(n_193), .Y(n_304) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_237), .B(n_251), .Y(n_305) );
AOI22x1_ASAP7_75t_L g306 ( .A1(n_257), .A2(n_197), .B1(n_193), .B2(n_203), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_244), .A2(n_193), .B1(n_205), .B2(n_207), .Y(n_307) );
BUFx12f_ASAP7_75t_L g308 ( .A(n_256), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_219), .A2(n_190), .B(n_179), .C(n_184), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_224), .B(n_13), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_220), .B(n_13), .Y(n_311) );
OR2x6_ASAP7_75t_SL g312 ( .A(n_218), .B(n_14), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_256), .A2(n_187), .B1(n_169), .B2(n_184), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_274), .A2(n_265), .B1(n_253), .B2(n_222), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
AOI21x1_ASAP7_75t_L g316 ( .A1(n_299), .A2(n_264), .B(n_269), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_304), .A2(n_226), .B(n_224), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_280), .B(n_248), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_281), .B(n_266), .Y(n_321) );
AOI221x1_ASAP7_75t_L g322 ( .A1(n_290), .A2(n_258), .B1(n_255), .B2(n_226), .C(n_267), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_302), .A2(n_226), .B(n_236), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_298), .A2(n_226), .B(n_236), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_290), .A2(n_246), .B(n_247), .C(n_245), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_275), .B(n_294), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_280), .A2(n_240), .B(n_254), .C(n_250), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_284), .A2(n_222), .B(n_235), .C(n_253), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_310), .A2(n_263), .B1(n_221), .B2(n_268), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_271), .B(n_268), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_271), .B(n_261), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_SL g332 ( .A1(n_309), .A2(n_264), .B(n_172), .C(n_174), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_297), .A2(n_261), .B(n_259), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_292), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_283), .A2(n_235), .B(n_221), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_303), .B(n_15), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_16), .Y(n_337) );
AOI221x1_ASAP7_75t_L g338 ( .A1(n_307), .A2(n_179), .B1(n_174), .B2(n_172), .C(n_187), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_306), .A2(n_187), .B(n_169), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_312), .B(n_17), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_326), .B(n_289), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_316), .A2(n_285), .B(n_279), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_323), .A2(n_296), .B(n_276), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_320), .B(n_295), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_332), .A2(n_324), .B(n_317), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_322), .B(n_310), .C(n_305), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_318), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_319), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_334), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_320), .B(n_286), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_319), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_339), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_341), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_328), .B(n_272), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_311), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_338), .A2(n_288), .B(n_273), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_330), .A2(n_300), .B(n_313), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_327), .A2(n_300), .B(n_313), .Y(n_364) );
NOR2x1_ASAP7_75t_SL g365 ( .A(n_314), .B(n_337), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_321), .A2(n_278), .B1(n_308), .B2(n_293), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_327), .A2(n_287), .B(n_293), .Y(n_367) );
AO31x2_ASAP7_75t_L g368 ( .A1(n_335), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_368) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_336), .B(n_278), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_325), .A2(n_333), .B(n_329), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_351), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_351), .Y(n_373) );
AOI33xp33_ASAP7_75t_L g374 ( .A1(n_353), .A2(n_332), .A3(n_21), .B1(n_22), .B2(n_23), .B3(n_18), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_357), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_287), .B(n_277), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_189), .B(n_25), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_277), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_345), .A2(n_272), .B(n_189), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_23), .B(n_189), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_345), .A2(n_27), .B(n_29), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_345), .A2(n_31), .B(n_33), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_359), .B(n_103), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_368), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_347), .B(n_34), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_35), .Y(n_387) );
AND2x4_ASAP7_75t_SL g388 ( .A(n_343), .B(n_36), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_368), .B(n_38), .Y(n_391) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_352), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_359), .B(n_39), .Y(n_393) );
CKINVDCx11_ASAP7_75t_R g394 ( .A(n_355), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_370), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_368), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_368), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_368), .B(n_40), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_347), .B(n_43), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
AO21x2_ASAP7_75t_L g403 ( .A1(n_349), .A2(n_44), .B(n_46), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_343), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_354), .B(n_47), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_343), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_344), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_49), .B(n_52), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_342), .B(n_53), .Y(n_410) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_370), .B(n_66), .Y(n_411) );
INVxp33_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_344), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_354), .B(n_67), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_365), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_350), .B(n_68), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_365), .A2(n_69), .B(n_70), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_372), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_410), .A2(n_358), .B1(n_356), .B2(n_364), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_418), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_367), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_382), .B(n_366), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_418), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_374), .B(n_350), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_373), .B(n_367), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_418), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g432 ( .A(n_384), .B(n_364), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_382), .B(n_367), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_380), .A2(n_362), .B(n_371), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_385), .B(n_367), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_412), .A2(n_369), .B1(n_360), .B2(n_371), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_389), .B(n_350), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_395), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_385), .B(n_360), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_396), .B(n_363), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_396), .B(n_363), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_398), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_363), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_410), .B(n_369), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_410), .B(n_346), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_401), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_378), .B(n_361), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_389), .B(n_361), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_390), .B(n_362), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_399), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_402), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_390), .B(n_346), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_409), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_375), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_391), .B(n_361), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_375), .B(n_361), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_375), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_397), .B(n_361), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_379), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_379), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_391), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_399), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_399), .B(n_346), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_379), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_378), .B(n_71), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_378), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_374), .B(n_96), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_392), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_377), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_416), .A2(n_72), .B(n_73), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_404), .B(n_74), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_387), .B(n_76), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_404), .B(n_77), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_407), .Y(n_481) );
NOR2x1p5_ASAP7_75t_L g482 ( .A(n_416), .B(n_78), .Y(n_482) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_380), .A2(n_79), .B(n_81), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_397), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_407), .B(n_82), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_377), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_387), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_413), .B(n_83), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_406), .B(n_84), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_406), .B(n_85), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_413), .B(n_86), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_384), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_411), .A2(n_88), .B(n_89), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_411), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_384), .B(n_90), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_415), .B(n_92), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_380), .A2(n_93), .B(n_94), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_377), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_417), .B(n_95), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_386), .B(n_400), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_454), .B(n_393), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_492), .B(n_393), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_467), .B(n_400), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_454), .B(n_393), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_482), .B(n_393), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_495), .B(n_387), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_421), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_467), .B(n_400), .Y(n_513) );
NOR2xp67_ASAP7_75t_SL g514 ( .A(n_489), .B(n_386), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_440), .B(n_393), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_468), .B(n_386), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_425), .B(n_384), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_494), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_458), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_440), .B(n_384), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_423), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_469), .B(n_380), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_468), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_433), .B(n_408), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_494), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_433), .B(n_408), .Y(n_526) );
OR2x6_ASAP7_75t_L g527 ( .A(n_492), .B(n_376), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_494), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_443), .B(n_408), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_458), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_443), .B(n_377), .Y(n_531) );
INVxp33_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_463), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_445), .B(n_377), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_427), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_427), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_472), .B(n_414), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_445), .B(n_403), .Y(n_539) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_432), .B(n_388), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_435), .B(n_403), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_463), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_478), .B(n_394), .Y(n_543) );
AND2x4_ASAP7_75t_SL g544 ( .A(n_495), .B(n_419), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_474), .B(n_419), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_435), .B(n_403), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_463), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_423), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_423), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_424), .B(n_403), .Y(n_550) );
CKINVDCx14_ASAP7_75t_R g551 ( .A(n_495), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_424), .B(n_405), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_481), .B(n_405), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_496), .B(n_414), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_419), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_498), .B(n_376), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_498), .B(n_502), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_429), .B(n_420), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_502), .B(n_388), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_484), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_444), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_466), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_479), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_426), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_422), .B(n_388), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_429), .B(n_420), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_448), .B(n_420), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_460), .B(n_420), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_460), .B(n_381), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_444), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_487), .B(n_381), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_426), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_447), .B(n_381), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_447), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_450), .B(n_381), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_450), .B(n_437), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_442), .B(n_381), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_455), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_442), .B(n_383), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_455), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_495), .A2(n_383), .B(n_476), .C(n_432), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_457), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_426), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_431), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_457), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_451), .B(n_383), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_459), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_431), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_456), .B(n_383), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_456), .B(n_383), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_456), .B(n_459), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_456), .B(n_431), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_471), .B(n_438), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_478), .B(n_471), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_439), .B(n_461), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_439), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_452), .B(n_449), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_489), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_438), .B(n_453), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_439), .B(n_461), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_452), .B(n_449), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_490), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_441), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_441), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_441), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_446), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_482), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_446), .Y(n_610) );
AND2x4_ASAP7_75t_SL g611 ( .A(n_600), .B(n_438), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_523), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_596), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_543), .A2(n_473), .B(n_428), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_551), .B(n_438), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_506), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_557), .B(n_449), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_523), .B(n_453), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_512), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_515), .B(n_453), .Y(n_620) );
OAI21xp33_ASAP7_75t_SL g621 ( .A1(n_540), .A2(n_501), .B(n_477), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_561), .B(n_461), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_594), .B(n_446), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_535), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_536), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g626 ( .A1(n_510), .A2(n_476), .B(n_462), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_538), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_507), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_571), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_515), .B(n_520), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_575), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_579), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_581), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_520), .B(n_453), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_533), .B(n_464), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_563), .B(n_430), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_583), .B(n_464), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_582), .A2(n_462), .B(n_500), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_596), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_503), .B(n_430), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_542), .B(n_466), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_586), .B(n_430), .Y(n_642) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_609), .B(n_466), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_542), .B(n_466), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
INVx4_ASAP7_75t_L g646 ( .A(n_544), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_503), .B(n_430), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_509), .B(n_436), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_566), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_509), .B(n_436), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_540), .A2(n_499), .B1(n_483), .B2(n_501), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_519), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_592), .B(n_436), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_605), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_592), .B(n_436), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_577), .B(n_434), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_601), .B(n_434), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_560), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_606), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_560), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_547), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_600), .B(n_485), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_530), .B(n_465), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_599), .B(n_485), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_514), .Y(n_665) );
AOI22x1_ASAP7_75t_L g666 ( .A1(n_511), .A2(n_493), .B1(n_497), .B2(n_491), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_598), .B(n_465), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_601), .B(n_434), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_545), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_603), .B(n_497), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_598), .B(n_465), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_600), .B(n_491), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_607), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_593), .B(n_488), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_610), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_597), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_521), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_597), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_604), .B(n_477), .Y(n_680) );
NAND2x1p5_ASAP7_75t_L g681 ( .A(n_504), .B(n_480), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_511), .A2(n_499), .B1(n_483), .B2(n_480), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_552), .B(n_488), .Y(n_683) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_521), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_595), .A2(n_483), .B1(n_499), .B2(n_486), .Y(n_685) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_532), .B(n_470), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_608), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_552), .B(n_475), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_548), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_548), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_602), .B(n_470), .Y(n_692) );
INVx3_ASAP7_75t_SL g693 ( .A(n_504), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_593), .B(n_470), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_602), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_504), .B(n_475), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_559), .B(n_475), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_555), .B(n_486), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_508), .B(n_486), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_508), .B(n_500), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_513), .B(n_500), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_513), .B(n_516), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_549), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_529), .B(n_522), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_532), .B(n_565), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_549), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_564), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_505), .B(n_525), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_516), .B(n_537), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_564), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_522), .B(n_556), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_531), .B(n_534), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_531), .B(n_534), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_529), .B(n_524), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_517), .B(n_584), .Y(n_715) );
OAI22x1_ASAP7_75t_L g716 ( .A1(n_612), .A2(n_505), .B1(n_518), .B2(n_528), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_618), .B(n_524), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_649), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_714), .B(n_526), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_630), .B(n_526), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_712), .B(n_573), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_695), .B(n_591), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_711), .B(n_578), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_693), .B(n_591), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_712), .B(n_589), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_713), .B(n_709), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_658), .B(n_590), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_711), .B(n_578), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_684), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_620), .B(n_590), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_646), .B(n_505), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_616), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g733 ( .A(n_646), .B(n_518), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_619), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_669), .B(n_553), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_634), .B(n_567), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_713), .B(n_589), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_635), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_702), .B(n_585), .Y(n_739) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_621), .B(n_582), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_704), .B(n_567), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_624), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_625), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_627), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_656), .B(n_576), .Y(n_745) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_621), .B(n_527), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_629), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_705), .A2(n_539), .B1(n_546), .B2(n_541), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_631), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_614), .A2(n_568), .B(n_554), .C(n_572), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_708), .B(n_518), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_667), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_652), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_632), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_660), .B(n_525), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_628), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_715), .B(n_573), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_656), .B(n_576), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_640), .B(n_558), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_647), .B(n_558), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_633), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_645), .Y(n_762) );
OAI211xp5_ASAP7_75t_SL g763 ( .A1(n_614), .A2(n_562), .B(n_525), .C(n_528), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g764 ( .A1(n_643), .A2(n_580), .B(n_528), .C(n_587), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_663), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_648), .B(n_527), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_661), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_657), .B(n_574), .Y(n_768) );
INVx2_ASAP7_75t_SL g769 ( .A(n_611), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_657), .B(n_574), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_665), .A2(n_539), .B1(n_541), .B2(n_546), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_671), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_650), .B(n_527), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_688), .B(n_585), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_654), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_617), .B(n_562), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_688), .B(n_584), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_692), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_659), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_708), .B(n_527), .Y(n_780) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_668), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_673), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_675), .Y(n_783) );
OR2x6_ASAP7_75t_L g784 ( .A(n_681), .B(n_562), .Y(n_784) );
AOI322xp5_ASAP7_75t_L g785 ( .A1(n_638), .A2(n_550), .A3(n_569), .B1(n_570), .B2(n_580), .C1(n_587), .C2(n_626), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_677), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_636), .B(n_569), .Y(n_787) );
OAI32xp33_ASAP7_75t_L g788 ( .A1(n_756), .A2(n_679), .A3(n_626), .B1(n_615), .B2(n_638), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_781), .B(n_697), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_723), .B(n_613), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_729), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_729), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_781), .B(n_668), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_775), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_735), .A2(n_637), .B1(n_639), .B2(n_651), .C(n_680), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_719), .B(n_720), .Y(n_796) );
NOR2xp33_ASAP7_75t_SL g797 ( .A(n_733), .B(n_666), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_779), .Y(n_798) );
AOI21xp33_ASAP7_75t_SL g799 ( .A1(n_733), .A2(n_679), .B(n_682), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_782), .Y(n_800) );
NOR2x1_ASAP7_75t_L g801 ( .A(n_756), .B(n_644), .Y(n_801) );
OAI32xp33_ASAP7_75t_L g802 ( .A1(n_726), .A2(n_623), .A3(n_683), .B1(n_672), .B2(n_662), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_783), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_735), .B(n_637), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_764), .A2(n_686), .B(n_642), .Y(n_805) );
NAND2x1p5_ASAP7_75t_L g806 ( .A(n_731), .B(n_641), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_740), .A2(n_664), .B1(n_670), .B2(n_550), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_741), .B(n_696), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_732), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_734), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_717), .B(n_694), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_740), .A2(n_716), .B(n_784), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_748), .B(n_698), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_730), .B(n_655), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_742), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_727), .B(n_653), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_743), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_723), .B(n_642), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_728), .B(n_701), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_744), .Y(n_820) );
AOI322xp5_ASAP7_75t_L g821 ( .A1(n_728), .A2(n_674), .A3(n_682), .B1(n_685), .B2(n_570), .C1(n_641), .C2(n_644), .Y(n_821) );
A2O1A1Ixp33_ASAP7_75t_L g822 ( .A1(n_785), .A2(n_686), .B(n_685), .C(n_699), .Y(n_822) );
XNOR2x1_ASAP7_75t_L g823 ( .A(n_767), .B(n_700), .Y(n_823) );
AO22x1_ASAP7_75t_L g824 ( .A1(n_731), .A2(n_710), .B1(n_676), .B2(n_678), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_747), .Y(n_825) );
INVxp67_ASAP7_75t_L g826 ( .A(n_718), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_765), .B(n_690), .Y(n_827) );
AOI21xp33_ASAP7_75t_R g828 ( .A1(n_746), .A2(n_622), .B(n_687), .Y(n_828) );
O2A1O1Ixp33_ASAP7_75t_L g829 ( .A1(n_822), .A2(n_753), .B(n_763), .C(n_750), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_795), .B(n_758), .Y(n_830) );
OR2x2_ASAP7_75t_L g831 ( .A(n_793), .B(n_770), .Y(n_831) );
INVxp33_ASAP7_75t_L g832 ( .A(n_801), .Y(n_832) );
NOR3x1_ASAP7_75t_L g833 ( .A(n_824), .B(n_769), .C(n_745), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_822), .A2(n_761), .B1(n_754), .B2(n_749), .C(n_762), .Y(n_834) );
OAI22xp5_ASAP7_75t_SL g835 ( .A1(n_806), .A2(n_784), .B1(n_780), .B2(n_765), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_807), .B(n_745), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_826), .Y(n_837) );
INVx1_ASAP7_75t_SL g838 ( .A(n_823), .Y(n_838) );
OAI211xp5_ASAP7_75t_SL g839 ( .A1(n_821), .A2(n_771), .B(n_750), .C(n_758), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_794), .B(n_768), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_788), .A2(n_770), .B1(n_768), .B2(n_722), .C(n_738), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_812), .A2(n_784), .B(n_780), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_797), .A2(n_751), .B(n_763), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_826), .Y(n_844) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_807), .A2(n_755), .B1(n_776), .B2(n_766), .C(n_773), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_802), .A2(n_736), .B1(n_778), .B2(n_772), .C(n_752), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g847 ( .A1(n_828), .A2(n_759), .B1(n_760), .B2(n_776), .C(n_787), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_798), .Y(n_848) );
INVx2_ASAP7_75t_SL g849 ( .A(n_823), .Y(n_849) );
O2A1O1Ixp5_ASAP7_75t_L g850 ( .A1(n_805), .A2(n_751), .B(n_786), .C(n_725), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_799), .B(n_724), .Y(n_851) );
AOI31xp33_ASAP7_75t_L g852 ( .A1(n_806), .A2(n_721), .A3(n_737), .B(n_739), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_804), .A2(n_777), .B1(n_774), .B2(n_757), .Y(n_853) );
AOI211xp5_ASAP7_75t_SL g854 ( .A1(n_813), .A2(n_622), .B(n_691), .C(n_703), .Y(n_854) );
NOR3xp33_ASAP7_75t_L g855 ( .A(n_791), .B(n_706), .C(n_707), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_789), .A2(n_689), .B1(n_796), .B2(n_819), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_796), .A2(n_790), .B(n_818), .C(n_792), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_800), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_803), .A2(n_815), .B1(n_809), .B2(n_810), .C(n_825), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_817), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g861 ( .A1(n_820), .A2(n_827), .B(n_808), .C(n_816), .Y(n_861) );
AOI221x1_ASAP7_75t_L g862 ( .A1(n_839), .A2(n_842), .B1(n_843), .B2(n_830), .C(n_835), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_851), .A2(n_838), .B(n_850), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_849), .B(n_851), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_833), .B(n_832), .Y(n_865) );
OAI211xp5_ASAP7_75t_SL g866 ( .A1(n_834), .A2(n_841), .B(n_829), .C(n_846), .Y(n_866) );
OAI211xp5_ASAP7_75t_L g867 ( .A1(n_847), .A2(n_861), .B(n_845), .C(n_836), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_866), .B(n_859), .C(n_852), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_864), .B(n_844), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_865), .B(n_837), .Y(n_870) );
NAND3xp33_ASAP7_75t_SL g871 ( .A(n_863), .B(n_854), .C(n_857), .Y(n_871) );
NOR3xp33_ASAP7_75t_L g872 ( .A(n_871), .B(n_867), .C(n_862), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_870), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_868), .A2(n_856), .B1(n_860), .B2(n_858), .C(n_848), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_873), .Y(n_875) );
AOI211x1_ASAP7_75t_L g876 ( .A1(n_874), .A2(n_869), .B(n_853), .C(n_840), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_876), .B(n_872), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_875), .A2(n_840), .B1(n_831), .B2(n_855), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_877), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_879), .B(n_878), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_880), .B(n_827), .Y(n_881) );
OR2x6_ASAP7_75t_L g882 ( .A(n_881), .B(n_808), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_811), .B1(n_814), .B2(n_872), .Y(n_883) );
endmodule