module fake_jpeg_6230_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_15),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_24),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_16),
.B1(n_21),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_24),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_58),
.B1(n_39),
.B2(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_58),
.C(n_50),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_44),
.B1(n_40),
.B2(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_88),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_57),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_63),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_47),
.B(n_60),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_66),
.B(n_61),
.Y(n_106)
);

NAND2x1_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_47),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_77),
.B(n_66),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_74),
.B(n_78),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_106),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_112),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_69),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_108),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_70),
.B1(n_64),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_107),
.B1(n_45),
.B2(n_51),
.Y(n_121)
);

XOR2x2_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_55),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_62),
.B1(n_52),
.B2(n_53),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_121),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_96),
.B1(n_92),
.B2(n_94),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_130),
.B1(n_100),
.B2(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_93),
.B1(n_88),
.B2(n_86),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_119),
.B(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_93),
.C(n_84),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_127),
.C(n_129),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_93),
.B(n_53),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_128),
.B(n_131),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_80),
.B1(n_45),
.B2(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_110),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_24),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_51),
.B1(n_42),
.B2(n_45),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_42),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_148),
.B1(n_19),
.B2(n_17),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_100),
.B1(n_80),
.B2(n_42),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_138),
.B1(n_141),
.B2(n_23),
.Y(n_159)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_146),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_104),
.B1(n_113),
.B2(n_83),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_87),
.C(n_19),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_87),
.Y(n_152)
);

NOR4xp25_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_132),
.C(n_117),
.D(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_83),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_105),
.C(n_29),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_105),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_134),
.B(n_9),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_29),
.C(n_23),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_141),
.C(n_148),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_140),
.B(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_23),
.C(n_17),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_147),
.C(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_137),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_22),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_22),
.C(n_12),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_20),
.B1(n_10),
.B2(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_183),
.C(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_181),
.Y(n_184)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_8),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_173),
.A2(n_160),
.B1(n_153),
.B2(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_155),
.C(n_1),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_0),
.C(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_175),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_199),
.B(n_205),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_194),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_182),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_0),
.Y(n_212)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_1),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_176),
.CI(n_8),
.CON(n_203),
.SN(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_193),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_176),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_210),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_186),
.A3(n_190),
.B1(n_8),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_202),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_213),
.B(n_3),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_200),
.C(n_2),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_218),
.C(n_5),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_201),
.C(n_203),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_5),
.B(n_6),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_2),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_5),
.B(n_6),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_212),
.C(n_4),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_3),
.B(n_4),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_223),
.B(n_224),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_219),
.B(n_6),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_7),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.C(n_222),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_7),
.Y(n_230)
);


endmodule