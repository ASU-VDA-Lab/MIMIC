module fake_jpeg_15986_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_1),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_56),
.B(n_63),
.C(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_88),
.B1(n_49),
.B2(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_50),
.B1(n_47),
.B2(n_62),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_91),
.B(n_55),
.C(n_52),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_50),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_85),
.C(n_2),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_98),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_109),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_59),
.B1(n_58),
.B2(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_1),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_49),
.B1(n_65),
.B2(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_85),
.B(n_88),
.C(n_3),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_96),
.C(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_117),
.C(n_125),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_126),
.B1(n_122),
.B2(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_25),
.C(n_44),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_110),
.B(n_97),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_131),
.B(n_133),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_113),
.B1(n_107),
.B2(n_92),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_26),
.B1(n_43),
.B2(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_22),
.B1(n_37),
.B2(n_36),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_132),
.C(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_118),
.B1(n_123),
.B2(n_120),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_142),
.B1(n_5),
.B2(n_6),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_131),
.B1(n_128),
.B2(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_24),
.B(n_27),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_18),
.B(n_35),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_115),
.B1(n_119),
.B2(n_7),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_134),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_143),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_145),
.B1(n_150),
.B2(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_46),
.Y(n_154)
);

AOI211xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_34),
.B(n_32),
.C(n_31),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_29),
.B(n_28),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_30),
.B(n_8),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_7),
.B(n_8),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_9),
.B(n_10),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_162)
);


endmodule