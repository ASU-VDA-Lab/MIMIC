module fake_jpeg_11604_n_514 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_63),
.Y(n_115)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_29),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_67),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_66),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_1),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_1),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_89),
.Y(n_144)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_95),
.Y(n_156)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_125),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_35),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_148),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_135),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_55),
.Y(n_140)
);

INVx5_ASAP7_75t_SL g193 ( 
.A(n_140),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_69),
.Y(n_148)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_154),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_177),
.Y(n_230)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_162),
.Y(n_250)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_165),
.B(n_170),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_87),
.B1(n_82),
.B2(n_81),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_202),
.B1(n_210),
.B2(n_150),
.Y(n_225)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_61),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_168),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_100),
.B1(n_59),
.B2(n_61),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_169),
.A2(n_185),
.B1(n_204),
.B2(n_20),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_108),
.B(n_54),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_65),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_173),
.B(n_174),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_127),
.B(n_78),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_76),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_91),
.B1(n_70),
.B2(n_34),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_178),
.B(n_92),
.Y(n_252)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_179),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_115),
.B(n_101),
.C(n_94),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_27),
.C(n_42),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_66),
.B(n_69),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_146),
.B(n_123),
.Y(n_231)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_96),
.B1(n_90),
.B2(n_88),
.Y(n_185)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_37),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_26),
.Y(n_194)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_48),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_212),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_103),
.A2(n_75),
.B1(n_74),
.B2(n_111),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_35),
.Y(n_203)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_120),
.A2(n_45),
.B1(n_48),
.B2(n_24),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_20),
.B1(n_56),
.B2(n_68),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_31),
.B1(n_32),
.B2(n_139),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_119),
.A2(n_69),
.B1(n_55),
.B2(n_19),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_207),
.B1(n_24),
.B2(n_38),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_137),
.A2(n_19),
.B1(n_31),
.B2(n_32),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_104),
.A2(n_24),
.B1(n_38),
.B2(n_32),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_36),
.A3(n_27),
.B1(n_42),
.B2(n_20),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_118),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_150),
.B1(n_149),
.B2(n_114),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_237),
.B1(n_244),
.B2(n_246),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_217),
.A2(n_207),
.B1(n_206),
.B2(n_161),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_240),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_195),
.B(n_171),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_245),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_252),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_149),
.B1(n_143),
.B2(n_136),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_121),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_143),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_247),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_136),
.B1(n_134),
.B2(n_130),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_134),
.B1(n_130),
.B2(n_114),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_168),
.B(n_164),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_118),
.B1(n_139),
.B2(n_172),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_175),
.B(n_2),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_31),
.B1(n_38),
.B2(n_27),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_261),
.B1(n_192),
.B2(n_195),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_178),
.A2(n_36),
.B1(n_42),
.B2(n_27),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

O2A1O1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_193),
.B(n_206),
.C(n_166),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_277),
.B1(n_286),
.B2(n_291),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_224),
.B(n_196),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_272),
.B(n_281),
.Y(n_336)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_191),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_289),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_292),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_201),
.B1(n_162),
.B2(n_187),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_192),
.C(n_191),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_222),
.C(n_243),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_251),
.B(n_199),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_240),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_247),
.B(n_186),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_294),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_287),
.A2(n_243),
.B(n_239),
.Y(n_328)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_232),
.B(n_176),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_290),
.B(n_295),
.Y(n_337)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

BUFx4f_ASAP7_75t_SL g293 ( 
.A(n_242),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_293),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_240),
.B(n_179),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_297),
.B(n_298),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_304),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_219),
.A2(n_201),
.B1(n_189),
.B2(n_187),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_234),
.B1(n_258),
.B2(n_189),
.Y(n_333)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_276),
.A2(n_225),
.B1(n_241),
.B2(n_237),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_226),
.CI(n_236),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_293),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_331),
.C(n_280),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_217),
.B1(n_231),
.B2(n_230),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_217),
.B1(n_248),
.B2(n_260),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_274),
.A2(n_249),
.B1(n_257),
.B2(n_256),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_283),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_302),
.Y(n_322)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_282),
.Y(n_323)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

AOI32xp33_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_296),
.A3(n_284),
.B1(n_294),
.B2(n_275),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_326),
.B(n_270),
.Y(n_357)
);

CKINVDCx10_ASAP7_75t_R g347 ( 
.A(n_328),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_250),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_334),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_229),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_333),
.A2(n_339),
.B1(n_299),
.B2(n_271),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_258),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_286),
.A2(n_234),
.B1(n_42),
.B2(n_36),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_279),
.B(n_216),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_266),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_287),
.A2(n_279),
.B(n_298),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_343),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_267),
.B1(n_265),
.B2(n_263),
.Y(n_344)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_262),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_348),
.B(n_360),
.Y(n_382)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_357),
.C(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_317),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_364),
.C(n_366),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_293),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_369),
.Y(n_391)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_304),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_330),
.B(n_292),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_324),
.B(n_278),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_363),
.B(n_367),
.Y(n_397)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_289),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_300),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_310),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_273),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_332),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_373),
.Y(n_400)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_310),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_374),
.A2(n_350),
.B1(n_351),
.B2(n_365),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_311),
.B(n_211),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_2),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_340),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_367),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_388),
.B1(n_398),
.B2(n_380),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_346),
.A2(n_335),
.B1(n_319),
.B2(n_309),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_384),
.A2(n_407),
.B1(n_371),
.B2(n_360),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_329),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_329),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_356),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_343),
.B(n_335),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_390),
.A2(n_362),
.B(n_340),
.Y(n_421)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_311),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_396),
.B(n_338),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_403),
.B1(n_406),
.B2(n_380),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g401 ( 
.A(n_345),
.B(n_321),
.CI(n_353),
.CON(n_401),
.SN(n_401)
);

FAx1_ASAP7_75t_SL g414 ( 
.A(n_401),
.B(n_364),
.CI(n_375),
.CON(n_414),
.SN(n_414)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_350),
.A2(n_342),
.B1(n_314),
.B2(n_307),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_368),
.A2(n_318),
.B1(n_328),
.B2(n_305),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_369),
.A2(n_339),
.B1(n_314),
.B2(n_313),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_374),
.B1(n_373),
.B2(n_355),
.Y(n_408)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_428),
.B1(n_431),
.B2(n_383),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_354),
.B1(n_347),
.B2(n_376),
.Y(n_411)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_378),
.A2(n_354),
.B1(n_361),
.B2(n_352),
.Y(n_412)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_366),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_427),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_414),
.B(n_425),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_378),
.A2(n_313),
.B1(n_305),
.B2(n_372),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_415),
.A2(n_418),
.B1(n_422),
.B2(n_426),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_416),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_362),
.B1(n_338),
.B2(n_327),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_422),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_393),
.B(n_392),
.Y(n_438)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_423),
.B(n_432),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_327),
.C(n_176),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_392),
.C(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_426),
.B(n_405),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_332),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_406),
.A2(n_180),
.B(n_80),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_180),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_430),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_38),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_404),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_4),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_421),
.A2(n_403),
.B(n_388),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_418),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_435),
.A2(n_437),
.B1(n_444),
.B2(n_415),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_410),
.A2(n_399),
.B1(n_398),
.B2(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_407),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_428),
.A2(n_381),
.B1(n_379),
.B2(n_395),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_449),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_401),
.C(n_397),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_413),
.C(n_427),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_453),
.B(n_454),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_425),
.C(n_430),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_457),
.B1(n_439),
.B2(n_461),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_419),
.Y(n_456)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_456),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_465),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_409),
.A3(n_419),
.B1(n_389),
.B2(n_395),
.C(n_428),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_458),
.B(n_462),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_SL g459 ( 
.A(n_448),
.B(n_414),
.C(n_401),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_459),
.B(n_451),
.Y(n_473)
);

INVx13_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_429),
.C(n_414),
.Y(n_462)
);

INVx13_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_463),
.A2(n_446),
.B(n_438),
.Y(n_472)
);

A2O1A1O1Ixp25_ASAP7_75t_L g466 ( 
.A1(n_448),
.A2(n_389),
.B(n_431),
.C(n_385),
.D(n_402),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_466),
.A2(n_434),
.B(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_402),
.C(n_5),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_452),
.C(n_5),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_467),
.A2(n_440),
.B1(n_443),
.B2(n_450),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_472),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_482),
.Y(n_483)
);

AOI21xp33_ASAP7_75t_L g492 ( 
.A1(n_473),
.A2(n_479),
.B(n_459),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_462),
.A2(n_443),
.B(n_435),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_475),
.B(n_478),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_476),
.A2(n_464),
.B1(n_455),
.B2(n_463),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_441),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_441),
.Y(n_479)
);

AO21x1_ASAP7_75t_L g484 ( 
.A1(n_479),
.A2(n_461),
.B(n_456),
.Y(n_484)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_453),
.C(n_454),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_486),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_478),
.C(n_471),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_492),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_477),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_488),
.B(n_491),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_468),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_482),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_480),
.B(n_436),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_469),
.C(n_481),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_4),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_460),
.Y(n_496)
);

AOI322xp5_ASAP7_75t_L g502 ( 
.A1(n_496),
.A2(n_489),
.A3(n_484),
.B1(n_493),
.B2(n_483),
.C1(n_490),
.C2(n_452),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_485),
.Y(n_501)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_500),
.B(n_6),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_497),
.A2(n_495),
.A3(n_500),
.B1(n_494),
.B2(n_498),
.C1(n_8),
.C2(n_9),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_504),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_5),
.B(n_6),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_508),
.B(n_509),
.Y(n_510)
);

O2A1O1Ixp33_ASAP7_75t_SL g509 ( 
.A1(n_506),
.A2(n_14),
.B(n_7),
.C(n_8),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_507),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_6),
.C(n_9),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_10),
.B(n_11),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_12),
.B(n_13),
.Y(n_514)
);


endmodule