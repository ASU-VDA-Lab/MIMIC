module fake_jpeg_28783_n_513 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_513);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_64),
.Y(n_115)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_65),
.Y(n_124)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_78),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_28),
.B(n_0),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_10),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_90),
.Y(n_157)
);

BUFx2_ASAP7_75t_R g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_103),
.B(n_119),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_105),
.A2(n_87),
.B1(n_84),
.B2(n_72),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_46),
.B1(n_37),
.B2(n_34),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_106),
.A2(n_20),
.B1(n_19),
.B2(n_21),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_18),
.B1(n_42),
.B2(n_46),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_107),
.A2(n_142),
.B1(n_99),
.B2(n_42),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_131),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_27),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_0),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_159),
.C(n_20),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_136),
.B(n_153),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_42),
.B1(n_18),
.B2(n_49),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_22),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_51),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_12),
.B(n_10),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_34),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_188),
.Y(n_229)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_167),
.Y(n_241)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_179),
.Y(n_227)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_101),
.B(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_180),
.B(n_197),
.Y(n_238)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_185),
.A2(n_192),
.B1(n_210),
.B2(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_186),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_42),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_196),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_126),
.A2(n_42),
.B1(n_76),
.B2(n_73),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_211),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_115),
.B(n_21),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_213),
.C(n_218),
.Y(n_246)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_199),
.Y(n_237)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_200),
.Y(n_253)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_204),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_31),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_209),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_208),
.A2(n_142),
.B1(n_127),
.B2(n_150),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_31),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_132),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_109),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_31),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_140),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_120),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_49),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_41),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_123),
.B1(n_160),
.B2(n_158),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_222),
.A2(n_224),
.B1(n_259),
.B2(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_171),
.A2(n_111),
.B1(n_160),
.B2(n_137),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_107),
.C(n_111),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_165),
.C(n_200),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_240),
.B(n_238),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_206),
.B(n_170),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_178),
.B(n_41),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_255),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_189),
.B(n_9),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_0),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_121),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_199),
.B(n_39),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_258),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_191),
.B(n_39),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_185),
.A2(n_127),
.B1(n_137),
.B2(n_139),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_128),
.B1(n_112),
.B2(n_163),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_156),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_268),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_192),
.A2(n_156),
.B1(n_150),
.B2(n_71),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_175),
.B(n_19),
.Y(n_268)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

BUFx4f_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_274),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_43),
.B(n_194),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_273),
.A2(n_307),
.B(n_258),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_277),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_288),
.Y(n_327)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_181),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_281),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_283),
.B1(n_264),
.B2(n_221),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_229),
.A2(n_162),
.B1(n_215),
.B2(n_214),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_226),
.Y(n_341)
);

AOI32xp33_ASAP7_75t_L g287 ( 
.A1(n_223),
.A2(n_206),
.A3(n_184),
.B1(n_165),
.B2(n_205),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_287),
.A2(n_306),
.B(n_257),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_219),
.B1(n_169),
.B2(n_183),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_31),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_295),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_242),
.A2(n_219),
.B1(n_120),
.B2(n_169),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_310),
.B1(n_311),
.B2(n_221),
.Y(n_326)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_31),
.C(n_43),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_300),
.C(n_231),
.Y(n_320)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_43),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_266),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_43),
.Y(n_298)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_43),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_301),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_233),
.B(n_1),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_242),
.B(n_1),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_1),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_244),
.B(n_2),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_304),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_248),
.B(n_229),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_230),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_305),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_232),
.B(n_2),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_261),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_3),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_241),
.B(n_265),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_250),
.B1(n_228),
.B2(n_241),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_317),
.A2(n_344),
.B1(n_245),
.B2(n_249),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_341),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_326),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_285),
.B(n_268),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_324),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_345),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_328),
.B(n_348),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_246),
.A3(n_223),
.B1(n_234),
.B2(n_237),
.Y(n_331)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_232),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_340),
.C(n_343),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_276),
.A2(n_239),
.B1(n_224),
.B2(n_267),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_335),
.A2(n_346),
.B1(n_299),
.B2(n_293),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_273),
.A2(n_226),
.B(n_243),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_235),
.C(n_251),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_235),
.C(n_251),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_276),
.A2(n_288),
.B1(n_275),
.B2(n_287),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_225),
.C(n_247),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_284),
.A2(n_288),
.B1(n_297),
.B2(n_307),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_272),
.B(n_293),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_301),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_253),
.B(n_264),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

OR2x4_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_311),
.Y(n_353)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_288),
.B1(n_272),
.B2(n_292),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_355),
.A2(n_317),
.B1(n_345),
.B2(n_329),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_371),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

AOI21xp33_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_334),
.B(n_331),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_343),
.C(n_340),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_347),
.B(n_303),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_364),
.Y(n_383)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_332),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_336),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

AO22x1_ASAP7_75t_SL g371 ( 
.A1(n_327),
.A2(n_346),
.B1(n_335),
.B2(n_324),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_327),
.A2(n_270),
.B1(n_274),
.B2(n_253),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_376),
.Y(n_390)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_323),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_378),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_315),
.B(n_338),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_281),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_380),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_312),
.B(n_225),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_381),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_278),
.Y(n_382)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_386),
.B(n_402),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_388),
.C(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_368),
.C(n_356),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_341),
.C(n_320),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_382),
.B(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_394),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_354),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_399),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_342),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_354),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_411),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_405),
.A2(n_408),
.B1(n_374),
.B2(n_333),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_279),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_407),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_355),
.A2(n_325),
.B1(n_339),
.B2(n_321),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_351),
.A2(n_350),
.B(n_353),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_410),
.A2(n_392),
.B(n_408),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_393),
.B(n_356),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_391),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_362),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_384),
.A2(n_350),
.B1(n_351),
.B2(n_367),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_416),
.A2(n_423),
.B1(n_395),
.B2(n_406),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_409),
.Y(n_419)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_422),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_384),
.A2(n_367),
.B1(n_371),
.B2(n_357),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_424),
.A2(n_433),
.B1(n_406),
.B2(n_404),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_405),
.A2(n_392),
.B1(n_396),
.B2(n_400),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_425),
.A2(n_310),
.B1(n_260),
.B2(n_247),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_426),
.B(n_430),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_401),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_368),
.C(n_373),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_435),
.C(n_403),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_394),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_410),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_436),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_389),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_432),
.B(n_434),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_411),
.A2(n_398),
.B1(n_390),
.B2(n_404),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_349),
.B(n_380),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_365),
.C(n_318),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_318),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_439),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_443),
.C(n_448),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_321),
.C(n_403),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_422),
.A2(n_391),
.B1(n_385),
.B2(n_409),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_452),
.C(n_435),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_385),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_291),
.C(n_278),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_420),
.C(n_424),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g450 ( 
.A(n_413),
.B(n_295),
.CI(n_269),
.CON(n_450),
.SN(n_450)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_375),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_455),
.A2(n_419),
.B1(n_423),
.B2(n_434),
.Y(n_458)
);

INVx13_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_458),
.A2(n_465),
.B1(n_445),
.B2(n_438),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_440),
.B(n_426),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_461),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_444),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_5),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_421),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_469),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_453),
.A2(n_418),
.B1(n_416),
.B2(n_412),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_452),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_425),
.C(n_433),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_437),
.B(n_413),
.CI(n_428),
.CON(n_470),
.SN(n_470)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_447),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_471),
.B(n_364),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_436),
.C(n_245),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_472),
.A2(n_442),
.B(n_449),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_473),
.B(n_484),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_476),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_465),
.A2(n_456),
.B1(n_451),
.B2(n_454),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_477),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_448),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_464),
.A2(n_455),
.B1(n_446),
.B2(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_479),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_458),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_3),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_472),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_489),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_464),
.B1(n_459),
.B2(n_457),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_485),
.B(n_466),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_494),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_483),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_495),
.B(n_470),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_491),
.C(n_488),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_477),
.C(n_466),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_498),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_490),
.A2(n_470),
.B(n_459),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_492),
.A2(n_482),
.B1(n_484),
.B2(n_469),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_499),
.A2(n_479),
.B1(n_488),
.B2(n_462),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_504),
.Y(n_507)
);

AOI322xp5_ASAP7_75t_L g505 ( 
.A1(n_500),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_491),
.C1(n_480),
.C2(n_457),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_6),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_506),
.B(n_501),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_508),
.A2(n_507),
.B(n_505),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_503),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_7),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_7),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_7),
.Y(n_513)
);


endmodule