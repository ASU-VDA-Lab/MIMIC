module real_jpeg_24275_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_358, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_358;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_8),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_4),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_182),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_4),
.A2(n_111),
.B1(n_112),
.B2(n_182),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_4),
.A2(n_174),
.B1(n_182),
.B2(n_199),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_42),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_68),
.B1(n_92),
.B2(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_111),
.B(n_115),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_SL g151 ( 
.A(n_6),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_7),
.A2(n_51),
.B1(n_111),
.B2(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_7),
.A2(n_51),
.B1(n_174),
.B2(n_199),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_65),
.B1(n_111),
.B2(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_10),
.A2(n_65),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_73),
.B1(n_111),
.B2(n_112),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_11),
.A2(n_73),
.B1(n_199),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_132),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_111),
.B1(n_112),
.B2(n_132),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_12),
.A2(n_132),
.B1(n_199),
.B2(n_218),
.Y(n_288)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_13),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_155),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_15),
.A2(n_111),
.B1(n_112),
.B2(n_155),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_15),
.A2(n_155),
.B1(n_173),
.B2(n_200),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_16),
.A2(n_76),
.B1(n_111),
.B2(n_112),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_16),
.A2(n_76),
.B1(n_177),
.B2(n_266),
.Y(n_265)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_17),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_355),
.C(n_356),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_351),
.B(n_354),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_337),
.B(n_350),
.Y(n_22)
);

OAI321xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_302),
.A3(n_330),
.B1(n_335),
.B2(n_336),
.C(n_358),
.Y(n_23)
);

AOI311xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_249),
.A3(n_293),
.B(n_296),
.C(n_297),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_204),
.C(n_244),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_167),
.B(n_203),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_136),
.B(n_166),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_105),
.B(n_135),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_79),
.B(n_104),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_54),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_31),
.B(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_52),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_32),
.A2(n_33),
.B1(n_52),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_35),
.B(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_38),
.B(n_44),
.C(n_53),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_36),
.A2(n_60),
.A3(n_111),
.B1(n_116),
.B2(n_127),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_38),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_38),
.B(n_177),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_38),
.A2(n_174),
.B(n_176),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_39),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_39),
.A2(n_45),
.B1(n_224),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_39),
.A2(n_242),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_40),
.A2(n_63),
.B1(n_64),
.B2(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_40),
.A2(n_163),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_40),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_40),
.A2(n_63),
.B(n_163),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_45),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_45),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_66),
.C(n_67),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_118),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_58),
.A2(n_118),
.B1(n_143),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_58),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_58),
.A2(n_118),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_58),
.A2(n_118),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_110),
.B1(n_117),
.B2(n_120),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_59),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_59),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_61),
.B1(n_111),
.B2(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_63),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_78),
.B1(n_83),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_68),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_68),
.A2(n_130),
.B(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_68),
.A2(n_129),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_69),
.B(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_69),
.A2(n_77),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_74),
.B(n_156),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B(n_103),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_86),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_102),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_125),
.B1(n_133),
.B2(n_134),
.Y(n_107)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_112),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_149),
.A3(n_173),
.B1(n_176),
.B2(n_178),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_117),
.A2(n_213),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_118),
.A2(n_191),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_118),
.B(n_237),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_118),
.A2(n_277),
.B(n_313),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_124),
.C(n_133),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_157),
.B2(n_158),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_160),
.C(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_146),
.C(n_152),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_153),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_147),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_147),
.A2(n_196),
.B1(n_202),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_147),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_147),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_147),
.A2(n_196),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_147),
.A2(n_196),
.B(n_265),
.Y(n_355)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_148),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_148),
.A2(n_197),
.B1(n_216),
.B2(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_148),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_150),
.B1(n_174),
.B2(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_162),
.B(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_169),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_188),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_187),
.C(n_188),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_179),
.B1(n_183),
.B2(n_184),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_183),
.Y(n_209)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.C(n_195),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_196),
.B(n_288),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_196),
.A2(n_323),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_197),
.A2(n_233),
.B(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_197),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_205),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_227),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_206),
.B(n_227),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_219),
.C(n_220),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_208),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_212),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_213),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_219),
.B(n_220),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_223),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_227),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_239),
.CI(n_243),
.CON(n_227),
.SN(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_238),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_235),
.C(n_238),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_245),
.B(n_246),
.Y(n_299)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_250),
.A2(n_294),
.B(n_298),
.C(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_272),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_251),
.B(n_295),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_259),
.CI(n_271),
.CON(n_251),
.SN(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_256),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_258),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_258),
.A2(n_281),
.B(n_285),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_270),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_263),
.C(n_267),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_264),
.B(n_308),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_265),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_268),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_292),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_280),
.B1(n_290),
.B2(n_291),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_304),
.B1(n_316),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_290),
.C(n_292),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_289),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_318),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_303),
.B(n_318),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_316),
.C(n_317),
.Y(n_303)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_315),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_306),
.B1(n_320),
.B2(n_328),
.Y(n_319)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_328),
.C(n_329),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_311),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_321),
.C(n_325),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_329),
.Y(n_318)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_349),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_338),
.B(n_349),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_348),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_343),
.C(n_345),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_352),
.B(n_353),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_352),
.Y(n_356)
);


endmodule