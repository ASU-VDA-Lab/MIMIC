module fake_jpeg_28339_n_48 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_48);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx2_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_30),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_1),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.C(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_41),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_14),
.C(n_17),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_31),
.C(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_40),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_45),
.B(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);


endmodule