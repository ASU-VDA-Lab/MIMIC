module fake_jpeg_14745_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_41),
.B(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_0),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_57),
.Y(n_102)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_66),
.Y(n_110)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_73),
.B(n_84),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_18),
.B1(n_36),
.B2(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_101),
.B1(n_109),
.B2(n_107),
.Y(n_150)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_21),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_97),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_30),
.B1(n_36),
.B2(n_27),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_100),
.B1(n_122),
.B2(n_37),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_36),
.B1(n_39),
.B2(n_26),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_45),
.A2(n_25),
.B1(n_37),
.B2(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_112),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_40),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_51),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_118),
.Y(n_144)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_41),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_64),
.A2(n_32),
.B1(n_39),
.B2(n_20),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_128),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_15),
.B(n_33),
.C(n_31),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_130),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_133),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_145),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g136 ( 
.A(n_87),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_136),
.Y(n_195)
);

OR2x2_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_31),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_142),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_157),
.Y(n_204)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_23),
.C(n_22),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_165),
.C(n_89),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_92),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_154),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_128),
.B(n_149),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_8),
.B1(n_11),
.B2(n_3),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_155),
.B1(n_161),
.B2(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_8),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_0),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_82),
.A2(n_13),
.B1(n_8),
.B2(n_5),
.Y(n_155)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_102),
.B(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_167),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_98),
.A2(n_96),
.B1(n_75),
.B2(n_71),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_86),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_7),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_166),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_0),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_94),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_101),
.B(n_1),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_144),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_173),
.B(n_206),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_74),
.B1(n_85),
.B2(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_197),
.Y(n_220)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_99),
.B1(n_111),
.B2(n_117),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_99),
.B1(n_111),
.B2(n_117),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_1),
.B1(n_123),
.B2(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_123),
.A2(n_1),
.B1(n_168),
.B2(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_202),
.B(n_136),
.Y(n_210)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_138),
.B(n_143),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_137),
.B(n_148),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_124),
.C(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_132),
.B(n_146),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_159),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_126),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_210),
.Y(n_244)
);

OR2x4_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_136),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_223),
.B(n_226),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_193),
.B(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_190),
.A2(n_159),
.B1(n_182),
.B2(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_172),
.B(n_205),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_172),
.A2(n_203),
.B(n_184),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.C(n_171),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_179),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_199),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_183),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_197),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_204),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_200),
.B(n_188),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_186),
.B(n_174),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_216),
.B(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_241),
.Y(n_279)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_176),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_209),
.B1(n_213),
.B2(n_218),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_170),
.C(n_174),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_170),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_219),
.B1(n_235),
.B2(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_181),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_181),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_209),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_235),
.C(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_263),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_234),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_211),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_284),
.B1(n_258),
.B2(n_256),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_271),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_216),
.B1(n_239),
.B2(n_221),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_274),
.B1(n_280),
.B2(n_281),
.Y(n_291)
);

OR2x6_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_231),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_276),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_232),
.B(n_222),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_215),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_245),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_251),
.C(n_244),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_243),
.B1(n_262),
.B2(n_240),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_290),
.A2(n_272),
.B1(n_279),
.B2(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_242),
.C(n_246),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_248),
.C(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_248),
.C(n_252),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_263),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_270),
.B(n_254),
.CI(n_240),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_304),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_287),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_307),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_273),
.B1(n_286),
.B2(n_268),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_269),
.B(n_280),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_308),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_273),
.B(n_277),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_273),
.B1(n_276),
.B2(n_275),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_311),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_273),
.C(n_278),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_273),
.B(n_275),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_298),
.B(n_213),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_302),
.C(n_299),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_289),
.C(n_293),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_292),
.C(n_211),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_311),
.B1(n_309),
.B2(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_319),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_314),
.C(n_318),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_315),
.B1(n_321),
.B2(n_320),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_327),
.Y(n_330)
);


endmodule