module real_jpeg_5935_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_1),
.A2(n_129),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_1),
.A2(n_129),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_49),
.B1(n_154),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_49),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_2),
.A2(n_49),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_2),
.A2(n_257),
.B(n_260),
.C(n_263),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_2),
.B(n_184),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_2),
.B(n_55),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_297),
.C(n_300),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_2),
.B(n_119),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_2),
.B(n_294),
.C(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_2),
.B(n_28),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_24),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_3),
.A2(n_24),
.B1(n_34),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_3),
.A2(n_24),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_4),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_81),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_81),
.B1(n_128),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_81),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_9),
.Y(n_259)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_11),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_421),
.B(n_424),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_417),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_139),
.B(n_416),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_18),
.B(n_132),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.C(n_130),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_19),
.B(n_413),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_84),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_20),
.A2(n_186),
.B1(n_187),
.B2(n_197),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_20),
.B(n_146),
.C(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_20),
.B(n_238),
.C(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_20),
.A2(n_197),
.B1(n_238),
.B2(n_341),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_20),
.A2(n_197),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_226)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_23),
.Y(n_127)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_46),
.B1(n_51),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_51),
.B1(n_126),
.B2(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_27),
.A2(n_46),
.B(n_51),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_27),
.A2(n_51),
.B(n_133),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_30),
.Y(n_320)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g261 ( 
.A(n_33),
.Y(n_261)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_39),
.Y(n_263)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_49),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_52),
.A2(n_84),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_52),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_52),
.B(n_226),
.C(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_52),
.A2(n_391),
.B1(n_393),
.B2(n_400),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_78),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_53),
.B(n_156),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_54),
.A2(n_65),
.B1(n_149),
.B2(n_155),
.Y(n_148)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_55),
.A2(n_201),
.B(n_205),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_55),
.B(n_150),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_55),
.A2(n_66),
.B1(n_78),
.B2(n_201),
.Y(n_237)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_57),
.Y(n_299)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_58),
.Y(n_221)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_59),
.Y(n_169)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_66),
.B(n_156),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_70),
.Y(n_295)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_75),
.Y(n_203)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_84),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B1(n_119),
.B2(n_120),
.Y(n_84)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_85),
.Y(n_394)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_93),
.B(n_225),
.Y(n_395)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_109),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_94),
.A2(n_109),
.B1(n_188),
.B2(n_194),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_94),
.A2(n_109),
.B1(n_188),
.B2(n_194),
.Y(n_238)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_105),
.Y(n_325)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_109),
.A2(n_394),
.B(n_395),
.Y(n_393)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_125),
.B(n_130),
.Y(n_413)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_131),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_132),
.B(n_419),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_132),
.B(n_419),
.Y(n_420)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_411),
.B(n_415),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_382),
.B(n_408),
.Y(n_140)
);

OAI211xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_271),
.B(n_376),
.C(n_381),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_243),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_143),
.A2(n_243),
.B(n_377),
.C(n_380),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_227),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_144),
.B(n_227),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_198),
.C(n_212),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_145),
.B(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_185),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_158),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_147),
.A2(n_148),
.B1(n_158),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_147),
.A2(n_148),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_147),
.A2(n_148),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_148),
.B(n_265),
.C(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_148),
.B(n_333),
.C(n_335),
.Y(n_346)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_158),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_166),
.B1(n_174),
.B2(n_181),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_160),
.A2(n_182),
.B(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_163),
.Y(n_301)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_218),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_167),
.A2(n_218),
.B1(n_266),
.B2(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_173),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_178),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_186),
.A2(n_187),
.B1(n_222),
.B2(n_292),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_186),
.B(n_292),
.C(n_315),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_186),
.A2(n_187),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_187),
.B(n_226),
.C(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_207),
.B2(n_211),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_211),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_207),
.A2(n_233),
.B(n_234),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_208),
.B(n_218),
.Y(n_326)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_224),
.C(n_226),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_215),
.A2(n_222),
.B1(n_292),
.B2(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_222),
.A2(n_292),
.B1(n_293),
.B2(n_302),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_224),
.A2(n_226),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_226),
.A2(n_250),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_226),
.A2(n_250),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_226),
.A2(n_250),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_226),
.B(n_387),
.C(n_392),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_241),
.B2(n_242),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_235),
.B(n_240),
.C(n_242),
.Y(n_407)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_238),
.A2(n_337),
.B1(n_338),
.B2(n_341),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_238),
.Y(n_341)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_239),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_239),
.A2(n_397),
.B1(n_401),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_244),
.B(n_246),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.C(n_254),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_247),
.A2(n_248),
.B1(n_252),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_252),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_254),
.B(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_255),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_256),
.A2(n_264),
.B1(n_265),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_265),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_268),
.Y(n_280)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_360),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_345),
.B(n_359),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_330),
.B(n_344),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_312),
.B(n_329),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_304),
.B(n_311),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_289),
.B(n_303),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_286),
.B(n_288),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_290),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_339),
.C(n_341),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_314),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_328),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_326),
.B2(n_327),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_343),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_343),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_335),
.B1(n_336),
.B2(n_342),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_347),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_355),
.C(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_351),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_370),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_369),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_369),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_368),
.C(n_372),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_378),
.B(n_379),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_373),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_403),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_396),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_396),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_392),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.C(n_402),
.Y(n_396)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_397),
.Y(n_406)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_407),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_414),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

BUFx4f_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_422),
.Y(n_425)
);

INVx13_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);


endmodule