module fake_jpeg_15629_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_17),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_39),
.B1(n_33),
.B2(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_58),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_30),
.B1(n_27),
.B2(n_42),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_17),
.B1(n_24),
.B2(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_65),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_31),
.C(n_36),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_71),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_46),
.B1(n_49),
.B2(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_30),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_19),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_47),
.C(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_34),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_56),
.B1(n_65),
.B2(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_78),
.B1(n_86),
.B2(n_57),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_19),
.B1(n_33),
.B2(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_84),
.B1(n_94),
.B2(n_66),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

OAI22x1_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_47),
.B1(n_41),
.B2(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_78),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_49),
.B(n_3),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_57),
.B(n_29),
.C(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_88),
.B1(n_94),
.B2(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_25),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_63),
.B1(n_74),
.B2(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_90),
.B1(n_89),
.B2(n_83),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_72),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_92),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_99),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_20),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_87),
.C(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_116),
.B1(n_128),
.B2(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_125),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_64),
.C(n_45),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_128),
.C(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_64),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_100),
.A3(n_103),
.B1(n_104),
.B2(n_97),
.C(n_29),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_108),
.C(n_109),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_132),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_95),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_110),
.C(n_111),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_140),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_98),
.B1(n_123),
.B2(n_114),
.C(n_115),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

BUFx12f_ASAP7_75t_SL g135 ( 
.A(n_127),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_138),
.B1(n_54),
.B2(n_53),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_18),
.B(n_21),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_20),
.C(n_28),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_126),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_139),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_150),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_119),
.C(n_118),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_2),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_151),
.B(n_18),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_143),
.B1(n_26),
.B2(n_25),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_28),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_158),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_148),
.Y(n_161)
);

NOR2x1_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_139),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C(n_10),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_26),
.B(n_23),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_156),
.B(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_170),
.B1(n_161),
.B2(n_23),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

AOI31xp33_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_11),
.A3(n_12),
.B(n_13),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_167),
.C(n_21),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_172),
.A3(n_11),
.B1(n_7),
.B2(n_5),
.C(n_21),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_5),
.C(n_7),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_54),
.Y(n_179)
);


endmodule