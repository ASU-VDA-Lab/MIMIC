module fake_netlist_5_1000_n_4355 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_422, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_441, n_450, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_4355);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_422;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_441;
input n_450;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_4355;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_3241;
wire n_4129;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2955;
wire n_2899;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_880;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_956;
wire n_564;
wire n_4240;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_4109;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3039;
wire n_3019;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_1860;
wire n_2543;
wire n_4155;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_556;
wire n_3036;
wire n_2482;
wire n_3695;
wire n_3891;
wire n_4145;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1705;
wire n_659;
wire n_1294;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3937;
wire n_3696;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_4315;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2561;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_3298;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_696;
wire n_550;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_475;
wire n_1070;
wire n_777;
wire n_1547;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_521;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_1587;
wire n_1473;
wire n_680;
wire n_2682;
wire n_553;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1556;
wire n_1384;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2980;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_3191;
wire n_571;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3837;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_3915;
wire n_2370;
wire n_3496;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3735;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_4067;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_593;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_3781;
wire n_1385;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_4353;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4161;
wire n_647;
wire n_3433;
wire n_4024;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_3392;
wire n_3430;
wire n_3975;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_561;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_4151;
wire n_4148;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_4252;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4331;
wire n_4160;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_3989;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_558;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_702;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_3981;
wire n_2108;
wire n_3640;
wire n_728;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_809;
wire n_3923;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2825;
wire n_2813;
wire n_1888;
wire n_2009;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_2064;
wire n_784;
wire n_3978;
wire n_4325;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_776;
wire n_1798;
wire n_2022;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_3416;
wire n_525;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_744;
wire n_590;
wire n_629;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_498;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3113;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4078;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_568;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_3205;
wire n_4156;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_524;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4154;
wire n_535;
wire n_3396;
wire n_3701;
wire n_940;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_514;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_636;
wire n_3741;
wire n_660;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_2029;
wire n_750;
wire n_995;
wire n_3221;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_3990;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_473;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_974;
wire n_2565;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_3149;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_3466;
wire n_3458;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_3960;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2477;
wire n_761;
wire n_2277;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3905;
wire n_4329;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2879;
wire n_2474;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_512;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3077;
wire n_3929;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2424;
wire n_2255;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_860;
wire n_3229;
wire n_4213;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4084;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_513;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3618;
wire n_3592;
wire n_4031;
wire n_495;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4339;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4060;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_1630;
wire n_2122;
wire n_716;
wire n_2512;
wire n_3589;
wire n_4102;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_3993;
wire n_2216;
wire n_531;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_890;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_950;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_3847;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3548;
wire n_912;
wire n_968;
wire n_3569;
wire n_4348;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_3953;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_483;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_762;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3231;
wire n_3105;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4286;
wire n_3864;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3866;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_3255;
wire n_2675;
wire n_2743;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4047;
wire n_543;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_470;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_918;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_540;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2393;
wire n_2318;
wire n_3689;
wire n_2020;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2471;
wire n_2298;
wire n_1807;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3861;
wire n_3780;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_4117;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_661;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_510;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1603;
wire n_1232;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4062;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_2492;
wire n_1998;
wire n_1105;
wire n_1019;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_4336;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_3324;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_2409;
wire n_917;
wire n_601;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_3839;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_3972;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_500;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_541;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_536;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_827;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_3968;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2430;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_703;
wire n_980;
wire n_1115;
wire n_698;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3239;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3172;
wire n_2598;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_737;
wire n_4050;
wire n_3700;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_760;
wire n_3858;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_481;
wire n_2772;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_4178;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_4092;
wire n_930;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_622;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_682;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_4015;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3265;
wire n_3050;
wire n_1857;
wire n_4056;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_479;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_839;
wire n_3551;
wire n_3903;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_598;
wire n_685;
wire n_608;
wire n_1367;
wire n_928;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_499;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_517;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_4287;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4270;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_722;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_471;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_502;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_585;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3921;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_3930;
wire n_730;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_795;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_695;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_657;
wire n_4320;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_491;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4245;
wire n_4288;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_1181;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_3225;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_3799;
wire n_4119;
wire n_1254;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4009;
wire n_3159;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_99),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_10),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_57),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_335),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_57),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_332),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_129),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_198),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_316),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_249),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_342),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_16),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_342),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_113),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_183),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_407),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_350),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_143),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_268),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_78),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_303),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_267),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_304),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_386),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_260),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_184),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_221),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_166),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_351),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_295),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_374),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_206),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_197),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_213),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_107),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_10),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_22),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_168),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_379),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_167),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_312),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_425),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_89),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_206),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_295),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_98),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_469),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_437),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_48),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_343),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_3),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_163),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_133),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_307),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_432),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_345),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_37),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_375),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_344),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_66),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_90),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_440),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_133),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_154),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_284),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_24),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_239),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_219),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_100),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_450),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_308),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_358),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_104),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_214),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_384),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_243),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_333),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_421),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_148),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_352),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_353),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_122),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_50),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_424),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_94),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_216),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_213),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_276),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_199),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_349),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_257),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_76),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_217),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_291),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_385),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_323),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_304),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_368),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_173),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_346),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_464),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_17),
.Y(n_579)
);

CKINVDCx14_ASAP7_75t_R g580 ( 
.A(n_243),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_250),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_92),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_451),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_284),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_66),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_5),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_37),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_252),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_38),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_417),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_68),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_297),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_467),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_222),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_111),
.Y(n_595)
);

HB1xp67_ASAP7_75t_SL g596 ( 
.A(n_336),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_107),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_221),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_24),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_270),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_44),
.Y(n_601)
);

BUFx2_ASAP7_75t_SL g602 ( 
.A(n_289),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_371),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_291),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_76),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_290),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_298),
.Y(n_607)
);

BUFx2_ASAP7_75t_R g608 ( 
.A(n_103),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_234),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_106),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_55),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_197),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_323),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_277),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_98),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_240),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_59),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_234),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_86),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_367),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_128),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_341),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_217),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_227),
.Y(n_624)
);

BUFx8_ASAP7_75t_SL g625 ( 
.A(n_135),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_328),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_293),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_29),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_130),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_86),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_383),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_124),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_427),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_281),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_391),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_204),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_271),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_168),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_223),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_463),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_167),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_64),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_224),
.Y(n_643)
);

BUFx5_ASAP7_75t_L g644 ( 
.A(n_263),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_47),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_303),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_321),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_299),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_103),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_179),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_71),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_444),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_287),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_81),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_183),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_63),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_152),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_433),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_458),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_460),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_53),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_156),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_413),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_398),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_117),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_33),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_11),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_276),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_380),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_238),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_468),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_128),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_166),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_403),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_208),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_282),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_46),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_321),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_236),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_419),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_347),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_144),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_302),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_406),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_441),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_260),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_237),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_275),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_77),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_14),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_382),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_58),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_4),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_72),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_11),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_443),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_6),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_191),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_117),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_269),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_74),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_93),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_190),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_115),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_397),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_429),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_139),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_334),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_393),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_453),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_80),
.Y(n_711)
);

INVxp33_ASAP7_75t_SL g712 ( 
.A(n_180),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_68),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_395),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_126),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_233),
.Y(n_716)
);

BUFx5_ASAP7_75t_L g717 ( 
.A(n_194),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_320),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_307),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_246),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_355),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_205),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_311),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_290),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_235),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_465),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_240),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_363),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_466),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_312),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_141),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_74),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_241),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_296),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_118),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_47),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_269),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_362),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_114),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_258),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_343),
.Y(n_741)
);

XNOR2x1_ASAP7_75t_L g742 ( 
.A(n_311),
.B(n_239),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_381),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_32),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_420),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_262),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_116),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_22),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_378),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_200),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_169),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_360),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_387),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_271),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_428),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_169),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_81),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_408),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_185),
.Y(n_759)
);

CKINVDCx14_ASAP7_75t_R g760 ( 
.A(n_92),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_159),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_26),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_50),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_12),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_120),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_131),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_118),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_388),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_729),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_644),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_617),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_678),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_644),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_644),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_644),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_644),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_625),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_748),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_644),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_644),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_476),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_543),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_717),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_543),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_517),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_717),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_489),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_729),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_717),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_717),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_526),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_717),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_490),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_717),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_717),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_767),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_767),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_497),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_707),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_588),
.Y(n_804)
);

INVx4_ASAP7_75t_R g805 ( 
.A(n_596),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_472),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_588),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_767),
.Y(n_809)
);

INVxp33_ASAP7_75t_L g810 ( 
.A(n_742),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_505),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_767),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_767),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_767),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_767),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_767),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_528),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_475),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_528),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_588),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_742),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_528),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_528),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_528),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_588),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_528),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_535),
.Y(n_827)
);

CKINVDCx16_ASAP7_75t_R g828 ( 
.A(n_748),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_535),
.Y(n_829)
);

INVxp33_ASAP7_75t_SL g830 ( 
.A(n_478),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_602),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_535),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_535),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_514),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_532),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_535),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_703),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_470),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_522),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_470),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_473),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_535),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_556),
.Y(n_844)
);

INVxp33_ASAP7_75t_SL g845 ( 
.A(n_479),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_487),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_531),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_602),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_534),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_473),
.Y(n_850)
);

INVxp33_ASAP7_75t_SL g851 ( 
.A(n_481),
.Y(n_851)
);

INVxp33_ASAP7_75t_L g852 ( 
.A(n_474),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_556),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_556),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_556),
.Y(n_855)
);

INVxp33_ASAP7_75t_L g856 ( 
.A(n_474),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_556),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_556),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_570),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_570),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_570),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_703),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_703),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_570),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_570),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_580),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_760),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_570),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_595),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_538),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_763),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_595),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_595),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_595),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_763),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_547),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_595),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_488),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_567),
.B(n_0),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_488),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_504),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_763),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_471),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_504),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_595),
.Y(n_885)
);

BUFx2_ASAP7_75t_SL g886 ( 
.A(n_567),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_618),
.Y(n_887)
);

INVxp33_ASAP7_75t_SL g888 ( 
.A(n_482),
.Y(n_888)
);

INVxp33_ASAP7_75t_SL g889 ( 
.A(n_483),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_618),
.Y(n_890)
);

INVxp33_ASAP7_75t_L g891 ( 
.A(n_477),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_618),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_618),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_471),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_763),
.B(n_0),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_618),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_618),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_492),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_672),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_672),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_532),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_672),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_672),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_549),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_672),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_552),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_512),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_672),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_555),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_682),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_558),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_575),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_577),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_682),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_682),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_557),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_910),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_898),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_868),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_868),
.Y(n_921)
);

OA21x2_ASAP7_75t_L g922 ( 
.A1(n_817),
.A2(n_578),
.B(n_557),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_772),
.A2(n_652),
.B(n_502),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_910),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_817),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_779),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_819),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_784),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_784),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_784),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_771),
.Y(n_931)
);

OAI22x1_ASAP7_75t_L g932 ( 
.A1(n_769),
.A2(n_553),
.B1(n_628),
.B2(n_480),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_810),
.A2(n_518),
.B1(n_559),
.B2(n_503),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_819),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_784),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_784),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_822),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_786),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_783),
.B(n_512),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_822),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_790),
.A2(n_754),
.B1(n_627),
.B2(n_712),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_786),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_786),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_823),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_804),
.B(n_512),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_808),
.B(n_631),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_823),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_786),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_824),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_820),
.B(n_631),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_825),
.B(n_631),
.Y(n_951)
);

CKINVDCx16_ASAP7_75t_R g952 ( 
.A(n_828),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_824),
.Y(n_953)
);

AND2x4_ASAP7_75t_SL g954 ( 
.A(n_846),
.B(n_471),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_786),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_826),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_840),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_840),
.Y(n_958)
);

OA21x2_ASAP7_75t_L g959 ( 
.A1(n_826),
.A2(n_583),
.B(n_578),
.Y(n_959)
);

OAI22x1_ASAP7_75t_SL g960 ( 
.A1(n_778),
.A2(n_591),
.B1(n_598),
.B2(n_585),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_827),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_837),
.B(n_603),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_772),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_835),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_827),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_829),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_829),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_773),
.B(n_678),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_785),
.A2(n_652),
.B(n_502),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_862),
.B(n_603),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_832),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_807),
.B(n_523),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_832),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_833),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_818),
.B(n_561),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_863),
.B(n_583),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_773),
.B(n_907),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_835),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_785),
.Y(n_979)
);

OA21x2_ASAP7_75t_L g980 ( 
.A1(n_833),
.A2(n_660),
.B(n_658),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_866),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_821),
.A2(n_604),
.B1(n_715),
.B2(n_656),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_836),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_871),
.B(n_658),
.Y(n_984)
);

INVx6_ASAP7_75t_L g985 ( 
.A(n_901),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_789),
.B(n_752),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_882),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_797),
.B(n_755),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_875),
.B(n_660),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_867),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_836),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_802),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_843),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_SL g994 ( 
.A1(n_787),
.A2(n_744),
.B1(n_751),
.B2(n_693),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_803),
.A2(n_484),
.B1(n_486),
.B2(n_485),
.Y(n_995)
);

OA21x2_ASAP7_75t_L g996 ( 
.A1(n_843),
.A2(n_671),
.B(n_663),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_844),
.A2(n_671),
.B(n_663),
.Y(n_997)
);

NOR2x1_ASAP7_75t_L g998 ( 
.A(n_895),
.B(n_681),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_882),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_811),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_853),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_838),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_853),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_854),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_854),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_855),
.B(n_681),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_916),
.B(n_684),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_886),
.B(n_678),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_886),
.B(n_586),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_855),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_857),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_834),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_857),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_770),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_858),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_876),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_858),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_859),
.Y(n_1020)
);

INVx6_ASAP7_75t_L g1021 ( 
.A(n_883),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_SL g1022 ( 
.A(n_894),
.B(n_608),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_831),
.B(n_586),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_830),
.B(n_682),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_859),
.Y(n_1025)
);

INVx6_ASAP7_75t_L g1026 ( 
.A(n_852),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_860),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_845),
.B(n_851),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_860),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_861),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_770),
.Y(n_1031)
);

CKINVDCx6p67_ASAP7_75t_R g1032 ( 
.A(n_906),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_861),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_864),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_864),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_879),
.A2(n_711),
.B1(n_548),
.B2(n_493),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_839),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_841),
.B(n_684),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_847),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_865),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_865),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_918),
.Y(n_1042)
);

OA21x2_ASAP7_75t_L g1043 ( 
.A1(n_923),
.A2(n_775),
.B(n_774),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_918),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_977),
.B(n_849),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_924),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_945),
.B(n_842),
.Y(n_1048)
);

OA21x2_ASAP7_75t_L g1049 ( 
.A1(n_923),
.A2(n_775),
.B(n_774),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_1018),
.B(n_870),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_924),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_925),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1004),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_925),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_929),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1032),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1026),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_969),
.A2(n_777),
.B(n_776),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_929),
.Y(n_1059)
);

INVx6_ASAP7_75t_L g1060 ( 
.A(n_1016),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_1016),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_1026),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1032),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1039),
.Y(n_1064)
);

CKINVDCx16_ASAP7_75t_R g1065 ( 
.A(n_952),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1004),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_917),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_976),
.B(n_543),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_1039),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_945),
.B(n_850),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_917),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_952),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_R g1073 ( 
.A(n_981),
.B(n_888),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_920),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_920),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_956),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_956),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_919),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_926),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_972),
.B(n_904),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1026),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1036),
.A2(n_909),
.B1(n_912),
.B2(n_911),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_992),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_945),
.B(n_946),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_977),
.B(n_962),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_945),
.B(n_878),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_981),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_975),
.B(n_913),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_992),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_R g1090 ( 
.A(n_990),
.B(n_999),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1026),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_921),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_969),
.A2(n_777),
.B(n_776),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_921),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_961),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1014),
.B(n_889),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_929),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_961),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_939),
.B(n_848),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_927),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_927),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_967),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_978),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_990),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_934),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_999),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1008),
.A2(n_781),
.B(n_780),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_964),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1036),
.A2(n_491),
.B1(n_500),
.B2(n_499),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_967),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1021),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_934),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_964),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_978),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_962),
.B(n_869),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_978),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_978),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_931),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_962),
.B(n_869),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1014),
.A2(n_794),
.B1(n_745),
.B2(n_620),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_937),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_937),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_931),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1021),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_1023),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_940),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1010),
.B(n_880),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_940),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1021),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_929),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_944),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_944),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_962),
.B(n_970),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1021),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_970),
.B(n_872),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_947),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_985),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_947),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_960),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_971),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_929),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_935),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1010),
.B(n_881),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_935),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_960),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1001),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1037),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_949),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_949),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_953),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_953),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_965),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_968),
.B(n_884),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_965),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_986),
.B(n_988),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_935),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_954),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_946),
.B(n_685),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_946),
.B(n_685),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1037),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_971),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_968),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_966),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_966),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_954),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_974),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_963),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_973),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_R g1169 ( 
.A(n_1022),
.B(n_593),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1011),
.B(n_856),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_970),
.B(n_872),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_974),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_995),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_983),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_983),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_993),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_1028),
.B(n_633),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_970),
.B(n_873),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_933),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_933),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_982),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_935),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_982),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_993),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1002),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_946),
.B(n_873),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_994),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_973),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_985),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_991),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_985),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1002),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1013),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1013),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1015),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_935),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_950),
.B(n_874),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_R g1198 ( 
.A(n_1011),
.B(n_635),
.Y(n_1198)
);

AND3x2_ASAP7_75t_L g1199 ( 
.A(n_1023),
.B(n_540),
.C(n_496),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_938),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_950),
.B(n_874),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_985),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_932),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_950),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_976),
.B(n_891),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1008),
.A2(n_781),
.B(n_780),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_938),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_991),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1015),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1017),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_932),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_938),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_950),
.B(n_877),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1017),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_951),
.B(n_877),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_941),
.A2(n_501),
.B1(n_509),
.B2(n_506),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_976),
.B(n_914),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_976),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1020),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_984),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_984),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1020),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1029),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_951),
.B(n_640),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_951),
.B(n_726),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_984),
.Y(n_1226)
);

CKINVDCx16_ASAP7_75t_R g1227 ( 
.A(n_951),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1029),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_984),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_938),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1030),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_938),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1030),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1003),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1034),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_963),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_943),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1034),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_989),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1035),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_989),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1035),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_989),
.B(n_696),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_989),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1024),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1003),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1009),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1033),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1033),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1033),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_943),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1009),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1009),
.B(n_480),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_943),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_998),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1005),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1009),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_922),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1041),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1041),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1005),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1038),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1038),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_922),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1038),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_943),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1041),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1038),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1155),
.B(n_998),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1217),
.Y(n_1270)
);

INVxp33_ASAP7_75t_L g1271 ( 
.A(n_1050),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1105),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1099),
.B(n_510),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1084),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1133),
.B(n_1016),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1227),
.B(n_659),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1084),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1217),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1084),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1170),
.B(n_664),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1244),
.B(n_1016),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1243),
.A2(n_959),
.B1(n_980),
.B2(n_922),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1046),
.B(n_1080),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1243),
.A2(n_959),
.B1(n_980),
.B2(n_922),
.Y(n_1284)
);

AND2x6_ASAP7_75t_L g1285 ( 
.A(n_1247),
.B(n_696),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1078),
.Y(n_1286)
);

INVx5_ASAP7_75t_L g1287 ( 
.A(n_1060),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1105),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1137),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1244),
.B(n_1016),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_1204),
.B(n_753),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1228),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1170),
.B(n_669),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1243),
.A2(n_980),
.B1(n_996),
.B2(n_959),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1228),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1158),
.A2(n_980),
.B1(n_996),
.B2(n_959),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1204),
.B(n_1016),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1218),
.A2(n_758),
.B1(n_753),
.B2(n_628),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1247),
.B(n_758),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1231),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1205),
.B(n_996),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1231),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1042),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1042),
.Y(n_1304)
);

OR2x6_ASAP7_75t_L g1305 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1085),
.B(n_1162),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1045),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1088),
.B(n_513),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1045),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1137),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1048),
.B(n_1031),
.Y(n_1311)
);

AND2x6_ASAP7_75t_L g1312 ( 
.A(n_1158),
.B(n_543),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1072),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1047),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1048),
.B(n_1031),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1205),
.Y(n_1316)
);

INVxp33_ASAP7_75t_L g1317 ( 
.A(n_1106),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1186),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1245),
.B(n_515),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1047),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1059),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1090),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1091),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1048),
.B(n_1031),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1159),
.A2(n_997),
.B1(n_996),
.B2(n_725),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1051),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1115),
.B(n_997),
.C(n_788),
.Y(n_1327)
);

OA22x2_ASAP7_75t_L g1328 ( 
.A1(n_1203),
.A2(n_553),
.B1(n_477),
.B2(n_495),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1043),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1218),
.B(n_1220),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1070),
.B(n_1031),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1051),
.Y(n_1332)
);

AND2x6_ASAP7_75t_L g1333 ( 
.A(n_1159),
.B(n_543),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1043),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1052),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_L g1336 ( 
.A(n_1082),
.B(n_1065),
.C(n_1096),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1197),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1245),
.B(n_516),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1052),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1070),
.B(n_1031),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1255),
.B(n_521),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1201),
.Y(n_1342)
);

AND2x6_ASAP7_75t_L g1343 ( 
.A(n_1070),
.B(n_543),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1127),
.B(n_997),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1054),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1054),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1076),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1086),
.B(n_1031),
.Y(n_1348)
);

INVx5_ASAP7_75t_L g1349 ( 
.A(n_1060),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1127),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1213),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1076),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1220),
.B(n_674),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1086),
.B(n_494),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1221),
.B(n_680),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_706),
.B1(n_709),
.B2(n_691),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1215),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1086),
.B(n_494),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1143),
.B(n_997),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1077),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1077),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1226),
.B(n_957),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1258),
.A2(n_725),
.B1(n_730),
.B2(n_682),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1095),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1264),
.A2(n_714),
.B1(n_721),
.B2(n_710),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1095),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1226),
.B(n_1229),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1043),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1043),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1098),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1049),
.Y(n_1371)
);

NOR3xp33_ASAP7_75t_L g1372 ( 
.A(n_1109),
.B(n_525),
.C(n_524),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1229),
.B(n_957),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1068),
.A2(n_725),
.B1(n_730),
.B2(n_682),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1125),
.B(n_592),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1098),
.Y(n_1376)
);

CKINVDCx16_ASAP7_75t_R g1377 ( 
.A(n_1073),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1102),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1083),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1102),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1110),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1110),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1140),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1140),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1161),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1161),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1091),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1168),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1059),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1239),
.B(n_728),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1064),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1059),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1179),
.A2(n_507),
.B1(n_550),
.B2(n_471),
.Y(n_1393)
);

AND3x2_ASAP7_75t_L g1394 ( 
.A(n_1211),
.B(n_540),
.C(n_496),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1239),
.B(n_738),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1241),
.A2(n_1252),
.B1(n_1262),
.B2(n_1257),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1057),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1049),
.Y(n_1398)
);

AND2x2_ASAP7_75t_SL g1399 ( 
.A(n_1049),
.B(n_572),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1168),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1188),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1188),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1108),
.B(n_592),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1190),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1241),
.B(n_1198),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1190),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1208),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1208),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1216),
.B(n_530),
.C(n_529),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1143),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1062),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1234),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1234),
.Y(n_1413)
);

AND2x6_ASAP7_75t_L g1414 ( 
.A(n_1153),
.B(n_572),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1060),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1153),
.B(n_957),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1119),
.B(n_957),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1246),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1246),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1135),
.B(n_957),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1064),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1107),
.A2(n_788),
.B(n_782),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1068),
.A2(n_1178),
.B1(n_1171),
.B2(n_1101),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1256),
.Y(n_1424)
);

INVx4_ASAP7_75t_L g1425 ( 
.A(n_1059),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1256),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1100),
.B(n_958),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1112),
.B(n_958),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1261),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1261),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1108),
.B(n_1113),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1068),
.A2(n_1122),
.B1(n_1126),
.B2(n_1121),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1059),
.Y(n_1433)
);

AND2x6_ASAP7_75t_L g1434 ( 
.A(n_1053),
.B(n_1066),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1049),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1068),
.A2(n_730),
.B1(n_725),
.B2(n_958),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1058),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1255),
.B(n_533),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1113),
.B(n_1147),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1058),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1068),
.A2(n_730),
.B1(n_725),
.B2(n_958),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1147),
.B(n_743),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1058),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1079),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1253),
.B(n_695),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1128),
.B(n_958),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1104),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1058),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1253),
.B(n_782),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1097),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1160),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1160),
.B(n_1252),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1067),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1189),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1093),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1173),
.A2(n_768),
.B1(n_749),
.B2(n_539),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1093),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1093),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1189),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1263),
.A2(n_590),
.B1(n_572),
.B2(n_791),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1071),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1263),
.B(n_805),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1097),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1093),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1074),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1131),
.B(n_987),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1097),
.Y(n_1468)
);

AND2x6_ASAP7_75t_L g1469 ( 
.A(n_1248),
.B(n_572),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1132),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1136),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1055),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1081),
.B(n_537),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1075),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1138),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1092),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1094),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1249),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1148),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1120),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1265),
.A2(n_1268),
.B1(n_1173),
.B2(n_1177),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1191),
.Y(n_1482)
);

AND3x2_ASAP7_75t_L g1483 ( 
.A(n_1149),
.B(n_623),
.C(n_607),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1250),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1265),
.B(n_541),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1259),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1268),
.B(n_572),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1260),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1225),
.B(n_542),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1150),
.B(n_987),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1267),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1151),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1152),
.B(n_791),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1154),
.B(n_987),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1068),
.A2(n_730),
.B1(n_725),
.B2(n_987),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1163),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1055),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1164),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1166),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1172),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1174),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1191),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1202),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_SL g1504 ( 
.A(n_1169),
.B(n_565),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1175),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1202),
.B(n_544),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1176),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1199),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1179),
.B(n_695),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1111),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1184),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1185),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_L g1513 ( 
.A(n_1068),
.B(n_705),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1224),
.B(n_572),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1192),
.B(n_987),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1468),
.Y(n_1516)
);

NAND3x1_ASAP7_75t_L g1517 ( 
.A(n_1336),
.B(n_1372),
.C(n_1456),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1274),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1316),
.B(n_1305),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1269),
.B(n_1193),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1316),
.B(n_1194),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1305),
.B(n_1195),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1273),
.B(n_1209),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1277),
.B(n_1274),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1274),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1431),
.B(n_1069),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1279),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1403),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1279),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1272),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1468),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1363),
.B(n_1124),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1272),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1277),
.B(n_1146),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1510),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1277),
.B(n_1283),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1295),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1295),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1303),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1449),
.B(n_1210),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1303),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1379),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1288),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1304),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1288),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1431),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1304),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1350),
.B(n_1069),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1449),
.B(n_1214),
.Y(n_1549)
);

AO22x2_ASAP7_75t_L g1550 ( 
.A1(n_1480),
.A2(n_498),
.B1(n_508),
.B2(n_495),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1318),
.B(n_1219),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1307),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1305),
.B(n_1222),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1307),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1451),
.Y(n_1555)
);

OR2x2_ASAP7_75t_SL g1556 ( 
.A(n_1377),
.B(n_1180),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1292),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1292),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1318),
.B(n_1223),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1270),
.A2(n_1181),
.B1(n_1146),
.B2(n_1187),
.Y(n_1560)
);

INVx4_ASAP7_75t_SL g1561 ( 
.A(n_1285),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1350),
.B(n_1124),
.Y(n_1562)
);

BUFx4f_ASAP7_75t_L g1563 ( 
.A(n_1286),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1300),
.Y(n_1564)
);

AO22x2_ASAP7_75t_L g1565 ( 
.A1(n_1509),
.A2(n_508),
.B1(n_511),
.B2(n_498),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1322),
.B(n_1181),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1300),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1302),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_L g1569 ( 
.A(n_1323),
.B(n_1083),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1309),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1410),
.B(n_1129),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1305),
.B(n_1270),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1310),
.B(n_1107),
.Y(n_1573)
);

AO22x2_ASAP7_75t_L g1574 ( 
.A1(n_1509),
.A2(n_511),
.B1(n_520),
.B2(n_519),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1309),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1305),
.B(n_1233),
.Y(n_1576)
);

OAI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1410),
.A2(n_1187),
.B1(n_1183),
.B2(n_1165),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1510),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1403),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1439),
.B(n_1129),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1302),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1278),
.B(n_1235),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1278),
.B(n_1238),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1319),
.B(n_1044),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1338),
.B(n_1044),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1478),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1341),
.B(n_1438),
.Y(n_1587)
);

OR2x2_ASAP7_75t_SL g1588 ( 
.A(n_1377),
.B(n_1139),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1314),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1306),
.B(n_1165),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1314),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1306),
.B(n_1103),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1337),
.B(n_1240),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1310),
.B(n_1206),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1478),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1468),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1484),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1484),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1468),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1337),
.B(n_1242),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1498),
.A2(n_1114),
.B1(n_1116),
.B2(n_1103),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1468),
.Y(n_1602)
);

OAI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1365),
.A2(n_1116),
.B1(n_1117),
.B2(n_1114),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1320),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1447),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1320),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1447),
.B(n_1056),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1313),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1486),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1506),
.B(n_1117),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1342),
.B(n_1206),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1289),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1289),
.B(n_1354),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1379),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1351),
.B(n_1212),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1472),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1444),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1445),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1310),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1291),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1310),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1357),
.B(n_1212),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1326),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1354),
.B(n_1134),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1354),
.B(n_1055),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1486),
.Y(n_1627)
);

OAI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1456),
.A2(n_520),
.B1(n_536),
.B2(n_527),
.C(n_519),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1472),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1488),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1393),
.A2(n_1308),
.B1(n_1409),
.B2(n_1489),
.C(n_1365),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1326),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1488),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1444),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1491),
.Y(n_1635)
);

INVx8_ASAP7_75t_L g1636 ( 
.A(n_1285),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1491),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1367),
.B(n_1056),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1454),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1360),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1360),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1332),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1354),
.B(n_1358),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1286),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1358),
.B(n_1130),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1357),
.B(n_1399),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1498),
.B(n_1251),
.Y(n_1647)
);

INVx4_ASAP7_75t_SL g1648 ( 
.A(n_1285),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1358),
.B(n_1130),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1399),
.B(n_1097),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1387),
.B(n_1063),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1361),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1399),
.B(n_1097),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1358),
.B(n_1130),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1361),
.Y(n_1655)
);

AO22x2_ASAP7_75t_L g1656 ( 
.A1(n_1299),
.A2(n_527),
.B1(n_546),
.B2(n_536),
.Y(n_1656)
);

AO22x2_ASAP7_75t_L g1657 ( 
.A1(n_1299),
.A2(n_546),
.B1(n_574),
.B2(n_564),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1310),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1364),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1391),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1364),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1472),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1370),
.Y(n_1663)
);

OR2x2_ASAP7_75t_SL g1664 ( 
.A(n_1375),
.B(n_1139),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1450),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1370),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1376),
.Y(n_1667)
);

AO22x2_ASAP7_75t_L g1668 ( 
.A1(n_1299),
.A2(n_574),
.B1(n_582),
.B2(n_564),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1391),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1376),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1454),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1378),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1378),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1460),
.B(n_1141),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1499),
.B(n_1501),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1332),
.Y(n_1676)
);

AO22x2_ASAP7_75t_L g1677 ( 
.A1(n_1299),
.A2(n_599),
.B1(n_610),
.B2(n_582),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1497),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1291),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1499),
.B(n_1200),
.Y(n_1680)
);

AND2x6_ASAP7_75t_L g1681 ( 
.A(n_1435),
.B(n_590),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1381),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1381),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1501),
.B(n_1200),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1335),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1470),
.B(n_1141),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1460),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1383),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1301),
.B(n_1142),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1317),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1375),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1383),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1301),
.A2(n_1157),
.B1(n_1141),
.B2(n_1156),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1335),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1482),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1452),
.B(n_1063),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1485),
.B(n_1089),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1386),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1339),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1386),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1482),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1334),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1388),
.Y(n_1703)
);

AND2x6_ASAP7_75t_L g1704 ( 
.A(n_1435),
.B(n_590),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1445),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1502),
.B(n_1089),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1339),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1388),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1271),
.B(n_1144),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1400),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1473),
.B(n_1087),
.C(n_1145),
.Y(n_1711)
);

AO22x2_ASAP7_75t_L g1712 ( 
.A1(n_1459),
.A2(n_610),
.B1(n_614),
.B2(n_599),
.Y(n_1712)
);

AO22x2_ASAP7_75t_L g1713 ( 
.A1(n_1459),
.A2(n_614),
.B1(n_624),
.B2(n_616),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1505),
.B(n_1251),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1505),
.B(n_1512),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1450),
.Y(n_1716)
);

INVx6_ASAP7_75t_L g1717 ( 
.A(n_1391),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1400),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1470),
.B(n_1144),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1512),
.B(n_1251),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1502),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1345),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1401),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1280),
.B(n_1118),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1345),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1401),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1402),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1344),
.B(n_1142),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1330),
.B(n_1144),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1402),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1346),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1346),
.Y(n_1732)
);

INVx5_ASAP7_75t_L g1733 ( 
.A(n_1334),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1450),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1413),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1344),
.B(n_1142),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1347),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1321),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1396),
.B(n_1156),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1471),
.B(n_1156),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1421),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1413),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1481),
.B(n_1200),
.Y(n_1743)
);

INVx4_ASAP7_75t_SL g1744 ( 
.A(n_1285),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1453),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1503),
.B(n_1212),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1450),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1453),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1497),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1462),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1347),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1462),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1321),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1359),
.A2(n_624),
.B1(n_626),
.B2(n_616),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1466),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1497),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1352),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1466),
.Y(n_1758)
);

OAI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1328),
.A2(n_730),
.B1(n_701),
.B2(n_623),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1474),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1334),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1293),
.A2(n_665),
.B1(n_676),
.B2(n_630),
.C(n_626),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1546),
.B(n_1397),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1733),
.B(n_1587),
.Y(n_1764)
);

AO22x1_ASAP7_75t_L g1765 ( 
.A1(n_1584),
.A2(n_1145),
.B1(n_1087),
.B2(n_1123),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1530),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1607),
.B(n_1492),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1523),
.B(n_1492),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1687),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1530),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1631),
.A2(n_1503),
.B1(n_1421),
.B2(n_1087),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1562),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1517),
.A2(n_1405),
.B1(n_1463),
.B2(n_1504),
.Y(n_1774)
);

NAND2x1p5_ASAP7_75t_L g1775 ( 
.A(n_1733),
.B(n_1321),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1566),
.B(n_1411),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1733),
.B(n_1518),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1532),
.A2(n_1291),
.B1(n_1285),
.B2(n_1471),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1533),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1532),
.A2(n_1291),
.B1(n_1285),
.B2(n_1475),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1733),
.B(n_1511),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1533),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1643),
.A2(n_1291),
.B1(n_1285),
.B2(n_1475),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1761),
.Y(n_1785)
);

AND2x6_ASAP7_75t_SL g1786 ( 
.A(n_1696),
.B(n_630),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1687),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1517),
.A2(n_1355),
.B1(n_1390),
.B2(n_1353),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1695),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1560),
.A2(n_1496),
.B1(n_1500),
.B2(n_1479),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1551),
.B(n_1500),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1536),
.A2(n_1392),
.B(n_1389),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1518),
.B(n_1507),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1643),
.A2(n_1507),
.B1(n_1511),
.B2(n_1479),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1543),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1761),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1572),
.B(n_1474),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1691),
.B(n_1476),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1526),
.B(n_1421),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1536),
.A2(n_1392),
.B(n_1389),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1559),
.B(n_1476),
.Y(n_1801)
);

NOR2xp67_ASAP7_75t_L g1802 ( 
.A(n_1711),
.B(n_1118),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1593),
.B(n_1477),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1600),
.B(n_1477),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1605),
.B(n_1442),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1539),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1542),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_SL g1808 ( 
.A1(n_1743),
.A2(n_1422),
.B(n_1423),
.C(n_1282),
.Y(n_1808)
);

BUFx4f_ASAP7_75t_L g1809 ( 
.A(n_1660),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1556),
.A2(n_1123),
.B1(n_1508),
.B2(n_571),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1518),
.B(n_1362),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1585),
.B(n_1328),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1539),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1545),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1540),
.B(n_1493),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1557),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1541),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1541),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_L g1819 ( 
.A1(n_1638),
.A2(n_1328),
.B(n_1395),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1558),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1564),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1549),
.B(n_1493),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1516),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1675),
.B(n_1359),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1643),
.A2(n_1487),
.B1(n_1416),
.B2(n_1373),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1646),
.A2(n_1653),
.B(n_1650),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1690),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1715),
.B(n_1334),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1544),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1695),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1628),
.A2(n_1298),
.B(n_1276),
.C(n_1356),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1544),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1646),
.A2(n_1432),
.B1(n_1325),
.B2(n_1368),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1567),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1638),
.A2(n_1508),
.B1(n_1434),
.B2(n_1514),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1542),
.A2(n_1615),
.B1(n_1609),
.B2(n_1669),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1516),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1745),
.B(n_1448),
.Y(n_1838)
);

INVxp67_ASAP7_75t_SL g1839 ( 
.A(n_1761),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1748),
.B(n_1448),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1738),
.B(n_1389),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1568),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1525),
.B(n_1281),
.Y(n_1843)
);

BUFx12f_ASAP7_75t_L g1844 ( 
.A(n_1644),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1547),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1702),
.A2(n_1650),
.B1(n_1653),
.B2(n_1761),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1525),
.B(n_1290),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1572),
.A2(n_1434),
.B1(n_1343),
.B2(n_1312),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1548),
.B(n_1394),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1750),
.B(n_1368),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1738),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1581),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1572),
.A2(n_1434),
.B1(n_1343),
.B2(n_1312),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1752),
.B(n_1368),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1755),
.A2(n_1334),
.B1(n_1369),
.B2(n_1368),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1701),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1614),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1525),
.B(n_1297),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1537),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1758),
.B(n_1368),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1618),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1760),
.B(n_1369),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1580),
.B(n_1483),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1592),
.B(n_1590),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1521),
.B(n_1369),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1738),
.Y(n_1866)
);

NOR3xp33_ASAP7_75t_L g1867 ( 
.A(n_1697),
.B(n_1324),
.C(n_1315),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1555),
.B(n_1369),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1538),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1519),
.B(n_1275),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1639),
.Y(n_1871)
);

BUFx5_ASAP7_75t_L g1872 ( 
.A(n_1681),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1547),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1615),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1640),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1521),
.B(n_1369),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1521),
.B(n_1398),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1689),
.A2(n_1327),
.B(n_1417),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1641),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1586),
.B(n_1398),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1595),
.B(n_1398),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1528),
.B(n_1398),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1696),
.B(n_1513),
.C(n_551),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1634),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1701),
.Y(n_1886)
);

OR2x6_ASAP7_75t_L g1887 ( 
.A(n_1519),
.B(n_1398),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1519),
.A2(n_1434),
.B1(n_1343),
.B2(n_1312),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1610),
.B(n_1448),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1611),
.A2(n_1461),
.B1(n_1434),
.B2(n_1333),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1552),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1627),
.B(n_1448),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1614),
.B(n_1352),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1522),
.B(n_1434),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1630),
.B(n_1448),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1614),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1579),
.B(n_1440),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1633),
.B(n_1366),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1516),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1693),
.A2(n_1443),
.B1(n_1455),
.B2(n_1440),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1552),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1619),
.B(n_1443),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1635),
.B(n_1366),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1753),
.B(n_1380),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1626),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1637),
.B(n_1380),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1626),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1705),
.B(n_507),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1609),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1554),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1582),
.B(n_1382),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1651),
.B(n_507),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1621),
.A2(n_1457),
.B1(n_1458),
.B2(n_1455),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1644),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1554),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1753),
.B(n_1382),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1652),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1753),
.B(n_1384),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1582),
.B(n_1384),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1535),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_SL g1921 ( 
.A(n_1706),
.B(n_1434),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1582),
.B(n_1385),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1671),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1571),
.A2(n_1331),
.B1(n_1340),
.B2(n_1311),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1583),
.B(n_1385),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1617),
.B(n_1404),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1570),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1583),
.B(n_1404),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1655),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1583),
.B(n_1406),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1721),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1721),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1608),
.B(n_1406),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1709),
.B(n_1407),
.Y(n_1935)
);

INVx3_ASAP7_75t_L g1936 ( 
.A(n_1658),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1762),
.A2(n_560),
.B1(n_562),
.B2(n_554),
.C(n_545),
.Y(n_1937)
);

NAND2x1p5_ASAP7_75t_L g1938 ( 
.A(n_1658),
.B(n_1596),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1535),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1659),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1709),
.B(n_1407),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1570),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1661),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1658),
.Y(n_1944)
);

OR2x6_ASAP7_75t_L g1945 ( 
.A(n_1636),
.B(n_1457),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1578),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1669),
.A2(n_566),
.B1(n_606),
.B2(n_587),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1621),
.A2(n_1343),
.B1(n_1333),
.B2(n_1312),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1746),
.B(n_1408),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1571),
.A2(n_1348),
.B1(n_1343),
.B2(n_1427),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1626),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1578),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1575),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1625),
.B(n_507),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1575),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1617),
.B(n_1408),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1663),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1589),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1746),
.B(n_1412),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1759),
.B(n_1412),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1617),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1666),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1759),
.B(n_1418),
.Y(n_1963)
);

A2O1A1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1754),
.A2(n_1327),
.B(n_1374),
.C(n_1284),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_SL g1965 ( 
.A(n_1741),
.B(n_550),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1754),
.B(n_1418),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1729),
.B(n_1419),
.Y(n_1967)
);

OAI22xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1534),
.A2(n_1724),
.B1(n_1660),
.B2(n_1717),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1729),
.B(n_1419),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1667),
.B(n_1424),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1534),
.A2(n_1343),
.B1(n_1446),
.B2(n_1428),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1670),
.B(n_1672),
.Y(n_1972)
);

INVx5_ASAP7_75t_L g1973 ( 
.A(n_1636),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1679),
.A2(n_1343),
.B1(n_1490),
.B2(n_1467),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1673),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1797),
.B(n_1613),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1795),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1769),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1814),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1864),
.A2(n_1625),
.B1(n_1577),
.B2(n_1569),
.Y(n_1980)
);

AND3x1_ASAP7_75t_SL g1981 ( 
.A(n_1937),
.B(n_676),
.C(n_665),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1887),
.Y(n_1982)
);

INVx5_ASAP7_75t_L g1983 ( 
.A(n_1887),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1861),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1797),
.B(n_1613),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1768),
.B(n_1679),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1801),
.B(n_1522),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1816),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1887),
.B(n_1660),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1766),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1766),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1887),
.B(n_1894),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1788),
.A2(n_1625),
.B1(n_1577),
.B2(n_1553),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1779),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1803),
.B(n_1522),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1823),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1804),
.B(n_1553),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1781),
.B(n_1601),
.Y(n_1998)
);

INVx4_ASAP7_75t_L g1999 ( 
.A(n_1809),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1884),
.Y(n_2000)
);

NOR2xp67_ASAP7_75t_L g2001 ( 
.A(n_1807),
.B(n_1743),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1823),
.Y(n_2002)
);

NOR3xp33_ASAP7_75t_SL g2003 ( 
.A(n_1819),
.B(n_1601),
.C(n_1739),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_R g2004 ( 
.A(n_1807),
.B(n_1717),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1799),
.B(n_1565),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1779),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1815),
.B(n_1603),
.Y(n_2007)
);

INVx5_ASAP7_75t_L g2008 ( 
.A(n_1945),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1827),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1909),
.Y(n_2010)
);

OR2x6_ASAP7_75t_L g2011 ( 
.A(n_1894),
.B(n_1717),
.Y(n_2011)
);

INVx1_ASAP7_75t_SL g2012 ( 
.A(n_1871),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1822),
.B(n_1553),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1797),
.B(n_1576),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1865),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1769),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1894),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1783),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1820),
.Y(n_2019)
);

AND3x1_ASAP7_75t_SL g2020 ( 
.A(n_1786),
.B(n_697),
.C(n_679),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1851),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1772),
.B(n_1576),
.Y(n_2022)
);

BUFx12f_ASAP7_75t_L g2023 ( 
.A(n_1909),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1787),
.Y(n_2024)
);

AND2x6_ASAP7_75t_SL g2025 ( 
.A(n_1776),
.B(n_1739),
.Y(n_2025)
);

INVx4_ASAP7_75t_L g2026 ( 
.A(n_1809),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1851),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1781),
.B(n_1576),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1851),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1787),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1783),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1767),
.B(n_1773),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1812),
.B(n_1912),
.Y(n_2033)
);

AOI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1776),
.A2(n_1563),
.B1(n_1649),
.B2(n_1645),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1773),
.B(n_1712),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1874),
.Y(n_2036)
);

BUFx4f_ASAP7_75t_SL g2037 ( 
.A(n_1844),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1821),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1834),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1789),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_SL g2041 ( 
.A(n_1810),
.B(n_568),
.C(n_563),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1874),
.Y(n_2042)
);

AND2x4_ASAP7_75t_SL g2043 ( 
.A(n_1946),
.B(n_1620),
.Y(n_2043)
);

BUFx12f_ASAP7_75t_L g2044 ( 
.A(n_1844),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1774),
.A2(n_1563),
.B1(n_1649),
.B2(n_1645),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1763),
.B(n_1664),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1789),
.B(n_1830),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1798),
.B(n_1588),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1791),
.B(n_1712),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1868),
.B(n_1798),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1876),
.Y(n_2051)
);

NOR3xp33_ASAP7_75t_L g2052 ( 
.A(n_1771),
.B(n_1831),
.C(n_1968),
.Y(n_2052)
);

AND3x2_ASAP7_75t_SL g2053 ( 
.A(n_1806),
.B(n_1713),
.C(n_1712),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1806),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1868),
.B(n_1713),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_R g2056 ( 
.A(n_1914),
.B(n_1636),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1813),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1934),
.B(n_1805),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_R g2059 ( 
.A(n_1914),
.B(n_1830),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_SL g2060 ( 
.A(n_1835),
.B(n_1674),
.C(n_1524),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1842),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1852),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1875),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1794),
.A2(n_1674),
.B1(n_1683),
.B2(n_1682),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_1947),
.B(n_573),
.C(n_569),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1856),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1856),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1813),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1886),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1879),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1917),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1923),
.B(n_1688),
.Y(n_2072)
);

AND3x1_ASAP7_75t_SL g2073 ( 
.A(n_1929),
.B(n_697),
.C(n_679),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1790),
.B(n_1692),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1866),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1817),
.Y(n_2076)
);

BUFx4f_ASAP7_75t_L g2077 ( 
.A(n_1849),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1817),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1886),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1863),
.A2(n_1645),
.B1(n_1654),
.B2(n_1649),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1885),
.B(n_1713),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1818),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1877),
.Y(n_2083)
);

BUFx12f_ASAP7_75t_L g2084 ( 
.A(n_1920),
.Y(n_2084)
);

NOR3xp33_ASAP7_75t_SL g2085 ( 
.A(n_1836),
.B(n_579),
.C(n_576),
.Y(n_2085)
);

OR2x6_ASAP7_75t_L g2086 ( 
.A(n_1857),
.B(n_1654),
.Y(n_2086)
);

BUFx12f_ASAP7_75t_L g2087 ( 
.A(n_1939),
.Y(n_2087)
);

OR2x6_ASAP7_75t_L g2088 ( 
.A(n_1857),
.B(n_1654),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1823),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1896),
.B(n_1620),
.Y(n_2090)
);

INVx8_ASAP7_75t_L g2091 ( 
.A(n_1823),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_1931),
.B(n_1698),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_1933),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_SL g2094 ( 
.A(n_1764),
.B(n_1883),
.C(n_584),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1837),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1818),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1829),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_1785),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1954),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1824),
.B(n_1656),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1940),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1943),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_1896),
.B(n_1561),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1837),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1932),
.B(n_1656),
.Y(n_2105)
);

A2O1A1Ixp33_ASAP7_75t_L g2106 ( 
.A1(n_1964),
.A2(n_1703),
.B(n_1708),
.C(n_1700),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1957),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1952),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1902),
.B(n_1710),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1828),
.B(n_1656),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1837),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1792),
.A2(n_1594),
.B(n_1573),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1908),
.B(n_1962),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1808),
.A2(n_1612),
.B(n_1420),
.Y(n_2114)
);

BUFx2_ASAP7_75t_L g2115 ( 
.A(n_1905),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1975),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1829),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1859),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1905),
.B(n_1907),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1869),
.Y(n_2120)
);

NOR3xp33_ASAP7_75t_SL g2121 ( 
.A(n_1764),
.B(n_589),
.C(n_581),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_1785),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1866),
.Y(n_2123)
);

NOR2x1_ASAP7_75t_L g2124 ( 
.A(n_1882),
.B(n_1596),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1832),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1770),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1832),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1902),
.B(n_1718),
.Y(n_2128)
);

CKINVDCx16_ASAP7_75t_R g2129 ( 
.A(n_1965),
.Y(n_2129)
);

INVx1_ASAP7_75t_SL g2130 ( 
.A(n_1911),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1845),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1866),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1845),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1873),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_R g2135 ( 
.A(n_1921),
.B(n_1629),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1897),
.B(n_1723),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1873),
.Y(n_2137)
);

OR2x6_ASAP7_75t_L g2138 ( 
.A(n_1907),
.B(n_1620),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1891),
.Y(n_2139)
);

BUFx4f_ASAP7_75t_L g2140 ( 
.A(n_1837),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1891),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1890),
.B(n_1726),
.Y(n_2142)
);

NOR3xp33_ASAP7_75t_SL g2143 ( 
.A(n_1870),
.B(n_597),
.C(n_594),
.Y(n_2143)
);

AND2x6_ASAP7_75t_L g2144 ( 
.A(n_1936),
.B(n_1629),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1867),
.B(n_1727),
.Y(n_2145)
);

BUFx4f_ASAP7_75t_L g2146 ( 
.A(n_1899),
.Y(n_2146)
);

BUFx4f_ASAP7_75t_L g2147 ( 
.A(n_1899),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1897),
.B(n_1657),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_1951),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1778),
.B(n_1730),
.Y(n_2150)
);

AOI211xp5_ASAP7_75t_L g2151 ( 
.A1(n_1765),
.A2(n_704),
.B(n_708),
.C(n_699),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1951),
.A2(n_1524),
.B1(n_1574),
.B2(n_1565),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1882),
.B(n_1657),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1901),
.Y(n_2154)
);

CKINVDCx20_ASAP7_75t_R g2155 ( 
.A(n_1899),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1899),
.Y(n_2156)
);

OR2x6_ASAP7_75t_L g2157 ( 
.A(n_1945),
.B(n_1620),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1972),
.B(n_1668),
.Y(n_2158)
);

BUFx5_ASAP7_75t_L g2159 ( 
.A(n_1872),
.Y(n_2159)
);

INVx4_ASAP7_75t_L g2160 ( 
.A(n_1936),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1901),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1919),
.B(n_1565),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1910),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1922),
.B(n_1735),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1910),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_1785),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1925),
.B(n_1574),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_1973),
.B(n_1945),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1928),
.B(n_1574),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1780),
.B(n_1742),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1973),
.B(n_1561),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1915),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_1945),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1915),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_1796),
.Y(n_2175)
);

NAND2xp33_ASAP7_75t_SL g2176 ( 
.A(n_1833),
.B(n_1516),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1808),
.A2(n_1612),
.B(n_1689),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1936),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1825),
.B(n_1826),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1930),
.B(n_1657),
.Y(n_2180)
);

INVxp67_ASAP7_75t_SL g2181 ( 
.A(n_1855),
.Y(n_2181)
);

INVx2_ASAP7_75t_SL g2182 ( 
.A(n_1893),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1944),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1927),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1935),
.B(n_1668),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_1838),
.B(n_1616),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1941),
.B(n_1668),
.Y(n_2187)
);

BUFx3_ASAP7_75t_L g2188 ( 
.A(n_1938),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1927),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_SL g2190 ( 
.A1(n_1784),
.A2(n_600),
.B1(n_605),
.B2(n_601),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1938),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1942),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_1973),
.B(n_1944),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_R g2194 ( 
.A(n_1944),
.B(n_1629),
.Y(n_2194)
);

OAI221xp5_ASAP7_75t_L g2195 ( 
.A1(n_1802),
.A2(n_708),
.B1(n_713),
.B2(n_704),
.C(n_699),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1973),
.B(n_1561),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1942),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1953),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1967),
.B(n_1677),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1953),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1973),
.Y(n_2201)
);

NOR3xp33_ASAP7_75t_SL g2202 ( 
.A(n_1870),
.B(n_611),
.C(n_609),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1955),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1893),
.B(n_1550),
.Y(n_2204)
);

OAI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_2007),
.A2(n_1924),
.B(n_1811),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2058),
.B(n_1677),
.Y(n_2206)
);

NAND2x1p5_ASAP7_75t_L g2207 ( 
.A(n_1983),
.B(n_1777),
.Y(n_2207)
);

NOR2x1_ASAP7_75t_L g2208 ( 
.A(n_1999),
.B(n_1961),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_2112),
.A2(n_1800),
.B(n_1843),
.Y(n_2209)
);

AO31x2_ASAP7_75t_L g2210 ( 
.A1(n_2114),
.A2(n_1846),
.A3(n_1913),
.B(n_1900),
.Y(n_2210)
);

AOI21x1_ASAP7_75t_SL g2211 ( 
.A1(n_2100),
.A2(n_2187),
.B(n_2185),
.Y(n_2211)
);

OAI21x1_ASAP7_75t_L g2212 ( 
.A1(n_2114),
.A2(n_1847),
.B(n_1843),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2058),
.B(n_1677),
.Y(n_2213)
);

NAND2x1p5_ASAP7_75t_L g2214 ( 
.A(n_1983),
.B(n_1777),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1977),
.Y(n_2215)
);

AND2x6_ASAP7_75t_L g2216 ( 
.A(n_2168),
.B(n_1961),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2050),
.B(n_2130),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2176),
.A2(n_1964),
.B(n_1878),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1992),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1979),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_1998),
.A2(n_1853),
.B1(n_1848),
.B2(n_1888),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2028),
.B(n_1550),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1990),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2059),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1998),
.A2(n_2001),
.B1(n_2048),
.B2(n_1993),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2032),
.B(n_1550),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2177),
.A2(n_1858),
.B(n_1847),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_2091),
.Y(n_2228)
);

OAI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_2007),
.A2(n_1811),
.B(n_1971),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1992),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1986),
.B(n_1955),
.Y(n_2231)
);

INVxp67_ASAP7_75t_SL g2232 ( 
.A(n_2015),
.Y(n_2232)
);

AO31x2_ASAP7_75t_L g2233 ( 
.A1(n_2177),
.A2(n_1969),
.A3(n_1963),
.B(n_1960),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1988),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_2052),
.B(n_1974),
.Y(n_2235)
);

AO31x2_ASAP7_75t_L g2236 ( 
.A1(n_2106),
.A2(n_1959),
.A3(n_1949),
.B(n_1966),
.Y(n_2236)
);

NAND2x1p5_ASAP7_75t_L g2237 ( 
.A(n_1983),
.B(n_2008),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1987),
.B(n_1958),
.Y(n_2238)
);

OAI21x1_ASAP7_75t_L g2239 ( 
.A1(n_2145),
.A2(n_1858),
.B(n_1594),
.Y(n_2239)
);

AOI211x1_ASAP7_75t_L g2240 ( 
.A1(n_2035),
.A2(n_720),
.B(n_723),
.C(n_713),
.Y(n_2240)
);

A2O1A1Ixp33_ASAP7_75t_L g2241 ( 
.A1(n_2003),
.A2(n_1850),
.B(n_1854),
.C(n_1840),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2176),
.A2(n_2179),
.B(n_2060),
.Y(n_2242)
);

OAI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_2145),
.A2(n_1950),
.B(n_1793),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1991),
.Y(n_2244)
);

A2O1A1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_2003),
.A2(n_1889),
.B(n_1862),
.C(n_1880),
.Y(n_2245)
);

AO31x2_ASAP7_75t_L g2246 ( 
.A1(n_2106),
.A2(n_1860),
.A3(n_1892),
.B(n_1881),
.Y(n_2246)
);

NOR2x1_ASAP7_75t_SL g2247 ( 
.A(n_1983),
.B(n_1782),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_2140),
.Y(n_2248)
);

AOI21x1_ASAP7_75t_L g2249 ( 
.A1(n_2179),
.A2(n_1916),
.B(n_1904),
.Y(n_2249)
);

OAI21x1_ASAP7_75t_L g2250 ( 
.A1(n_2074),
.A2(n_1573),
.B(n_1926),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2060),
.A2(n_1775),
.B(n_1904),
.Y(n_2251)
);

AOI21xp33_ASAP7_75t_L g2252 ( 
.A1(n_2049),
.A2(n_1793),
.B(n_1898),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2052),
.A2(n_1515),
.B(n_1494),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2142),
.A2(n_1775),
.B(n_1916),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2074),
.A2(n_1623),
.B(n_1647),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2036),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1995),
.B(n_1958),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1997),
.B(n_1872),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2142),
.A2(n_1918),
.B(n_1895),
.Y(n_2259)
);

AOI21x1_ASAP7_75t_L g2260 ( 
.A1(n_2150),
.A2(n_1918),
.B(n_1782),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2181),
.A2(n_1841),
.B(n_1839),
.Y(n_2261)
);

BUFx4f_ASAP7_75t_SL g2262 ( 
.A(n_2044),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2140),
.Y(n_2263)
);

AOI21x1_ASAP7_75t_SL g2264 ( 
.A1(n_2199),
.A2(n_1970),
.B(n_1906),
.Y(n_2264)
);

O2A1O1Ixp5_ASAP7_75t_L g2265 ( 
.A1(n_2150),
.A2(n_1956),
.B(n_1926),
.C(n_1736),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2019),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2038),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_2047),
.Y(n_2268)
);

AOI21x1_ASAP7_75t_SL g2269 ( 
.A1(n_2153),
.A2(n_1903),
.B(n_1684),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2170),
.A2(n_1956),
.B(n_1961),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2124),
.A2(n_1841),
.B(n_1714),
.Y(n_2271)
);

AOI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2181),
.A2(n_1596),
.B(n_1728),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2186),
.A2(n_1736),
.B(n_1728),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2033),
.B(n_1751),
.Y(n_2274)
);

AOI21x1_ASAP7_75t_L g2275 ( 
.A1(n_2170),
.A2(n_1720),
.B(n_1680),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2195),
.A2(n_701),
.B1(n_675),
.B2(n_550),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2021),
.A2(n_1678),
.B(n_1662),
.Y(n_2277)
);

OR2x6_ASAP7_75t_L g2278 ( 
.A(n_1989),
.B(n_2157),
.Y(n_2278)
);

OAI21x1_ASAP7_75t_L g2279 ( 
.A1(n_2021),
.A2(n_1678),
.B(n_1662),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_2047),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1994),
.Y(n_2281)
);

INVx4_ASAP7_75t_L g2282 ( 
.A(n_2091),
.Y(n_2282)
);

AO31x2_ASAP7_75t_L g2283 ( 
.A1(n_2186),
.A2(n_1589),
.A3(n_1604),
.B(n_1591),
.Y(n_2283)
);

OAI21x1_ASAP7_75t_L g2284 ( 
.A1(n_2027),
.A2(n_1678),
.B(n_1662),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2013),
.B(n_1591),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2146),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_2024),
.Y(n_2287)
);

AO21x1_ASAP7_75t_L g2288 ( 
.A1(n_2109),
.A2(n_1719),
.B(n_1686),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2022),
.A2(n_1425),
.B(n_1392),
.Y(n_2289)
);

O2A1O1Ixp5_ASAP7_75t_L g2290 ( 
.A1(n_2109),
.A2(n_2128),
.B(n_2136),
.C(n_2055),
.Y(n_2290)
);

NAND3x1_ASAP7_75t_L g2291 ( 
.A(n_1980),
.B(n_2048),
.C(n_2005),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2128),
.A2(n_1464),
.B(n_1425),
.Y(n_2292)
);

OAI21x1_ASAP7_75t_L g2293 ( 
.A1(n_2027),
.A2(n_1756),
.B(n_1749),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_1992),
.Y(n_2294)
);

O2A1O1Ixp5_ASAP7_75t_L g2295 ( 
.A1(n_2136),
.A2(n_1606),
.B(n_1624),
.C(n_1604),
.Y(n_2295)
);

AOI21xp33_ASAP7_75t_L g2296 ( 
.A1(n_2180),
.A2(n_2148),
.B(n_2110),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2162),
.B(n_1686),
.Y(n_2297)
);

AOI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_2193),
.A2(n_1464),
.B(n_1425),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2015),
.B(n_1732),
.Y(n_2299)
);

A2O1A1Ixp33_ASAP7_75t_L g2300 ( 
.A1(n_2195),
.A2(n_1513),
.B(n_639),
.C(n_646),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2046),
.A2(n_1719),
.B1(n_1740),
.B2(n_1686),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2039),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2051),
.B(n_2083),
.Y(n_2303)
);

A2O1A1Ixp33_ASAP7_75t_L g2304 ( 
.A1(n_2164),
.A2(n_639),
.B(n_646),
.C(n_607),
.Y(n_2304)
);

AOI21x1_ASAP7_75t_L g2305 ( 
.A1(n_2081),
.A2(n_1426),
.B(n_1424),
.Y(n_2305)
);

AOI21x1_ASAP7_75t_L g2306 ( 
.A1(n_2105),
.A2(n_1429),
.B(n_1426),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2051),
.B(n_1751),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_2025),
.B(n_1749),
.Y(n_2308)
);

CKINVDCx16_ASAP7_75t_R g2309 ( 
.A(n_2004),
.Y(n_2309)
);

OA22x2_ASAP7_75t_L g2310 ( 
.A1(n_2152),
.A2(n_723),
.B1(n_724),
.B2(n_720),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2168),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2083),
.B(n_1606),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2061),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2193),
.A2(n_1464),
.B(n_1433),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_2029),
.A2(n_1756),
.B(n_1749),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2099),
.B(n_1722),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2009),
.B(n_1722),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2143),
.B(n_1872),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2164),
.B(n_1725),
.Y(n_2319)
);

O2A1O1Ixp5_ASAP7_75t_L g2320 ( 
.A1(n_2158),
.A2(n_1632),
.B(n_1642),
.C(n_1624),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2146),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2064),
.A2(n_1433),
.B(n_1622),
.Y(n_2322)
);

OAI21x1_ASAP7_75t_L g2323 ( 
.A1(n_2029),
.A2(n_1756),
.B(n_1642),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2113),
.B(n_1725),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2167),
.B(n_1731),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2094),
.A2(n_1740),
.B(n_1719),
.Y(n_2326)
);

OAI21x1_ASAP7_75t_SL g2327 ( 
.A1(n_2045),
.A2(n_1948),
.B(n_1676),
.Y(n_2327)
);

AOI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2160),
.A2(n_1433),
.B(n_1622),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2062),
.Y(n_2329)
);

AO31x2_ASAP7_75t_L g2330 ( 
.A1(n_2127),
.A2(n_1632),
.A3(n_1685),
.B(n_1676),
.Y(n_2330)
);

OAI21x1_ASAP7_75t_L g2331 ( 
.A1(n_2075),
.A2(n_1694),
.B(n_1685),
.Y(n_2331)
);

A2O1A1Ixp33_ASAP7_75t_L g2332 ( 
.A1(n_2065),
.A2(n_654),
.B(n_698),
.C(n_647),
.Y(n_2332)
);

NAND2x1p5_ASAP7_75t_L g2333 ( 
.A(n_2008),
.B(n_1622),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_2075),
.A2(n_1699),
.B(n_1694),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2169),
.B(n_1757),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2063),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2014),
.B(n_1757),
.Y(n_2337)
);

O2A1O1Ixp5_ASAP7_75t_L g2338 ( 
.A1(n_2204),
.A2(n_1707),
.B(n_1731),
.C(n_1699),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_SL g2339 ( 
.A(n_2042),
.B(n_1622),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_1982),
.B(n_2017),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2014),
.B(n_1740),
.Y(n_2341)
);

OAI21x1_ASAP7_75t_L g2342 ( 
.A1(n_2123),
.A2(n_1732),
.B(n_1707),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2017),
.B(n_1737),
.Y(n_2343)
);

NOR2x1_ASAP7_75t_L g2344 ( 
.A(n_1999),
.B(n_1737),
.Y(n_2344)
);

OAI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2094),
.A2(n_1430),
.B(n_1429),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2006),
.Y(n_2346)
);

OA21x2_ASAP7_75t_L g2347 ( 
.A1(n_2126),
.A2(n_1294),
.B(n_1296),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2160),
.A2(n_2008),
.B(n_2157),
.Y(n_2348)
);

AOI21x1_ASAP7_75t_L g2349 ( 
.A1(n_2157),
.A2(n_1430),
.B(n_1458),
.Y(n_2349)
);

OAI21x1_ASAP7_75t_L g2350 ( 
.A1(n_2123),
.A2(n_1371),
.B(n_1329),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2059),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2132),
.A2(n_1982),
.B(n_2178),
.Y(n_2352)
);

AO21x1_ASAP7_75t_L g2353 ( 
.A1(n_2118),
.A2(n_2120),
.B(n_2071),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2132),
.A2(n_1371),
.B(n_1329),
.Y(n_2354)
);

AOI21xp33_ASAP7_75t_L g2355 ( 
.A1(n_2182),
.A2(n_2046),
.B(n_2034),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2178),
.A2(n_1371),
.B(n_1329),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2143),
.A2(n_1333),
.B(n_1312),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2070),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2098),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2072),
.B(n_612),
.Y(n_2360)
);

INVx3_ASAP7_75t_L g2361 ( 
.A(n_2171),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_L g2362 ( 
.A1(n_2183),
.A2(n_1465),
.B(n_1437),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2202),
.A2(n_1333),
.B(n_1312),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2202),
.B(n_2121),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_2067),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2072),
.B(n_613),
.Y(n_2366)
);

OAI22x1_ASAP7_75t_L g2367 ( 
.A1(n_2053),
.A2(n_731),
.B1(n_732),
.B2(n_724),
.Y(n_2367)
);

OAI22x1_ASAP7_75t_L g2368 ( 
.A1(n_2053),
.A2(n_732),
.B1(n_735),
.B2(n_731),
.Y(n_2368)
);

AOI221x1_ASAP7_75t_L g2369 ( 
.A1(n_2190),
.A2(n_746),
.B1(n_747),
.B2(n_741),
.C(n_735),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2008),
.A2(n_1599),
.B(n_1531),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_1989),
.A2(n_1599),
.B(n_1531),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2171),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_1989),
.A2(n_1599),
.B(n_1531),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2018),
.Y(n_2374)
);

AO21x1_ASAP7_75t_L g2375 ( 
.A1(n_2101),
.A2(n_746),
.B(n_741),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_L g2376 ( 
.A1(n_2183),
.A2(n_1465),
.B(n_1437),
.Y(n_2376)
);

OAI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2121),
.A2(n_1333),
.B(n_1312),
.Y(n_2377)
);

AOI21xp5_ASAP7_75t_L g2378 ( 
.A1(n_2196),
.A2(n_1599),
.B(n_1531),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1976),
.B(n_615),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2119),
.B(n_1665),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2196),
.A2(n_1602),
.B(n_1465),
.Y(n_2381)
);

AO21x1_ASAP7_75t_L g2382 ( 
.A1(n_2102),
.A2(n_750),
.B(n_747),
.Y(n_2382)
);

AO31x2_ASAP7_75t_L g2383 ( 
.A1(n_2131),
.A2(n_647),
.A3(n_698),
.B(n_654),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2133),
.A2(n_1437),
.B(n_1230),
.Y(n_2384)
);

OAI21x1_ASAP7_75t_L g2385 ( 
.A1(n_2137),
.A2(n_1230),
.B(n_1436),
.Y(n_2385)
);

OAI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2080),
.A2(n_1333),
.B(n_1681),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_1976),
.B(n_550),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2139),
.A2(n_1230),
.B(n_1441),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2065),
.A2(n_1333),
.B(n_1681),
.Y(n_2389)
);

BUFx12f_ASAP7_75t_L g2390 ( 
.A(n_2069),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2090),
.A2(n_1602),
.B(n_1872),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1985),
.B(n_619),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2012),
.B(n_1665),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2103),
.Y(n_2394)
);

OAI21x1_ASAP7_75t_L g2395 ( 
.A1(n_2141),
.A2(n_1495),
.B(n_1872),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1984),
.B(n_1665),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2077),
.A2(n_1602),
.B1(n_1716),
.B2(n_1665),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2079),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1985),
.B(n_621),
.Y(n_2399)
);

O2A1O1Ixp5_ASAP7_75t_L g2400 ( 
.A1(n_2107),
.A2(n_756),
.B(n_764),
.C(n_750),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2116),
.Y(n_2401)
);

AO32x2_ASAP7_75t_L g2402 ( 
.A1(n_2073),
.A2(n_2149),
.A3(n_1981),
.B1(n_2030),
.B2(n_2066),
.Y(n_2402)
);

OAI21x1_ASAP7_75t_L g2403 ( 
.A1(n_2154),
.A2(n_1872),
.B(n_1027),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2031),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2147),
.Y(n_2405)
);

AOI21x1_ASAP7_75t_SL g2406 ( 
.A1(n_2103),
.A2(n_1872),
.B(n_1744),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2119),
.B(n_1716),
.Y(n_2407)
);

OAI21x1_ASAP7_75t_L g2408 ( 
.A1(n_2163),
.A2(n_1027),
.B(n_1012),
.Y(n_2408)
);

A2O1A1Ixp33_ASAP7_75t_L g2409 ( 
.A1(n_2041),
.A2(n_702),
.B(n_764),
.C(n_756),
.Y(n_2409)
);

OAI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2092),
.A2(n_2175),
.B(n_2041),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2077),
.B(n_2115),
.Y(n_2411)
);

AND2x6_ASAP7_75t_L g2412 ( 
.A(n_2201),
.B(n_1602),
.Y(n_2412)
);

AOI21xp33_ASAP7_75t_L g2413 ( 
.A1(n_2151),
.A2(n_2088),
.B(n_2086),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2165),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2000),
.B(n_622),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2054),
.Y(n_2416)
);

AOI21x1_ASAP7_75t_L g2417 ( 
.A1(n_2098),
.A2(n_887),
.B(n_885),
.Y(n_2417)
);

A2O1A1Ixp33_ASAP7_75t_L g2418 ( 
.A1(n_2085),
.A2(n_1981),
.B(n_2147),
.C(n_2172),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2093),
.B(n_629),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_2173),
.Y(n_2420)
);

A2O1A1Ixp33_ASAP7_75t_L g2421 ( 
.A1(n_2085),
.A2(n_702),
.B(n_590),
.C(n_634),
.Y(n_2421)
);

AO21x1_ASAP7_75t_L g2422 ( 
.A1(n_2174),
.A2(n_887),
.B(n_885),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2184),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2016),
.B(n_2040),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2026),
.B(n_632),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2192),
.Y(n_2426)
);

A2O1A1Ixp33_ASAP7_75t_L g2427 ( 
.A1(n_2197),
.A2(n_590),
.B(n_637),
.C(n_636),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2004),
.Y(n_2428)
);

OAI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2122),
.A2(n_1704),
.B(n_1681),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2129),
.A2(n_1734),
.B1(n_1747),
.B2(n_1716),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2011),
.B(n_675),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2057),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2173),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2011),
.B(n_675),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2026),
.B(n_638),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_1978),
.B(n_641),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2198),
.A2(n_1012),
.B(n_793),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2068),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2010),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2076),
.B(n_2078),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2082),
.B(n_2096),
.Y(n_2441)
);

AOI21xp33_ASAP7_75t_L g2442 ( 
.A1(n_2086),
.A2(n_1747),
.B(n_1734),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2097),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2108),
.B(n_1716),
.Y(n_2444)
);

OAI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2122),
.A2(n_1704),
.B(n_1681),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2090),
.A2(n_2201),
.B(n_2138),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2117),
.B(n_642),
.Y(n_2447)
);

OAI21x1_ASAP7_75t_L g2448 ( 
.A1(n_2125),
.A2(n_892),
.B(n_890),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2134),
.A2(n_892),
.B(n_890),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2091),
.Y(n_2450)
);

OAI21x1_ASAP7_75t_L g2451 ( 
.A1(n_2161),
.A2(n_793),
.B(n_792),
.Y(n_2451)
);

OAI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2189),
.A2(n_1704),
.B(n_1414),
.Y(n_2452)
);

AOI21x1_ASAP7_75t_L g2453 ( 
.A1(n_2166),
.A2(n_896),
.B(n_893),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2155),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2090),
.A2(n_1349),
.B(n_1287),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2200),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2203),
.B(n_643),
.Y(n_2457)
);

A2O1A1Ixp33_ASAP7_75t_L g2458 ( 
.A1(n_2191),
.A2(n_590),
.B(n_648),
.C(n_645),
.Y(n_2458)
);

O2A1O1Ixp33_ASAP7_75t_L g2459 ( 
.A1(n_2108),
.A2(n_896),
.B(n_897),
.C(n_893),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2155),
.B(n_1734),
.Y(n_2460)
);

AOI21x1_ASAP7_75t_L g2461 ( 
.A1(n_2138),
.A2(n_2088),
.B(n_2086),
.Y(n_2461)
);

INVx4_ASAP7_75t_L g2462 ( 
.A(n_2011),
.Y(n_2462)
);

OAI21x1_ASAP7_75t_L g2463 ( 
.A1(n_2159),
.A2(n_899),
.B(n_897),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_SL g2464 ( 
.A1(n_2073),
.A2(n_900),
.B(n_899),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_1996),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2201),
.A2(n_2138),
.B(n_2191),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2088),
.A2(n_1747),
.B1(n_1734),
.B2(n_650),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2201),
.A2(n_1349),
.B(n_1287),
.Y(n_2468)
);

OAI21x1_ASAP7_75t_L g2469 ( 
.A1(n_2159),
.A2(n_795),
.B(n_792),
.Y(n_2469)
);

AOI221xp5_ASAP7_75t_L g2470 ( 
.A1(n_2020),
.A2(n_653),
.B1(n_655),
.B2(n_651),
.C(n_649),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_1996),
.Y(n_2471)
);

A2O1A1Ixp33_ASAP7_75t_L g2472 ( 
.A1(n_2188),
.A2(n_661),
.B(n_662),
.C(n_657),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2465),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2223),
.Y(n_2474)
);

AND2x4_ASAP7_75t_L g2475 ( 
.A(n_2219),
.B(n_2173),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2223),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2218),
.A2(n_2173),
.B(n_2159),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2256),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2297),
.B(n_2411),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2232),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_SL g2481 ( 
.A1(n_2225),
.A2(n_2135),
.B1(n_2020),
.B2(n_675),
.Y(n_2481)
);

INVx2_ASAP7_75t_SL g2482 ( 
.A(n_2287),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2244),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2232),
.Y(n_2484)
);

INVxp33_ASAP7_75t_L g2485 ( 
.A(n_2424),
.Y(n_2485)
);

OR2x6_ASAP7_75t_L g2486 ( 
.A(n_2278),
.B(n_2023),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2248),
.Y(n_2487)
);

AND2x4_ASAP7_75t_L g2488 ( 
.A(n_2219),
.B(n_2043),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2353),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2248),
.Y(n_2490)
);

INVxp67_ASAP7_75t_L g2491 ( 
.A(n_2359),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_2268),
.Y(n_2492)
);

INVx3_ASAP7_75t_SL g2493 ( 
.A(n_2256),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2242),
.A2(n_2159),
.B(n_2135),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2244),
.Y(n_2495)
);

BUFx4_ASAP7_75t_SL g2496 ( 
.A(n_2268),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2303),
.B(n_2144),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2281),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2287),
.Y(n_2499)
);

INVx5_ASAP7_75t_L g2500 ( 
.A(n_2278),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2296),
.B(n_2217),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2359),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2281),
.Y(n_2503)
);

CKINVDCx20_ASAP7_75t_R g2504 ( 
.A(n_2309),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2215),
.Y(n_2505)
);

AOI22xp5_ASAP7_75t_L g2506 ( 
.A1(n_2364),
.A2(n_2037),
.B1(n_2087),
.B2(n_2084),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2454),
.B(n_2156),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2220),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2346),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2276),
.A2(n_2037),
.B1(n_667),
.B2(n_668),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2222),
.B(n_2144),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2465),
.Y(n_2512)
);

NAND2xp33_ASAP7_75t_SL g2513 ( 
.A(n_2224),
.B(n_2056),
.Y(n_2513)
);

NOR2x1_ASAP7_75t_SL g2514 ( 
.A(n_2278),
.B(n_1996),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2319),
.B(n_2144),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2231),
.B(n_2226),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2439),
.B(n_666),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2234),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_L g2519 ( 
.A1(n_2235),
.A2(n_705),
.B1(n_673),
.B2(n_677),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2248),
.Y(n_2520)
);

INVx2_ASAP7_75t_SL g2521 ( 
.A(n_2398),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2365),
.B(n_670),
.Y(n_2522)
);

AO21x1_ASAP7_75t_L g2523 ( 
.A1(n_2235),
.A2(n_902),
.B(n_900),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_2364),
.A2(n_705),
.B1(n_686),
.B2(n_687),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2355),
.A2(n_2308),
.B1(n_2310),
.B2(n_2276),
.Y(n_2525)
);

AOI221xp5_ASAP7_75t_L g2526 ( 
.A1(n_2290),
.A2(n_689),
.B1(n_690),
.B2(n_688),
.C(n_683),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2398),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2299),
.B(n_2144),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2454),
.B(n_2308),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2266),
.Y(n_2530)
);

INVx3_ASAP7_75t_SL g2531 ( 
.A(n_2428),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2390),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2390),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2267),
.Y(n_2534)
);

OAI22xp5_ASAP7_75t_L g2535 ( 
.A1(n_2206),
.A2(n_694),
.B1(n_700),
.B2(n_692),
.Y(n_2535)
);

AOI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2291),
.A2(n_716),
.B1(n_719),
.B2(n_718),
.Y(n_2536)
);

INVx8_ASAP7_75t_L g2537 ( 
.A(n_2412),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2461),
.B(n_1996),
.Y(n_2538)
);

INVx2_ASAP7_75t_SL g2539 ( 
.A(n_2351),
.Y(n_2539)
);

CKINVDCx6p67_ASAP7_75t_R g2540 ( 
.A(n_2248),
.Y(n_2540)
);

OR2x6_ASAP7_75t_L g2541 ( 
.A(n_2237),
.B(n_2002),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2346),
.Y(n_2542)
);

BUFx2_ASAP7_75t_SL g2543 ( 
.A(n_2280),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2262),
.Y(n_2544)
);

BUFx12f_ASAP7_75t_L g2545 ( 
.A(n_2450),
.Y(n_2545)
);

CKINVDCx14_ASAP7_75t_R g2546 ( 
.A(n_2387),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2291),
.A2(n_722),
.B1(n_733),
.B2(n_727),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2307),
.B(n_2144),
.Y(n_2548)
);

INVx1_ASAP7_75t_SL g2549 ( 
.A(n_2340),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2262),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2230),
.B(n_2002),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2213),
.A2(n_2310),
.B1(n_2409),
.B2(n_2221),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_L g2553 ( 
.A(n_2263),
.Y(n_2553)
);

OAI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2409),
.A2(n_736),
.B1(n_737),
.B2(n_734),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2302),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2313),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2280),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2251),
.A2(n_2159),
.B(n_2194),
.Y(n_2558)
);

INVx3_ASAP7_75t_L g2559 ( 
.A(n_2465),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2300),
.A2(n_740),
.B1(n_757),
.B2(n_739),
.Y(n_2560)
);

HAxp5_ASAP7_75t_L g2561 ( 
.A(n_2470),
.B(n_759),
.CON(n_2561),
.SN(n_2561)
);

AOI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2292),
.A2(n_2159),
.B(n_2194),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2374),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2325),
.B(n_2335),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2300),
.A2(n_762),
.B1(n_765),
.B2(n_761),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2273),
.A2(n_2089),
.B(n_2002),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2393),
.Y(n_2567)
);

BUFx4f_ASAP7_75t_L g2568 ( 
.A(n_2263),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2329),
.Y(n_2569)
);

BUFx2_ASAP7_75t_L g2570 ( 
.A(n_2311),
.Y(n_2570)
);

INVx5_ASAP7_75t_L g2571 ( 
.A(n_2412),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_2263),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2374),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2259),
.A2(n_2089),
.B(n_2002),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2450),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2460),
.B(n_2111),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_2410),
.B(n_2056),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2336),
.B(n_2089),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_2450),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2460),
.B(n_2089),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2358),
.Y(n_2581)
);

CKINVDCx11_ASAP7_75t_R g2582 ( 
.A(n_2450),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2311),
.B(n_2111),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2404),
.Y(n_2584)
);

BUFx3_ASAP7_75t_L g2585 ( 
.A(n_2263),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2312),
.B(n_2095),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_SL g2587 ( 
.A1(n_2367),
.A2(n_766),
.B1(n_2104),
.B2(n_2095),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2286),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2431),
.A2(n_1744),
.B1(n_1648),
.B2(n_1414),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2404),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2340),
.B(n_2095),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2420),
.Y(n_2592)
);

OAI21x1_ASAP7_75t_L g2593 ( 
.A1(n_2209),
.A2(n_2212),
.B(n_2403),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2401),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2465),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2238),
.B(n_2095),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2383),
.B(n_2274),
.Y(n_2597)
);

INVx3_ASAP7_75t_L g2598 ( 
.A(n_2286),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2383),
.B(n_2104),
.Y(n_2599)
);

NOR2xp33_ASAP7_75t_R g2600 ( 
.A(n_2339),
.B(n_2104),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_2340),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2434),
.A2(n_1744),
.B1(n_1648),
.B2(n_1414),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2413),
.A2(n_705),
.B1(n_1414),
.B2(n_2104),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2416),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2393),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_2237),
.B(n_2111),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2383),
.B(n_2111),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2420),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2383),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2414),
.Y(n_2610)
);

NAND3xp33_ASAP7_75t_L g2611 ( 
.A(n_2369),
.B(n_796),
.C(n_795),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2257),
.B(n_1704),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2423),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2230),
.A2(n_705),
.B1(n_1414),
.B2(n_1704),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2254),
.A2(n_1648),
.B(n_1747),
.Y(n_2615)
);

CKINVDCx6p67_ASAP7_75t_R g2616 ( 
.A(n_2286),
.Y(n_2616)
);

OAI21xp33_ASAP7_75t_L g2617 ( 
.A1(n_2332),
.A2(n_798),
.B(n_796),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2286),
.Y(n_2618)
);

INVx1_ASAP7_75t_SL g2619 ( 
.A(n_2433),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2321),
.Y(n_2620)
);

OAI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2368),
.A2(n_1000),
.B1(n_903),
.B2(n_905),
.Y(n_2621)
);

INVx3_ASAP7_75t_SL g2622 ( 
.A(n_2380),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_2321),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2396),
.Y(n_2624)
);

INVx2_ASAP7_75t_SL g2625 ( 
.A(n_2321),
.Y(n_2625)
);

NAND2x2_ASAP7_75t_L g2626 ( 
.A(n_2425),
.B(n_1),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2294),
.B(n_2433),
.Y(n_2627)
);

BUFx3_ASAP7_75t_L g2628 ( 
.A(n_2321),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2416),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2405),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2294),
.B(n_348),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2240),
.A2(n_2332),
.B1(n_2304),
.B2(n_2421),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2471),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2396),
.Y(n_2634)
);

OR2x6_ASAP7_75t_L g2635 ( 
.A(n_2348),
.B(n_1000),
.Y(n_2635)
);

AOI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2322),
.A2(n_1349),
.B(n_1287),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2301),
.B(n_1000),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2426),
.Y(n_2638)
);

AOI222xp33_ASAP7_75t_L g2639 ( 
.A1(n_2360),
.A2(n_801),
.B1(n_799),
.B2(n_806),
.C1(n_800),
.C2(n_798),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2418),
.B(n_1000),
.Y(n_2640)
);

O2A1O1Ixp33_ASAP7_75t_L g2641 ( 
.A1(n_2421),
.A2(n_903),
.B(n_905),
.C(n_902),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2432),
.Y(n_2642)
);

BUFx12f_ASAP7_75t_L g2643 ( 
.A(n_2405),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2205),
.B(n_2229),
.Y(n_2644)
);

CKINVDCx6p67_ASAP7_75t_R g2645 ( 
.A(n_2405),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2233),
.B(n_908),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2443),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2405),
.Y(n_2648)
);

INVx2_ASAP7_75t_SL g2649 ( 
.A(n_2317),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2233),
.B(n_908),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2261),
.A2(n_1349),
.B(n_1287),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2418),
.B(n_1000),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2228),
.Y(n_2653)
);

CKINVDCx20_ASAP7_75t_R g2654 ( 
.A(n_2379),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2304),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2435),
.A2(n_1414),
.B1(n_705),
.B2(n_1469),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2258),
.A2(n_1349),
.B(n_1287),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2228),
.Y(n_2658)
);

INVx4_ASAP7_75t_L g2659 ( 
.A(n_2282),
.Y(n_2659)
);

BUFx3_ASAP7_75t_L g2660 ( 
.A(n_2444),
.Y(n_2660)
);

NAND3xp33_ASAP7_75t_L g2661 ( 
.A(n_2458),
.B(n_800),
.C(n_799),
.Y(n_2661)
);

NAND2x1p5_ASAP7_75t_L g2662 ( 
.A(n_2352),
.B(n_1142),
.Y(n_2662)
);

BUFx2_ASAP7_75t_L g2663 ( 
.A(n_2216),
.Y(n_2663)
);

OR2x6_ASAP7_75t_SL g2664 ( 
.A(n_2366),
.B(n_914),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2282),
.Y(n_2665)
);

CKINVDCx20_ASAP7_75t_R g2666 ( 
.A(n_2392),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_2375),
.A2(n_705),
.B1(n_1414),
.B2(n_1469),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2316),
.A2(n_2324),
.B1(n_2245),
.B2(n_2241),
.Y(n_2668)
);

OR2x6_ASAP7_75t_L g2669 ( 
.A(n_2288),
.B(n_1006),
.Y(n_2669)
);

BUFx3_ASAP7_75t_L g2670 ( 
.A(n_2444),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2432),
.Y(n_2671)
);

INVx3_ASAP7_75t_SL g2672 ( 
.A(n_2380),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2330),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2233),
.B(n_915),
.Y(n_2674)
);

OAI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2462),
.A2(n_915),
.B1(n_806),
.B2(n_809),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2330),
.Y(n_2676)
);

INVx4_ASAP7_75t_L g2677 ( 
.A(n_2412),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2415),
.B(n_2399),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2462),
.B(n_354),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2258),
.A2(n_1349),
.B(n_1287),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2361),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2438),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2341),
.B(n_705),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2438),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2456),
.Y(n_2685)
);

O2A1O1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2458),
.A2(n_809),
.B(n_812),
.C(n_801),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2394),
.B(n_356),
.Y(n_2687)
);

OR2x6_ASAP7_75t_L g2688 ( 
.A(n_2243),
.B(n_1006),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2394),
.B(n_705),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2361),
.B(n_357),
.Y(n_2690)
);

INVx2_ASAP7_75t_SL g2691 ( 
.A(n_2380),
.Y(n_2691)
);

OAI21x1_ASAP7_75t_L g2692 ( 
.A1(n_2209),
.A2(n_936),
.B(n_813),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2407),
.B(n_2337),
.Y(n_2693)
);

AOI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2289),
.A2(n_1415),
.B(n_1182),
.Y(n_2694)
);

CKINVDCx20_ASAP7_75t_R g2695 ( 
.A(n_2419),
.Y(n_2695)
);

CKINVDCx20_ASAP7_75t_R g2696 ( 
.A(n_2436),
.Y(n_2696)
);

INVx5_ASAP7_75t_L g2697 ( 
.A(n_2412),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2372),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2372),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2233),
.B(n_2),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2407),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_2382),
.A2(n_1469),
.B1(n_813),
.B2(n_814),
.Y(n_2702)
);

BUFx2_ASAP7_75t_L g2703 ( 
.A(n_2216),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2283),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2216),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2241),
.B(n_4),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2245),
.B(n_5),
.Y(n_2707)
);

OR2x6_ASAP7_75t_L g2708 ( 
.A(n_2466),
.B(n_1006),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2407),
.B(n_359),
.Y(n_2709)
);

OAI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2472),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2710)
);

BUFx8_ASAP7_75t_L g2711 ( 
.A(n_2402),
.Y(n_2711)
);

NAND2x1_ASAP7_75t_L g2712 ( 
.A(n_2216),
.B(n_1142),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2446),
.B(n_361),
.Y(n_2713)
);

HB1xp67_ASAP7_75t_L g2714 ( 
.A(n_2456),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2330),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2208),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2330),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_2216),
.B(n_364),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2472),
.B(n_365),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2447),
.B(n_812),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2283),
.Y(n_2721)
);

AND3x1_ASAP7_75t_SL g2722 ( 
.A(n_2211),
.B(n_7),
.C(n_8),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2430),
.Y(n_2723)
);

OAI21xp33_ASAP7_75t_L g2724 ( 
.A1(n_2427),
.A2(n_815),
.B(n_814),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2283),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2290),
.B(n_1006),
.Y(n_2726)
);

BUFx2_ASAP7_75t_L g2727 ( 
.A(n_2412),
.Y(n_2727)
);

NAND2xp33_ASAP7_75t_SL g2728 ( 
.A(n_2397),
.B(n_9),
.Y(n_2728)
);

NAND2x1_ASAP7_75t_L g2729 ( 
.A(n_2344),
.B(n_1182),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2457),
.B(n_366),
.Y(n_2730)
);

INVx1_ASAP7_75t_SL g2731 ( 
.A(n_2207),
.Y(n_2731)
);

NAND3xp33_ASAP7_75t_L g2732 ( 
.A(n_2427),
.B(n_816),
.C(n_815),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2440),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2207),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2508),
.Y(n_2735)
);

OAI21x1_ASAP7_75t_L g2736 ( 
.A1(n_2694),
.A2(n_2227),
.B(n_2306),
.Y(n_2736)
);

AO21x2_ASAP7_75t_L g2737 ( 
.A1(n_2726),
.A2(n_2318),
.B(n_2305),
.Y(n_2737)
);

OAI21x1_ASAP7_75t_L g2738 ( 
.A1(n_2694),
.A2(n_2227),
.B(n_2269),
.Y(n_2738)
);

INVx3_ASAP7_75t_L g2739 ( 
.A(n_2599),
.Y(n_2739)
);

OAI21x1_ASAP7_75t_SL g2740 ( 
.A1(n_2514),
.A2(n_2247),
.B(n_2349),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2502),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2480),
.Y(n_2742)
);

OA21x2_ASAP7_75t_L g2743 ( 
.A1(n_2489),
.A2(n_2295),
.B(n_2338),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2610),
.Y(n_2744)
);

NAND3xp33_ASAP7_75t_L g2745 ( 
.A(n_2526),
.B(n_2400),
.C(n_2326),
.Y(n_2745)
);

OAI21x1_ASAP7_75t_SL g2746 ( 
.A1(n_2523),
.A2(n_2260),
.B(n_2422),
.Y(n_2746)
);

OAI21x1_ASAP7_75t_L g2747 ( 
.A1(n_2593),
.A2(n_2558),
.B(n_2692),
.Y(n_2747)
);

AOI22x1_ASAP7_75t_L g2748 ( 
.A1(n_2587),
.A2(n_2214),
.B1(n_2464),
.B2(n_2389),
.Y(n_2748)
);

AO21x2_ASAP7_75t_L g2749 ( 
.A1(n_2646),
.A2(n_2318),
.B(n_2429),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2526),
.B(n_2253),
.Y(n_2750)
);

OAI21x1_ASAP7_75t_L g2751 ( 
.A1(n_2558),
.A2(n_2269),
.B(n_2264),
.Y(n_2751)
);

AO222x2_ASAP7_75t_L g2752 ( 
.A1(n_2664),
.A2(n_13),
.B1(n_15),
.B2(n_9),
.C1(n_12),
.C2(n_14),
.Y(n_2752)
);

OAI21x1_ASAP7_75t_L g2753 ( 
.A1(n_2651),
.A2(n_2264),
.B(n_2384),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2660),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2651),
.A2(n_2384),
.B(n_2239),
.Y(n_2755)
);

OAI21x1_ASAP7_75t_L g2756 ( 
.A1(n_2562),
.A2(n_2338),
.B(n_2249),
.Y(n_2756)
);

AND2x4_ASAP7_75t_L g2757 ( 
.A(n_2500),
.B(n_2283),
.Y(n_2757)
);

OAI21x1_ASAP7_75t_L g2758 ( 
.A1(n_2562),
.A2(n_2295),
.B(n_2250),
.Y(n_2758)
);

OAI21x1_ASAP7_75t_L g2759 ( 
.A1(n_2615),
.A2(n_2320),
.B(n_2270),
.Y(n_2759)
);

OAI21x1_ASAP7_75t_L g2760 ( 
.A1(n_2615),
.A2(n_2320),
.B(n_2270),
.Y(n_2760)
);

BUFx12f_ASAP7_75t_L g2761 ( 
.A(n_2544),
.Y(n_2761)
);

OAI21x1_ASAP7_75t_L g2762 ( 
.A1(n_2636),
.A2(n_2395),
.B(n_2275),
.Y(n_2762)
);

OR2x2_ASAP7_75t_L g2763 ( 
.A(n_2597),
.B(n_2236),
.Y(n_2763)
);

AOI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2481),
.A2(n_2252),
.B1(n_2327),
.B2(n_2255),
.Y(n_2764)
);

OAI21x1_ASAP7_75t_L g2765 ( 
.A1(n_2636),
.A2(n_2463),
.B(n_2271),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2484),
.Y(n_2766)
);

OAI222xp33_ASAP7_75t_L g2767 ( 
.A1(n_2481),
.A2(n_2214),
.B1(n_2285),
.B2(n_2441),
.C1(n_2467),
.C2(n_2333),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2536),
.A2(n_2386),
.B1(n_2377),
.B2(n_2345),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2494),
.A2(n_2477),
.B(n_2644),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_SL g2770 ( 
.A1(n_2706),
.A2(n_2445),
.B(n_2453),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2479),
.B(n_2529),
.Y(n_2771)
);

OAI21x1_ASAP7_75t_L g2772 ( 
.A1(n_2477),
.A2(n_2463),
.B(n_2362),
.Y(n_2772)
);

OAI21x1_ASAP7_75t_L g2773 ( 
.A1(n_2494),
.A2(n_2362),
.B(n_2448),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2525),
.A2(n_2333),
.B1(n_2373),
.B2(n_2371),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2501),
.B(n_2442),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_L g2776 ( 
.A(n_2501),
.B(n_2272),
.Y(n_2776)
);

OAI21x1_ASAP7_75t_L g2777 ( 
.A1(n_2566),
.A2(n_2680),
.B(n_2657),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2644),
.A2(n_2370),
.B(n_2452),
.Y(n_2778)
);

AO21x2_ASAP7_75t_L g2779 ( 
.A1(n_2646),
.A2(n_2391),
.B(n_2363),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_L g2780 ( 
.A1(n_2566),
.A2(n_2449),
.B(n_2448),
.Y(n_2780)
);

OAI21x1_ASAP7_75t_L g2781 ( 
.A1(n_2657),
.A2(n_2449),
.B(n_2265),
.Y(n_2781)
);

O2A1O1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_2710),
.A2(n_2655),
.B(n_2707),
.C(n_2706),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_L g2783 ( 
.A1(n_2710),
.A2(n_2343),
.B1(n_2357),
.B2(n_2211),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2668),
.B(n_2400),
.Y(n_2784)
);

OAI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2680),
.A2(n_2265),
.B(n_2385),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2607),
.Y(n_2786)
);

OAI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2519),
.A2(n_2459),
.B(n_2378),
.Y(n_2787)
);

OAI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2547),
.A2(n_2381),
.B(n_2437),
.Y(n_2788)
);

OAI21x1_ASAP7_75t_L g2789 ( 
.A1(n_2574),
.A2(n_2388),
.B(n_2408),
.Y(n_2789)
);

CKINVDCx20_ASAP7_75t_R g2790 ( 
.A(n_2504),
.Y(n_2790)
);

OAI21x1_ASAP7_75t_SL g2791 ( 
.A1(n_2707),
.A2(n_2417),
.B(n_2328),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2505),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2491),
.Y(n_2793)
);

CKINVDCx16_ASAP7_75t_R g2794 ( 
.A(n_2695),
.Y(n_2794)
);

AND2x4_ASAP7_75t_L g2795 ( 
.A(n_2500),
.B(n_2246),
.Y(n_2795)
);

OA21x2_ASAP7_75t_L g2796 ( 
.A1(n_2609),
.A2(n_2354),
.B(n_2350),
.Y(n_2796)
);

AO21x2_ASAP7_75t_L g2797 ( 
.A1(n_2650),
.A2(n_2376),
.B(n_2356),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2552),
.A2(n_2678),
.B1(n_2577),
.B2(n_2719),
.Y(n_2798)
);

OAI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2655),
.A2(n_2451),
.B(n_2279),
.Y(n_2799)
);

OAI21x1_ASAP7_75t_L g2800 ( 
.A1(n_2574),
.A2(n_2406),
.B(n_2323),
.Y(n_2800)
);

INVx3_ASAP7_75t_L g2801 ( 
.A(n_2538),
.Y(n_2801)
);

AO31x2_ASAP7_75t_L g2802 ( 
.A1(n_2673),
.A2(n_2455),
.A3(n_2298),
.B(n_2314),
.Y(n_2802)
);

OAI21x1_ASAP7_75t_L g2803 ( 
.A1(n_2676),
.A2(n_2406),
.B(n_2469),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2613),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2518),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2530),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2534),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2582),
.Y(n_2808)
);

AO21x2_ASAP7_75t_L g2809 ( 
.A1(n_2650),
.A2(n_2284),
.B(n_2277),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2555),
.Y(n_2810)
);

A2O1A1Ixp33_ASAP7_75t_L g2811 ( 
.A1(n_2728),
.A2(n_2402),
.B(n_2468),
.C(n_2293),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2556),
.Y(n_2812)
);

AO31x2_ASAP7_75t_L g2813 ( 
.A1(n_2715),
.A2(n_2236),
.A3(n_2246),
.B(n_2210),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2552),
.A2(n_2347),
.B1(n_816),
.B2(n_2334),
.Y(n_2814)
);

AND2x4_ASAP7_75t_L g2815 ( 
.A(n_2500),
.B(n_2246),
.Y(n_2815)
);

INVx2_ASAP7_75t_SL g2816 ( 
.A(n_2500),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2638),
.Y(n_2817)
);

A2O1A1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_2641),
.A2(n_2402),
.B(n_2315),
.C(n_2342),
.Y(n_2818)
);

HB1xp67_ASAP7_75t_L g2819 ( 
.A(n_2491),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2658),
.Y(n_2820)
);

OA21x2_ASAP7_75t_L g2821 ( 
.A1(n_2700),
.A2(n_2331),
.B(n_2236),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2668),
.B(n_13),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2714),
.Y(n_2823)
);

INVxp33_ASAP7_75t_SL g2824 ( 
.A(n_2496),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_SL g2825 ( 
.A(n_2478),
.B(n_2402),
.Y(n_2825)
);

HB1xp67_ASAP7_75t_L g2826 ( 
.A(n_2633),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_L g2827 ( 
.A1(n_2717),
.A2(n_2347),
.B(n_2236),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2549),
.B(n_2246),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2569),
.Y(n_2829)
);

NAND2x1p5_ASAP7_75t_L g2830 ( 
.A(n_2571),
.B(n_2347),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2499),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2535),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2516),
.B(n_2210),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2711),
.A2(n_2210),
.B1(n_20),
.B2(n_18),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2670),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2516),
.B(n_2210),
.Y(n_2836)
);

NAND2x1p5_ASAP7_75t_L g2837 ( 
.A(n_2571),
.B(n_1006),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2581),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2594),
.Y(n_2839)
);

OAI21x1_ASAP7_75t_L g2840 ( 
.A1(n_2662),
.A2(n_2725),
.B(n_2721),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2647),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2524),
.A2(n_1469),
.B(n_936),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2700),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2685),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2649),
.B(n_18),
.Y(n_2845)
);

INVx1_ASAP7_75t_SL g2846 ( 
.A(n_2531),
.Y(n_2846)
);

OR2x6_ASAP7_75t_L g2847 ( 
.A(n_2669),
.B(n_1007),
.Y(n_2847)
);

AOI21xp33_ASAP7_75t_SL g2848 ( 
.A1(n_2493),
.A2(n_19),
.B(n_20),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2685),
.Y(n_2849)
);

AO21x2_ASAP7_75t_L g2850 ( 
.A1(n_2674),
.A2(n_1469),
.B(n_19),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2474),
.Y(n_2851)
);

OAI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2632),
.A2(n_1469),
.B(n_936),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2632),
.A2(n_1469),
.B(n_928),
.Y(n_2853)
);

OAI21x1_ASAP7_75t_L g2854 ( 
.A1(n_2662),
.A2(n_370),
.B(n_369),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2576),
.B(n_2580),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2608),
.Y(n_2856)
);

OA21x2_ASAP7_75t_L g2857 ( 
.A1(n_2674),
.A2(n_21),
.B(n_23),
.Y(n_2857)
);

OAI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2538),
.A2(n_373),
.B(n_372),
.Y(n_2858)
);

BUFx3_ASAP7_75t_L g2859 ( 
.A(n_2527),
.Y(n_2859)
);

OA21x2_ASAP7_75t_L g2860 ( 
.A1(n_2704),
.A2(n_21),
.B(n_23),
.Y(n_2860)
);

OAI21x1_ASAP7_75t_L g2861 ( 
.A1(n_2712),
.A2(n_377),
.B(n_376),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2476),
.Y(n_2862)
);

AO21x2_ASAP7_75t_L g2863 ( 
.A1(n_2640),
.A2(n_25),
.B(n_26),
.Y(n_2863)
);

NOR2x1_ASAP7_75t_SL g2864 ( 
.A(n_2688),
.B(n_2708),
.Y(n_2864)
);

OAI21x1_ASAP7_75t_L g2865 ( 
.A1(n_2515),
.A2(n_390),
.B(n_389),
.Y(n_2865)
);

OAI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2730),
.A2(n_928),
.B(n_394),
.Y(n_2866)
);

OAI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2535),
.A2(n_928),
.B(n_396),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2483),
.Y(n_2868)
);

INVxp67_ASAP7_75t_L g2869 ( 
.A(n_2522),
.Y(n_2869)
);

INVxp67_ASAP7_75t_L g2870 ( 
.A(n_2539),
.Y(n_2870)
);

OA21x2_ASAP7_75t_L g2871 ( 
.A1(n_2704),
.A2(n_25),
.B(n_27),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2495),
.Y(n_2872)
);

OA21x2_ASAP7_75t_L g2873 ( 
.A1(n_2652),
.A2(n_2511),
.B(n_2515),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2498),
.Y(n_2874)
);

OA21x2_ASAP7_75t_L g2875 ( 
.A1(n_2511),
.A2(n_27),
.B(n_28),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2688),
.A2(n_1415),
.B(n_1196),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2564),
.B(n_28),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2503),
.Y(n_2878)
);

BUFx8_ASAP7_75t_L g2879 ( 
.A(n_2643),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2549),
.B(n_392),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2509),
.Y(n_2881)
);

OAI21x1_ASAP7_75t_L g2882 ( 
.A1(n_2528),
.A2(n_401),
.B(n_399),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2550),
.Y(n_2883)
);

OAI22x1_ASAP7_75t_L g2884 ( 
.A1(n_2567),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2884)
);

OAI21x1_ASAP7_75t_L g2885 ( 
.A1(n_2528),
.A2(n_2548),
.B(n_2612),
.Y(n_2885)
);

NAND3xp33_ASAP7_75t_L g2886 ( 
.A(n_2510),
.B(n_1019),
.C(n_1007),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2496),
.Y(n_2887)
);

NOR2x1_ASAP7_75t_SL g2888 ( 
.A(n_2688),
.B(n_1007),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2542),
.Y(n_2889)
);

HB1xp67_ASAP7_75t_L g2890 ( 
.A(n_2578),
.Y(n_2890)
);

BUFx6f_ASAP7_75t_L g2891 ( 
.A(n_2658),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2563),
.Y(n_2892)
);

OAI21x1_ASAP7_75t_L g2893 ( 
.A1(n_2548),
.A2(n_2612),
.B(n_2729),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2693),
.B(n_30),
.Y(n_2894)
);

AO31x2_ASAP7_75t_L g2895 ( 
.A1(n_2677),
.A2(n_928),
.A3(n_1236),
.B(n_1167),
.Y(n_2895)
);

CKINVDCx8_ASAP7_75t_R g2896 ( 
.A(n_2543),
.Y(n_2896)
);

OAI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2497),
.A2(n_404),
.B(n_402),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2601),
.Y(n_2898)
);

OAI21x1_ASAP7_75t_L g2899 ( 
.A1(n_2497),
.A2(n_409),
.B(n_405),
.Y(n_2899)
);

OR2x6_ASAP7_75t_L g2900 ( 
.A(n_2537),
.B(n_1007),
.Y(n_2900)
);

NAND2x1p5_ASAP7_75t_L g2901 ( 
.A(n_2571),
.B(n_1007),
.Y(n_2901)
);

OAI22xp33_ASAP7_75t_L g2902 ( 
.A1(n_2626),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2902)
);

CKINVDCx16_ASAP7_75t_R g2903 ( 
.A(n_2532),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2605),
.B(n_1019),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2637),
.A2(n_1415),
.B(n_1196),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2733),
.B(n_34),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2573),
.Y(n_2907)
);

AOI21xp33_ASAP7_75t_L g2908 ( 
.A1(n_2641),
.A2(n_34),
.B(n_35),
.Y(n_2908)
);

AOI221x1_ASAP7_75t_L g2909 ( 
.A1(n_2554),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.C(n_39),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2571),
.B(n_1019),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2584),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2590),
.Y(n_2912)
);

AOI222xp33_ASAP7_75t_L g2913 ( 
.A1(n_2510),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_2913)
);

OA21x2_ASAP7_75t_L g2914 ( 
.A1(n_2732),
.A2(n_40),
.B(n_41),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2601),
.B(n_42),
.Y(n_2915)
);

AO31x2_ASAP7_75t_L g2916 ( 
.A1(n_2677),
.A2(n_1236),
.A3(n_1167),
.B(n_45),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2604),
.Y(n_2917)
);

AOI22x1_ASAP7_75t_L g2918 ( 
.A1(n_2624),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2629),
.Y(n_2919)
);

AO21x1_ASAP7_75t_L g2920 ( 
.A1(n_2554),
.A2(n_43),
.B(n_46),
.Y(n_2920)
);

OAI21x1_ASAP7_75t_L g2921 ( 
.A1(n_2642),
.A2(n_414),
.B(n_412),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2671),
.Y(n_2922)
);

AOI21x1_ASAP7_75t_L g2923 ( 
.A1(n_2708),
.A2(n_48),
.B(n_49),
.Y(n_2923)
);

OAI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2682),
.A2(n_416),
.B(n_415),
.Y(n_2924)
);

OR2x2_ASAP7_75t_L g2925 ( 
.A(n_2485),
.B(n_2586),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2684),
.Y(n_2926)
);

AO21x2_ASAP7_75t_L g2927 ( 
.A1(n_2600),
.A2(n_2661),
.B(n_2586),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2731),
.Y(n_2928)
);

OAI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2596),
.A2(n_422),
.B(n_418),
.Y(n_2929)
);

AO21x2_ASAP7_75t_L g2930 ( 
.A1(n_2596),
.A2(n_2686),
.B(n_2724),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2689),
.Y(n_2931)
);

AOI221xp5_ASAP7_75t_L g2932 ( 
.A1(n_2560),
.A2(n_52),
.B1(n_49),
.B2(n_51),
.C(n_53),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2686),
.A2(n_1415),
.B(n_1196),
.Y(n_2933)
);

AOI21xp33_ASAP7_75t_SL g2934 ( 
.A1(n_2517),
.A2(n_51),
.B(n_52),
.Y(n_2934)
);

OA21x2_ASAP7_75t_L g2935 ( 
.A1(n_2617),
.A2(n_54),
.B(n_55),
.Y(n_2935)
);

AOI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2654),
.A2(n_2666),
.B1(n_2696),
.B2(n_2713),
.Y(n_2936)
);

OAI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2701),
.A2(n_426),
.B(n_423),
.Y(n_2937)
);

OAI21x1_ASAP7_75t_L g2938 ( 
.A1(n_2701),
.A2(n_431),
.B(n_430),
.Y(n_2938)
);

OAI21x1_ASAP7_75t_L g2939 ( 
.A1(n_2473),
.A2(n_438),
.B(n_435),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2731),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2734),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2734),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2627),
.B(n_439),
.Y(n_2943)
);

HB1xp67_ASAP7_75t_L g2944 ( 
.A(n_2619),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2592),
.Y(n_2945)
);

OAI21x1_ASAP7_75t_L g2946 ( 
.A1(n_2473),
.A2(n_446),
.B(n_442),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2507),
.B(n_54),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2591),
.B(n_56),
.Y(n_2948)
);

AOI221xp5_ASAP7_75t_L g2949 ( 
.A1(n_2560),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.C(n_60),
.Y(n_2949)
);

OAI21x1_ASAP7_75t_L g2950 ( 
.A1(n_2512),
.A2(n_449),
.B(n_447),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2723),
.B(n_60),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2561),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2711),
.Y(n_2953)
);

OAI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2486),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2619),
.Y(n_2955)
);

OAI21x1_ASAP7_75t_L g2956 ( 
.A1(n_2512),
.A2(n_455),
.B(n_454),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2570),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2559),
.A2(n_457),
.B(n_456),
.Y(n_2958)
);

INVx5_ASAP7_75t_L g2959 ( 
.A(n_2900),
.Y(n_2959)
);

INVx4_ASAP7_75t_L g2960 ( 
.A(n_2808),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_SL g2961 ( 
.A(n_2824),
.B(n_2634),
.Y(n_2961)
);

INVx4_ASAP7_75t_SL g2962 ( 
.A(n_2808),
.Y(n_2962)
);

INVxp67_ASAP7_75t_SL g2963 ( 
.A(n_2776),
.Y(n_2963)
);

CKINVDCx20_ASAP7_75t_R g2964 ( 
.A(n_2790),
.Y(n_2964)
);

NAND2xp33_ASAP7_75t_SL g2965 ( 
.A(n_2808),
.B(n_2698),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2896),
.Y(n_2966)
);

INVx4_ASAP7_75t_L g2967 ( 
.A(n_2808),
.Y(n_2967)
);

HB1xp67_ASAP7_75t_L g2968 ( 
.A(n_2843),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2750),
.A2(n_2713),
.B1(n_2486),
.B2(n_2546),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2890),
.B(n_2482),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2798),
.A2(n_2832),
.B1(n_2834),
.B2(n_2750),
.Y(n_2971)
);

AOI221xp5_ASAP7_75t_L g2972 ( 
.A1(n_2782),
.A2(n_2565),
.B1(n_2621),
.B2(n_2611),
.C(n_2683),
.Y(n_2972)
);

AO31x2_ASAP7_75t_L g2973 ( 
.A1(n_2888),
.A2(n_2727),
.A3(n_2663),
.B(n_2705),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2744),
.Y(n_2974)
);

NAND2xp33_ASAP7_75t_R g2975 ( 
.A(n_2824),
.B(n_2486),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2744),
.Y(n_2976)
);

AOI22xp33_ASAP7_75t_L g2977 ( 
.A1(n_2822),
.A2(n_2631),
.B1(n_2718),
.B2(n_2475),
.Y(n_2977)
);

OR2x2_ASAP7_75t_L g2978 ( 
.A(n_2735),
.B(n_2669),
.Y(n_2978)
);

AOI21xp33_ASAP7_75t_L g2979 ( 
.A1(n_2822),
.A2(n_2708),
.B(n_2720),
.Y(n_2979)
);

BUFx2_ASAP7_75t_L g2980 ( 
.A(n_2826),
.Y(n_2980)
);

AND2x2_ASAP7_75t_SL g2981 ( 
.A(n_2794),
.B(n_2703),
.Y(n_2981)
);

OAI221xp5_ASAP7_75t_L g2982 ( 
.A1(n_2952),
.A2(n_2565),
.B1(n_2506),
.B2(n_2603),
.C(n_2513),
.Y(n_2982)
);

AOI22x1_ASAP7_75t_L g2983 ( 
.A1(n_2913),
.A2(n_2884),
.B1(n_2752),
.B2(n_2867),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2771),
.B(n_2521),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_SL g2985 ( 
.A1(n_2752),
.A2(n_2722),
.B1(n_2537),
.B2(n_2718),
.Y(n_2985)
);

OAI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2832),
.A2(n_2589),
.B1(n_2602),
.B2(n_2697),
.Y(n_2986)
);

NAND2xp33_ASAP7_75t_L g2987 ( 
.A(n_2918),
.B(n_2658),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2804),
.Y(n_2988)
);

INVx4_ASAP7_75t_L g2989 ( 
.A(n_2820),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2846),
.B(n_2533),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2804),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2776),
.B(n_2669),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2920),
.A2(n_2631),
.B1(n_2475),
.B2(n_2627),
.Y(n_2993)
);

OAI22xp33_ASAP7_75t_L g2994 ( 
.A1(n_2909),
.A2(n_2697),
.B1(n_2537),
.B2(n_2672),
.Y(n_2994)
);

OR2x2_ASAP7_75t_L g2995 ( 
.A(n_2925),
.B(n_2763),
.Y(n_2995)
);

OAI211xp5_ASAP7_75t_L g2996 ( 
.A1(n_2934),
.A2(n_2639),
.B(n_2702),
.C(n_2667),
.Y(n_2996)
);

NAND2x1p5_ASAP7_75t_L g2997 ( 
.A(n_2875),
.B(n_2697),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2817),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_L g2999 ( 
.A1(n_2751),
.A2(n_2756),
.B(n_2747),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2761),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2775),
.B(n_2492),
.Y(n_3001)
);

AND2x2_ASAP7_75t_SL g3002 ( 
.A(n_2825),
.B(n_2557),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2896),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2745),
.A2(n_2679),
.B1(n_2709),
.B2(n_2687),
.Y(n_3004)
);

CKINVDCx11_ASAP7_75t_R g3005 ( 
.A(n_2790),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2775),
.B(n_2716),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2817),
.Y(n_3007)
);

AOI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2932),
.A2(n_2679),
.B1(n_2709),
.B2(n_2488),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2833),
.B(n_2635),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2829),
.Y(n_3010)
);

NAND2x1p5_ASAP7_75t_L g3011 ( 
.A(n_2875),
.B(n_2697),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2801),
.B(n_2551),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2829),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_L g3014 ( 
.A1(n_2866),
.A2(n_2687),
.B1(n_2690),
.B2(n_2635),
.Y(n_3014)
);

AND2x4_ASAP7_75t_L g3015 ( 
.A(n_2801),
.B(n_2551),
.Y(n_3015)
);

O2A1O1Ixp33_ASAP7_75t_SL g3016 ( 
.A1(n_2902),
.A2(n_2954),
.B(n_2887),
.C(n_2848),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2855),
.B(n_2622),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2823),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_2883),
.Y(n_3019)
);

AND2x4_ASAP7_75t_L g3020 ( 
.A(n_2801),
.B(n_2635),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2949),
.A2(n_2690),
.B1(n_2681),
.B2(n_2691),
.Y(n_3021)
);

AOI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2784),
.A2(n_2488),
.B1(n_2616),
.B2(n_2540),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2739),
.B(n_2559),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2754),
.B(n_2583),
.Y(n_3024)
);

BUFx2_ASAP7_75t_L g3025 ( 
.A(n_2835),
.Y(n_3025)
);

AND2x4_ASAP7_75t_L g3026 ( 
.A(n_2739),
.B(n_2595),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2841),
.Y(n_3027)
);

OAI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2768),
.A2(n_2606),
.B1(n_2541),
.B2(n_2699),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_SL g3029 ( 
.A1(n_2951),
.A2(n_2568),
.B1(n_2699),
.B2(n_2681),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2841),
.Y(n_3030)
);

BUFx3_ASAP7_75t_L g3031 ( 
.A(n_2761),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2784),
.A2(n_2681),
.B1(n_2639),
.B2(n_2585),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_2951),
.A2(n_2628),
.B1(n_2598),
.B2(n_2620),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2739),
.B(n_2595),
.Y(n_3034)
);

AND2x4_ASAP7_75t_L g3035 ( 
.A(n_2786),
.B(n_2541),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2786),
.B(n_2541),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2792),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2805),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2806),
.Y(n_3039)
);

CKINVDCx16_ASAP7_75t_R g3040 ( 
.A(n_2903),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2954),
.A2(n_2598),
.B1(n_2648),
.B2(n_2620),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_2793),
.Y(n_3042)
);

OAI221xp5_ASAP7_75t_L g3043 ( 
.A1(n_2764),
.A2(n_2656),
.B1(n_2568),
.B2(n_2606),
.C(n_2648),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2786),
.B(n_2606),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2831),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2898),
.B(n_2575),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_SL g3047 ( 
.A1(n_2935),
.A2(n_2490),
.B1(n_2520),
.B2(n_2487),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2856),
.B(n_2623),
.Y(n_3048)
);

AOI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2902),
.A2(n_2748),
.B1(n_2908),
.B2(n_2869),
.Y(n_3049)
);

CKINVDCx14_ASAP7_75t_R g3050 ( 
.A(n_2883),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2769),
.A2(n_2675),
.B(n_2614),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2819),
.B(n_2625),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2886),
.A2(n_2545),
.B1(n_2490),
.B2(n_2520),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2836),
.B(n_2487),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2764),
.A2(n_2645),
.B1(n_2665),
.B2(n_2653),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2787),
.A2(n_2490),
.B1(n_2520),
.B2(n_2487),
.Y(n_3056)
);

NAND2x1p5_ASAP7_75t_L g3057 ( 
.A(n_2875),
.B(n_2659),
.Y(n_3057)
);

INVx3_ASAP7_75t_L g3058 ( 
.A(n_2831),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2807),
.Y(n_3059)
);

AND2x4_ASAP7_75t_L g3060 ( 
.A(n_2928),
.B(n_2579),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2859),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2957),
.B(n_2553),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2774),
.A2(n_2659),
.B1(n_2572),
.B2(n_2588),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2788),
.A2(n_2572),
.B1(n_2588),
.B2(n_2553),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2936),
.B(n_2630),
.Y(n_3065)
);

NOR2x1p5_ASAP7_75t_L g3066 ( 
.A(n_2859),
.B(n_2553),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2810),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2812),
.Y(n_3068)
);

OAI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2935),
.A2(n_2588),
.B1(n_2618),
.B2(n_2572),
.Y(n_3069)
);

AOI221xp5_ASAP7_75t_L g3070 ( 
.A1(n_2767),
.A2(n_69),
.B1(n_65),
.B2(n_67),
.C(n_70),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2945),
.B(n_2618),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2944),
.B(n_2618),
.Y(n_3072)
);

CKINVDCx5p33_ASAP7_75t_R g3073 ( 
.A(n_2879),
.Y(n_3073)
);

OAI221xp5_ASAP7_75t_L g3074 ( 
.A1(n_2783),
.A2(n_2630),
.B1(n_69),
.B2(n_65),
.C(n_67),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2838),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_2879),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2839),
.Y(n_3077)
);

OR2x6_ASAP7_75t_SL g3078 ( 
.A(n_2953),
.B(n_2630),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_2940),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2741),
.Y(n_3080)
);

AO21x1_ASAP7_75t_L g3081 ( 
.A1(n_2904),
.A2(n_70),
.B(n_71),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2953),
.B(n_72),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_2783),
.A2(n_1025),
.B1(n_1040),
.B2(n_1019),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_2880),
.A2(n_2931),
.B1(n_2770),
.B2(n_2873),
.Y(n_3084)
);

OR2x2_ASAP7_75t_L g3085 ( 
.A(n_2885),
.B(n_2873),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2820),
.Y(n_3086)
);

CKINVDCx20_ASAP7_75t_R g3087 ( 
.A(n_2879),
.Y(n_3087)
);

CKINVDCx20_ASAP7_75t_R g3088 ( 
.A(n_2887),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2870),
.B(n_73),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2880),
.A2(n_1025),
.B1(n_1040),
.B2(n_1019),
.Y(n_3090)
);

AOI221xp5_ASAP7_75t_L g3091 ( 
.A1(n_2877),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.C(n_78),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2742),
.Y(n_3092)
);

OAI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2904),
.A2(n_80),
.B1(n_75),
.B2(n_79),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2885),
.B(n_79),
.Y(n_3094)
);

OAI221xp5_ASAP7_75t_L g3095 ( 
.A1(n_2814),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.C(n_85),
.Y(n_3095)
);

OAI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_2935),
.A2(n_2914),
.B1(n_2852),
.B2(n_2871),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2766),
.Y(n_3097)
);

NAND2xp33_ASAP7_75t_SL g3098 ( 
.A(n_2880),
.B(n_82),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_2873),
.B(n_83),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_2941),
.B(n_2942),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_SL g3101 ( 
.A(n_2943),
.B(n_1025),
.Y(n_3101)
);

BUFx8_ASAP7_75t_SL g3102 ( 
.A(n_2820),
.Y(n_3102)
);

BUFx8_ASAP7_75t_SL g3103 ( 
.A(n_2820),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_SL g3104 ( 
.A1(n_2811),
.A2(n_1040),
.B(n_1025),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2955),
.B(n_84),
.Y(n_3105)
);

NAND2xp33_ASAP7_75t_SL g3106 ( 
.A(n_2891),
.B(n_85),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_2891),
.Y(n_3107)
);

INVx3_ASAP7_75t_L g3108 ( 
.A(n_2891),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_2891),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2933),
.A2(n_1415),
.B(n_1196),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2844),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_2849),
.B(n_87),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_2900),
.Y(n_3113)
);

OAI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2914),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_SL g3115 ( 
.A(n_2943),
.B(n_1025),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_2828),
.B(n_88),
.Y(n_3116)
);

NAND2x1p5_ASAP7_75t_L g3117 ( 
.A(n_2857),
.B(n_1040),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_L g3118 ( 
.A(n_2943),
.Y(n_3118)
);

OR2x2_ASAP7_75t_L g3119 ( 
.A(n_2828),
.B(n_90),
.Y(n_3119)
);

AOI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_2930),
.A2(n_1040),
.B1(n_1196),
.B2(n_1182),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2862),
.B(n_91),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2814),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2931),
.B(n_95),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2862),
.Y(n_3124)
);

CKINVDCx11_ASAP7_75t_R g3125 ( 
.A(n_2900),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2874),
.Y(n_3126)
);

HB1xp67_ASAP7_75t_L g3127 ( 
.A(n_2821),
.Y(n_3127)
);

OR2x2_ASAP7_75t_L g3128 ( 
.A(n_2828),
.B(n_95),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2930),
.A2(n_99),
.B1(n_96),
.B2(n_97),
.Y(n_3129)
);

NAND2xp33_ASAP7_75t_SL g3130 ( 
.A(n_2845),
.B(n_96),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2874),
.B(n_97),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2893),
.B(n_100),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_2816),
.B(n_101),
.Y(n_3133)
);

OAI221xp5_ASAP7_75t_L g3134 ( 
.A1(n_2914),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.C(n_105),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_2894),
.A2(n_106),
.B1(n_102),
.B2(n_105),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_SL g3136 ( 
.A1(n_2863),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_3136)
);

AND2x4_ASAP7_75t_L g3137 ( 
.A(n_2816),
.B(n_108),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2907),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2863),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2907),
.B(n_112),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2795),
.B(n_112),
.Y(n_3141)
);

AOI221xp5_ASAP7_75t_L g3142 ( 
.A1(n_2906),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.C(n_116),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2851),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2868),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2872),
.Y(n_3145)
);

AND2x4_ASAP7_75t_L g3146 ( 
.A(n_2795),
.B(n_119),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2893),
.B(n_119),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_2927),
.A2(n_2791),
.B1(n_2947),
.B2(n_2815),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2927),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2778),
.A2(n_1415),
.B(n_1207),
.Y(n_3150)
);

BUFx4f_ASAP7_75t_SL g3151 ( 
.A(n_2948),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2811),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_3152)
);

OR2x6_ASAP7_75t_L g3153 ( 
.A(n_2795),
.B(n_2815),
.Y(n_3153)
);

INVx3_ASAP7_75t_L g3154 ( 
.A(n_3153),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3085),
.Y(n_3155)
);

AO21x2_ASAP7_75t_L g3156 ( 
.A1(n_3096),
.A2(n_2747),
.B(n_2840),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_3127),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2974),
.Y(n_3158)
);

AO21x2_ASAP7_75t_L g3159 ( 
.A1(n_3096),
.A2(n_2840),
.B(n_2758),
.Y(n_3159)
);

BUFx3_ASAP7_75t_L g3160 ( 
.A(n_3102),
.Y(n_3160)
);

OAI21x1_ASAP7_75t_L g3161 ( 
.A1(n_2999),
.A2(n_2777),
.B(n_2758),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2988),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_3127),
.Y(n_3163)
);

INVxp67_ASAP7_75t_SL g3164 ( 
.A(n_2968),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_3042),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2998),
.Y(n_3166)
);

AO21x2_ASAP7_75t_L g3167 ( 
.A1(n_3069),
.A2(n_2736),
.B(n_2738),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3007),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2968),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_3153),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2976),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2991),
.Y(n_3172)
);

BUFx6f_ASAP7_75t_L g3173 ( 
.A(n_2997),
.Y(n_3173)
);

INVx3_ASAP7_75t_L g3174 ( 
.A(n_3153),
.Y(n_3174)
);

OA21x2_ASAP7_75t_L g3175 ( 
.A1(n_3150),
.A2(n_2777),
.B(n_2756),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3010),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3013),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_3027),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3030),
.Y(n_3179)
);

OR2x2_ASAP7_75t_L g3180 ( 
.A(n_2963),
.B(n_2813),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_3124),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3037),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_3035),
.B(n_3036),
.Y(n_3183)
);

AO21x1_ASAP7_75t_SL g3184 ( 
.A1(n_3099),
.A2(n_2799),
.B(n_2864),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_3138),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2963),
.B(n_2878),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3038),
.Y(n_3187)
);

AND3x2_ASAP7_75t_L g3188 ( 
.A(n_2961),
.B(n_3070),
.C(n_3082),
.Y(n_3188)
);

INVx3_ASAP7_75t_L g3189 ( 
.A(n_2997),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3126),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_2980),
.B(n_2815),
.Y(n_3191)
);

BUFx3_ASAP7_75t_L g3192 ( 
.A(n_3103),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_3039),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2995),
.B(n_2757),
.Y(n_3194)
);

AND2x4_ASAP7_75t_L g3195 ( 
.A(n_3035),
.B(n_2757),
.Y(n_3195)
);

HB1xp67_ASAP7_75t_L g3196 ( 
.A(n_3042),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3079),
.B(n_2813),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_L g3198 ( 
.A(n_3040),
.B(n_2915),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3068),
.Y(n_3199)
);

BUFx2_ASAP7_75t_L g3200 ( 
.A(n_3078),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3059),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3075),
.Y(n_3202)
);

AO21x2_ASAP7_75t_L g3203 ( 
.A1(n_3069),
.A2(n_2736),
.B(n_2738),
.Y(n_3203)
);

BUFx4f_ASAP7_75t_SL g3204 ( 
.A(n_2964),
.Y(n_3204)
);

BUFx2_ASAP7_75t_L g3205 ( 
.A(n_3011),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3077),
.Y(n_3206)
);

OA21x2_ASAP7_75t_L g3207 ( 
.A1(n_3150),
.A2(n_2827),
.B(n_2751),
.Y(n_3207)
);

BUFx3_ASAP7_75t_L g3208 ( 
.A(n_3088),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3025),
.B(n_2757),
.Y(n_3209)
);

HB1xp67_ASAP7_75t_L g3210 ( 
.A(n_3018),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3067),
.Y(n_3211)
);

INVx2_ASAP7_75t_SL g3212 ( 
.A(n_3018),
.Y(n_3212)
);

OA21x2_ASAP7_75t_L g3213 ( 
.A1(n_3148),
.A2(n_3084),
.B(n_2992),
.Y(n_3213)
);

HB1xp67_ASAP7_75t_L g3214 ( 
.A(n_3079),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3092),
.Y(n_3215)
);

INVx5_ASAP7_75t_L g3216 ( 
.A(n_2959),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_3011),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_3057),
.Y(n_3218)
);

BUFx4f_ASAP7_75t_L g3219 ( 
.A(n_3118),
.Y(n_3219)
);

HB1xp67_ASAP7_75t_L g3220 ( 
.A(n_3100),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3097),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3080),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_2970),
.B(n_2821),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3144),
.Y(n_3224)
);

OAI21x1_ASAP7_75t_L g3225 ( 
.A1(n_3057),
.A2(n_2762),
.B(n_2760),
.Y(n_3225)
);

AOI21x1_ASAP7_75t_L g3226 ( 
.A1(n_3132),
.A2(n_2871),
.B(n_2860),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3143),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3145),
.Y(n_3228)
);

OAI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2971),
.A2(n_2923),
.B(n_2899),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_3036),
.B(n_2881),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3111),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3125),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3100),
.Y(n_3233)
);

AO21x1_ASAP7_75t_SL g3234 ( 
.A1(n_2992),
.A2(n_2892),
.B(n_2889),
.Y(n_3234)
);

AO21x2_ASAP7_75t_L g3235 ( 
.A1(n_3114),
.A2(n_2746),
.B(n_2762),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_3023),
.B(n_2821),
.Y(n_3236)
);

HB1xp67_ASAP7_75t_L g3237 ( 
.A(n_3054),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3117),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3034),
.Y(n_3239)
);

OR2x2_ASAP7_75t_L g3240 ( 
.A(n_3054),
.B(n_2813),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3117),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3094),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3023),
.B(n_2813),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3044),
.Y(n_3244)
);

NOR2x1_ASAP7_75t_L g3245 ( 
.A(n_3104),
.B(n_2860),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3026),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3026),
.Y(n_3247)
);

INVx1_ASAP7_75t_SL g3248 ( 
.A(n_3006),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3001),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3147),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3001),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3006),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3121),
.Y(n_3253)
);

OR2x2_ASAP7_75t_L g3254 ( 
.A(n_3009),
.B(n_2827),
.Y(n_3254)
);

NAND2x1_ASAP7_75t_L g3255 ( 
.A(n_2966),
.B(n_2860),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_2983),
.A2(n_2985),
.B1(n_3070),
.B2(n_3152),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3121),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3131),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3131),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3140),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_3012),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3140),
.Y(n_3262)
);

HB1xp67_ASAP7_75t_L g3263 ( 
.A(n_3052),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2978),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_3009),
.B(n_2857),
.Y(n_3265)
);

OR2x2_ASAP7_75t_L g3266 ( 
.A(n_3119),
.B(n_2749),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2981),
.B(n_2911),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3048),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3128),
.Y(n_3269)
);

INVx3_ASAP7_75t_L g3270 ( 
.A(n_3012),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3116),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3060),
.Y(n_3272)
);

INVx2_ASAP7_75t_SL g3273 ( 
.A(n_3045),
.Y(n_3273)
);

INVx1_ASAP7_75t_SL g3274 ( 
.A(n_3072),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3060),
.Y(n_3275)
);

INVxp33_ASAP7_75t_L g3276 ( 
.A(n_3005),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3062),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3116),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3141),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3141),
.Y(n_3280)
);

OAI21x1_ASAP7_75t_L g3281 ( 
.A1(n_3110),
.A2(n_2760),
.B(n_2759),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3071),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3146),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3146),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3024),
.B(n_2871),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3110),
.A2(n_2759),
.B(n_2755),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2973),
.Y(n_3287)
);

BUFx3_ASAP7_75t_L g3288 ( 
.A(n_3087),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_3046),
.B(n_2779),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3047),
.B(n_2857),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3045),
.B(n_3058),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_3015),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_3015),
.Y(n_3293)
);

INVx3_ASAP7_75t_L g3294 ( 
.A(n_2989),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3058),
.B(n_2779),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2973),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2973),
.Y(n_3297)
);

HB1xp67_ASAP7_75t_L g3298 ( 
.A(n_3086),
.Y(n_3298)
);

HB1xp67_ASAP7_75t_L g3299 ( 
.A(n_3086),
.Y(n_3299)
);

INVxp33_ASAP7_75t_L g3300 ( 
.A(n_2990),
.Y(n_3300)
);

INVxp67_ASAP7_75t_L g3301 ( 
.A(n_2984),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3047),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_2985),
.A2(n_2749),
.B1(n_2847),
.B2(n_2842),
.Y(n_3303)
);

HB1xp67_ASAP7_75t_L g3304 ( 
.A(n_3108),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3108),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3020),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3123),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3002),
.B(n_3017),
.Y(n_3308)
);

OAI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3074),
.A2(n_2899),
.B(n_2897),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3020),
.B(n_2830),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_2989),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3112),
.Y(n_3312)
);

CKINVDCx5p33_ASAP7_75t_R g3313 ( 
.A(n_3019),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3231),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3248),
.B(n_3105),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_L g3316 ( 
.A1(n_3256),
.A2(n_3074),
.B1(n_3049),
.B2(n_3134),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3188),
.A2(n_3134),
.B1(n_3095),
.B2(n_3098),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3305),
.Y(n_3318)
);

AOI221xp5_ASAP7_75t_L g3319 ( 
.A1(n_3229),
.A2(n_3016),
.B1(n_3130),
.B2(n_3091),
.C(n_3142),
.Y(n_3319)
);

AOI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3303),
.A2(n_2994),
.B1(n_3055),
.B2(n_3106),
.Y(n_3320)
);

OAI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3229),
.A2(n_3029),
.B1(n_3129),
.B2(n_3149),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3309),
.A2(n_3095),
.B1(n_2994),
.B2(n_2982),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3305),
.Y(n_3323)
);

AO31x2_ASAP7_75t_L g3324 ( 
.A1(n_3290),
.A2(n_3081),
.A3(n_3113),
.B(n_2818),
.Y(n_3324)
);

OAI221xp5_ASAP7_75t_L g3325 ( 
.A1(n_3309),
.A2(n_3091),
.B1(n_2969),
.B2(n_3142),
.C(n_3029),
.Y(n_3325)
);

OR2x6_ASAP7_75t_L g3326 ( 
.A(n_3232),
.B(n_2960),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3232),
.A2(n_3004),
.B1(n_2993),
.B2(n_3136),
.Y(n_3327)
);

OAI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_3232),
.A2(n_3008),
.B1(n_3114),
.B2(n_2975),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3302),
.A2(n_2982),
.B1(n_3122),
.B2(n_3136),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3183),
.B(n_2960),
.Y(n_3330)
);

OAI21x1_ASAP7_75t_L g3331 ( 
.A1(n_3255),
.A2(n_2755),
.B(n_2785),
.Y(n_3331)
);

AOI21x1_ASAP7_75t_L g3332 ( 
.A1(n_3200),
.A2(n_3137),
.B(n_3133),
.Y(n_3332)
);

OAI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_3232),
.A2(n_3083),
.B1(n_3022),
.B2(n_3063),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3183),
.B(n_2967),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3305),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_3302),
.A2(n_3093),
.B1(n_2972),
.B2(n_3139),
.Y(n_3336)
);

AOI221xp5_ASAP7_75t_L g3337 ( 
.A1(n_3290),
.A2(n_3253),
.B1(n_3260),
.B2(n_3259),
.C(n_3258),
.Y(n_3337)
);

OAI221xp5_ASAP7_75t_L g3338 ( 
.A1(n_3200),
.A2(n_3265),
.B1(n_3267),
.B2(n_3253),
.C(n_3260),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3245),
.A2(n_3051),
.B(n_3028),
.Y(n_3339)
);

BUFx4f_ASAP7_75t_SL g3340 ( 
.A(n_3288),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_3250),
.A2(n_3043),
.B1(n_2972),
.B2(n_3051),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3183),
.B(n_2967),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3231),
.Y(n_3343)
);

AOI22xp33_ASAP7_75t_L g3344 ( 
.A1(n_3250),
.A2(n_3043),
.B1(n_2979),
.B2(n_3028),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3250),
.A2(n_3014),
.B1(n_2986),
.B2(n_3065),
.Y(n_3345)
);

AOI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3242),
.A2(n_3115),
.B1(n_3101),
.B2(n_2987),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3178),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_3232),
.A2(n_3041),
.B1(n_3032),
.B2(n_3003),
.Y(n_3348)
);

OAI221xp5_ASAP7_75t_L g3349 ( 
.A1(n_3265),
.A2(n_3033),
.B1(n_3135),
.B2(n_2965),
.C(n_2966),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_3242),
.A2(n_3118),
.B1(n_3021),
.B2(n_3003),
.Y(n_3350)
);

OAI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3232),
.A2(n_3151),
.B1(n_3118),
.B2(n_3120),
.Y(n_3351)
);

AOI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_3242),
.A2(n_3151),
.B1(n_3064),
.B2(n_2977),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_3248),
.B(n_2912),
.Y(n_3353)
);

HB1xp67_ASAP7_75t_L g3354 ( 
.A(n_3214),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3183),
.B(n_3308),
.Y(n_3355)
);

HB1xp67_ASAP7_75t_L g3356 ( 
.A(n_3165),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3308),
.B(n_2962),
.Y(n_3357)
);

INVx3_ASAP7_75t_L g3358 ( 
.A(n_3294),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3231),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3245),
.A2(n_3133),
.B1(n_3137),
.B2(n_2850),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_3269),
.B(n_2917),
.Y(n_3361)
);

OAI22xp5_ASAP7_75t_L g3362 ( 
.A1(n_3279),
.A2(n_3053),
.B1(n_3056),
.B2(n_2959),
.Y(n_3362)
);

OAI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_3300),
.A2(n_2959),
.B1(n_3061),
.B2(n_3113),
.Y(n_3363)
);

OA21x2_ASAP7_75t_L g3364 ( 
.A1(n_3296),
.A2(n_2785),
.B(n_2753),
.Y(n_3364)
);

INVx1_ASAP7_75t_SL g3365 ( 
.A(n_3204),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3178),
.Y(n_3366)
);

INVx3_ASAP7_75t_L g3367 ( 
.A(n_3294),
.Y(n_3367)
);

OAI21x1_ASAP7_75t_L g3368 ( 
.A1(n_3255),
.A2(n_3225),
.B(n_3226),
.Y(n_3368)
);

AOI22xp33_ASAP7_75t_L g3369 ( 
.A1(n_3213),
.A2(n_3269),
.B1(n_3184),
.B2(n_3252),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3182),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3279),
.A2(n_2959),
.B1(n_3066),
.B2(n_3090),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3279),
.A2(n_3050),
.B1(n_3109),
.B2(n_3107),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3182),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3213),
.A2(n_3269),
.B1(n_3184),
.B2(n_3252),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3213),
.A2(n_3000),
.B1(n_3031),
.B2(n_2847),
.Y(n_3375)
);

OR2x2_ASAP7_75t_L g3376 ( 
.A(n_3266),
.B(n_2919),
.Y(n_3376)
);

NAND3xp33_ASAP7_75t_L g3377 ( 
.A(n_3258),
.B(n_2996),
.C(n_3089),
.Y(n_3377)
);

OAI211xp5_ASAP7_75t_L g3378 ( 
.A1(n_3213),
.A2(n_3226),
.B(n_3266),
.C(n_3262),
.Y(n_3378)
);

OAI21x1_ASAP7_75t_L g3379 ( 
.A1(n_3225),
.A2(n_2753),
.B(n_2800),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3178),
.Y(n_3380)
);

OA21x2_ASAP7_75t_L g3381 ( 
.A1(n_3296),
.A2(n_2800),
.B(n_2765),
.Y(n_3381)
);

AOI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3249),
.A2(n_3251),
.B1(n_3262),
.B2(n_3259),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3280),
.A2(n_2847),
.B1(n_2901),
.B2(n_2837),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3312),
.A2(n_2850),
.B1(n_2962),
.B2(n_2897),
.Y(n_3384)
);

OAI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3280),
.A2(n_2847),
.B1(n_3076),
.B2(n_3073),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_3276),
.A2(n_2996),
.B(n_2882),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3178),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_SL g3388 ( 
.A1(n_3208),
.A2(n_3198),
.B1(n_3288),
.B2(n_3216),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_SL g3389 ( 
.A1(n_3208),
.A2(n_2882),
.B1(n_2865),
.B2(n_2929),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3249),
.B(n_2922),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3280),
.A2(n_3284),
.B1(n_3283),
.B2(n_3278),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_3154),
.B(n_2962),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3251),
.A2(n_3278),
.B1(n_3271),
.B2(n_3283),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3312),
.A2(n_2865),
.B1(n_2929),
.B2(n_2737),
.Y(n_3394)
);

OAI211xp5_ASAP7_75t_L g3395 ( 
.A1(n_3218),
.A2(n_2926),
.B(n_2818),
.C(n_2905),
.Y(n_3395)
);

OA21x2_ASAP7_75t_L g3396 ( 
.A1(n_3297),
.A2(n_2765),
.B(n_2781),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3187),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3187),
.Y(n_3398)
);

AOI221xp5_ASAP7_75t_L g3399 ( 
.A1(n_3257),
.A2(n_3301),
.B1(n_3186),
.B2(n_3289),
.C(n_3244),
.Y(n_3399)
);

OAI221xp5_ASAP7_75t_L g3400 ( 
.A1(n_3218),
.A2(n_2910),
.B1(n_2901),
.B2(n_2837),
.C(n_2830),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3194),
.B(n_2737),
.Y(n_3401)
);

HB1xp67_ASAP7_75t_L g3402 ( 
.A(n_3196),
.Y(n_3402)
);

INVxp67_ASAP7_75t_L g3403 ( 
.A(n_3210),
.Y(n_3403)
);

OAI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_3283),
.A2(n_2910),
.B1(n_2876),
.B2(n_2743),
.Y(n_3404)
);

OR2x2_ASAP7_75t_L g3405 ( 
.A(n_3264),
.B(n_2802),
.Y(n_3405)
);

OAI33xp33_ASAP7_75t_L g3406 ( 
.A1(n_3197),
.A2(n_123),
.A3(n_125),
.B1(n_126),
.B2(n_127),
.B3(n_129),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3194),
.B(n_2809),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3199),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_SL g3409 ( 
.A1(n_3208),
.A2(n_2858),
.B1(n_2938),
.B2(n_2937),
.Y(n_3409)
);

AOI21xp33_ASAP7_75t_L g3410 ( 
.A1(n_3257),
.A2(n_2740),
.B(n_2937),
.Y(n_3410)
);

BUFx6f_ASAP7_75t_L g3411 ( 
.A(n_3160),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3199),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_3311),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3284),
.A2(n_2743),
.B1(n_2796),
.B2(n_2853),
.Y(n_3414)
);

OAI221xp5_ASAP7_75t_L g3415 ( 
.A1(n_3257),
.A2(n_2743),
.B1(n_127),
.B2(n_130),
.C(n_131),
.Y(n_3415)
);

INVx4_ASAP7_75t_L g3416 ( 
.A(n_3160),
.Y(n_3416)
);

AOI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3288),
.A2(n_2938),
.B1(n_2858),
.B2(n_2939),
.Y(n_3417)
);

OAI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3284),
.A2(n_2796),
.B1(n_2916),
.B2(n_2958),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3220),
.Y(n_3419)
);

OAI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3271),
.A2(n_2796),
.B1(n_2916),
.B2(n_2958),
.Y(n_3420)
);

INVx3_ASAP7_75t_L g3421 ( 
.A(n_3294),
.Y(n_3421)
);

OAI22xp5_ASAP7_75t_SL g3422 ( 
.A1(n_3160),
.A2(n_2946),
.B1(n_2950),
.B2(n_2939),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3311),
.Y(n_3423)
);

OAI211xp5_ASAP7_75t_L g3424 ( 
.A1(n_3254),
.A2(n_2950),
.B(n_2956),
.C(n_2946),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3271),
.A2(n_2916),
.B1(n_2956),
.B2(n_2854),
.Y(n_3425)
);

NAND3xp33_ASAP7_75t_L g3426 ( 
.A(n_3254),
.B(n_3295),
.C(n_3155),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3202),
.Y(n_3427)
);

OAI22xp33_ASAP7_75t_L g3428 ( 
.A1(n_3278),
.A2(n_2916),
.B1(n_2921),
.B2(n_2924),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3235),
.A2(n_2924),
.B1(n_2921),
.B2(n_2854),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3235),
.A2(n_2809),
.B1(n_2861),
.B2(n_2797),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3235),
.A2(n_2861),
.B1(n_2797),
.B2(n_2781),
.Y(n_3431)
);

AOI221xp5_ASAP7_75t_L g3432 ( 
.A1(n_3289),
.A2(n_125),
.B1(n_132),
.B2(n_134),
.C(n_135),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3219),
.A2(n_3306),
.B1(n_3192),
.B2(n_3233),
.Y(n_3433)
);

OAI221xp5_ASAP7_75t_L g3434 ( 
.A1(n_3205),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.C(n_137),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3237),
.B(n_2802),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_3235),
.A2(n_2772),
.B(n_2789),
.Y(n_3436)
);

OAI21x1_ASAP7_75t_L g3437 ( 
.A1(n_3161),
.A2(n_2772),
.B(n_2773),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3219),
.A2(n_2789),
.B(n_2773),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_SL g3439 ( 
.A1(n_3216),
.A2(n_2780),
.B1(n_138),
.B2(n_136),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3202),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3311),
.Y(n_3441)
);

INVx2_ASAP7_75t_SL g3442 ( 
.A(n_3192),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_3219),
.A2(n_2802),
.B1(n_2803),
.B2(n_2895),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3306),
.A2(n_2780),
.B1(n_2803),
.B2(n_2802),
.Y(n_3444)
);

OAI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3161),
.A2(n_2895),
.B(n_137),
.Y(n_3445)
);

OAI21xp33_ASAP7_75t_L g3446 ( 
.A1(n_3285),
.A2(n_138),
.B(n_139),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3370),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3373),
.Y(n_3448)
);

NAND3xp33_ASAP7_75t_L g3449 ( 
.A(n_3322),
.B(n_3297),
.C(n_3295),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3397),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3355),
.B(n_3154),
.Y(n_3451)
);

AND2x4_ASAP7_75t_L g3452 ( 
.A(n_3392),
.B(n_3154),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3341),
.B(n_3307),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3392),
.B(n_3154),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3318),
.Y(n_3455)
);

INVx3_ASAP7_75t_SL g3456 ( 
.A(n_3416),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3398),
.Y(n_3457)
);

INVxp67_ASAP7_75t_L g3458 ( 
.A(n_3377),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3408),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3323),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3412),
.Y(n_3461)
);

NOR2xp67_ASAP7_75t_L g3462 ( 
.A(n_3416),
.B(n_3170),
.Y(n_3462)
);

INVxp67_ASAP7_75t_L g3463 ( 
.A(n_3326),
.Y(n_3463)
);

INVxp67_ASAP7_75t_L g3464 ( 
.A(n_3326),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3335),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3330),
.B(n_3170),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3382),
.B(n_3315),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3334),
.B(n_3170),
.Y(n_3468)
);

INVx4_ASAP7_75t_SL g3469 ( 
.A(n_3411),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3342),
.B(n_3170),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3388),
.B(n_3174),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3427),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3337),
.B(n_3388),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3369),
.B(n_3174),
.Y(n_3474)
);

INVx4_ASAP7_75t_R g3475 ( 
.A(n_3442),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3440),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_3326),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3361),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3374),
.B(n_3174),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3356),
.B(n_3240),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3354),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3354),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3393),
.B(n_3386),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3357),
.B(n_3174),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3399),
.B(n_3307),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3314),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3343),
.Y(n_3487)
);

INVx2_ASAP7_75t_SL g3488 ( 
.A(n_3411),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3403),
.B(n_3307),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3401),
.B(n_3358),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3358),
.B(n_3261),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3347),
.Y(n_3492)
);

AOI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_3319),
.A2(n_3310),
.B1(n_3233),
.B2(n_3264),
.Y(n_3493)
);

NOR2x1_ASAP7_75t_SL g3494 ( 
.A(n_3332),
.B(n_3234),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3403),
.B(n_3285),
.Y(n_3495)
);

INVxp67_ASAP7_75t_L g3496 ( 
.A(n_3349),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3367),
.B(n_3261),
.Y(n_3497)
);

OR2x2_ASAP7_75t_L g3498 ( 
.A(n_3356),
.B(n_3402),
.Y(n_3498)
);

HB1xp67_ASAP7_75t_L g3499 ( 
.A(n_3402),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3366),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3390),
.Y(n_3501)
);

BUFx3_ASAP7_75t_L g3502 ( 
.A(n_3411),
.Y(n_3502)
);

CKINVDCx5p33_ASAP7_75t_R g3503 ( 
.A(n_3340),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3380),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3419),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3353),
.Y(n_3506)
);

INVx2_ASAP7_75t_SL g3507 ( 
.A(n_3411),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3367),
.B(n_3261),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3316),
.A2(n_3219),
.B1(n_3192),
.B2(n_3261),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3421),
.B(n_3270),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3359),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3387),
.Y(n_3512)
);

OR2x2_ASAP7_75t_L g3513 ( 
.A(n_3435),
.B(n_3240),
.Y(n_3513)
);

OAI222xp33_ASAP7_75t_L g3514 ( 
.A1(n_3325),
.A2(n_3320),
.B1(n_3328),
.B2(n_3339),
.C1(n_3321),
.C2(n_3317),
.Y(n_3514)
);

OR2x2_ASAP7_75t_L g3515 ( 
.A(n_3376),
.B(n_3180),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3421),
.B(n_3270),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3413),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3407),
.B(n_3423),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3441),
.B(n_3270),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3391),
.B(n_3270),
.Y(n_3520)
);

NOR2x1_ASAP7_75t_L g3521 ( 
.A(n_3363),
.B(n_3189),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3375),
.B(n_3292),
.Y(n_3522)
);

BUFx3_ASAP7_75t_L g3523 ( 
.A(n_3340),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3368),
.Y(n_3524)
);

HB1xp67_ASAP7_75t_L g3525 ( 
.A(n_3324),
.Y(n_3525)
);

OR2x2_ASAP7_75t_L g3526 ( 
.A(n_3324),
.B(n_3180),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3328),
.A2(n_3173),
.B1(n_3217),
.B2(n_3205),
.Y(n_3527)
);

OR2x2_ASAP7_75t_L g3528 ( 
.A(n_3324),
.B(n_3155),
.Y(n_3528)
);

HB1xp67_ASAP7_75t_L g3529 ( 
.A(n_3324),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3405),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3433),
.B(n_3292),
.Y(n_3531)
);

HB1xp67_ASAP7_75t_L g3532 ( 
.A(n_3362),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3345),
.B(n_3264),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3381),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3378),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3381),
.Y(n_3536)
);

OR2x2_ASAP7_75t_L g3537 ( 
.A(n_3426),
.B(n_3155),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3445),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3418),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3420),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3344),
.B(n_3244),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3396),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3446),
.B(n_3268),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3415),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3372),
.B(n_3292),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3425),
.Y(n_3546)
);

BUFx2_ASAP7_75t_L g3547 ( 
.A(n_3363),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3360),
.B(n_3292),
.Y(n_3548)
);

INVx2_ASAP7_75t_SL g3549 ( 
.A(n_3365),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3360),
.B(n_3293),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3396),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3352),
.B(n_3293),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3329),
.B(n_3268),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3364),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3329),
.B(n_3212),
.Y(n_3555)
);

BUFx3_ASAP7_75t_L g3556 ( 
.A(n_3422),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_3346),
.Y(n_3557)
);

AND2x4_ASAP7_75t_SL g3558 ( 
.A(n_3417),
.B(n_3209),
.Y(n_3558)
);

NAND3xp33_ASAP7_75t_L g3559 ( 
.A(n_3432),
.B(n_3173),
.C(n_3238),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3336),
.A2(n_3293),
.B1(n_3195),
.B2(n_3216),
.Y(n_3560)
);

OAI222xp33_ASAP7_75t_L g3561 ( 
.A1(n_3338),
.A2(n_3217),
.B1(n_3274),
.B2(n_3189),
.C1(n_3272),
.C2(n_3275),
.Y(n_3561)
);

INVxp67_ASAP7_75t_L g3562 ( 
.A(n_3348),
.Y(n_3562)
);

OR2x2_ASAP7_75t_L g3563 ( 
.A(n_3395),
.B(n_3212),
.Y(n_3563)
);

INVxp67_ASAP7_75t_L g3564 ( 
.A(n_3327),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3385),
.Y(n_3565)
);

OR2x2_ASAP7_75t_L g3566 ( 
.A(n_3414),
.B(n_3197),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3371),
.B(n_3293),
.Y(n_3567)
);

HB1xp67_ASAP7_75t_L g3568 ( 
.A(n_3404),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3364),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3384),
.B(n_3223),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3336),
.B(n_3239),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3331),
.Y(n_3572)
);

HB1xp67_ASAP7_75t_L g3573 ( 
.A(n_3400),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3434),
.B(n_3313),
.Y(n_3574)
);

AO21x2_ASAP7_75t_L g3575 ( 
.A1(n_3535),
.A2(n_3436),
.B(n_3351),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3514),
.A2(n_3406),
.B(n_3333),
.Y(n_3576)
);

OAI33xp33_ASAP7_75t_L g3577 ( 
.A1(n_3458),
.A2(n_3333),
.A3(n_3351),
.B1(n_3385),
.B2(n_3406),
.B3(n_3428),
.Y(n_3577)
);

AO21x2_ASAP7_75t_L g3578 ( 
.A1(n_3473),
.A2(n_3163),
.B(n_3157),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3544),
.B(n_3223),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3496),
.A2(n_3439),
.B1(n_3389),
.B2(n_3350),
.Y(n_3580)
);

OA21x2_ASAP7_75t_L g3581 ( 
.A1(n_3449),
.A2(n_3163),
.B(n_3157),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3447),
.Y(n_3582)
);

BUFx3_ASAP7_75t_L g3583 ( 
.A(n_3523),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3484),
.B(n_3195),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3484),
.B(n_3195),
.Y(n_3585)
);

OR2x2_ASAP7_75t_L g3586 ( 
.A(n_3571),
.B(n_3239),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_3454),
.B(n_3195),
.Y(n_3587)
);

AOI222xp33_ASAP7_75t_L g3588 ( 
.A1(n_3564),
.A2(n_3562),
.B1(n_3559),
.B2(n_3555),
.C1(n_3483),
.C2(n_3547),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3453),
.B(n_3277),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3454),
.B(n_3246),
.Y(n_3590)
);

AOI222xp33_ASAP7_75t_L g3591 ( 
.A1(n_3547),
.A2(n_3384),
.B1(n_3429),
.B2(n_3430),
.C1(n_3394),
.C2(n_3424),
.Y(n_3591)
);

OAI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3527),
.A2(n_3439),
.B(n_3410),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3557),
.A2(n_3389),
.B1(n_3429),
.B2(n_3409),
.Y(n_3593)
);

AND2x2_ASAP7_75t_SL g3594 ( 
.A(n_3477),
.B(n_3417),
.Y(n_3594)
);

NAND3xp33_ASAP7_75t_L g3595 ( 
.A(n_3532),
.B(n_3430),
.C(n_3431),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3452),
.B(n_3246),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3498),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3498),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3556),
.B(n_3173),
.Y(n_3599)
);

OR2x2_ASAP7_75t_L g3600 ( 
.A(n_3533),
.B(n_3263),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3452),
.B(n_3247),
.Y(n_3601)
);

INVxp67_ASAP7_75t_L g3602 ( 
.A(n_3477),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3447),
.Y(n_3603)
);

NAND3xp33_ASAP7_75t_L g3604 ( 
.A(n_3573),
.B(n_3431),
.C(n_3394),
.Y(n_3604)
);

BUFx2_ASAP7_75t_L g3605 ( 
.A(n_3523),
.Y(n_3605)
);

OA21x2_ASAP7_75t_L g3606 ( 
.A1(n_3542),
.A2(n_3163),
.B(n_3157),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3452),
.B(n_3247),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_3549),
.B(n_3503),
.Y(n_3608)
);

OR2x2_ASAP7_75t_L g3609 ( 
.A(n_3485),
.B(n_3274),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3519),
.Y(n_3610)
);

AND2x4_ASAP7_75t_L g3611 ( 
.A(n_3469),
.B(n_3189),
.Y(n_3611)
);

AOI221xp5_ASAP7_75t_L g3612 ( 
.A1(n_3556),
.A2(n_3428),
.B1(n_3221),
.B2(n_3215),
.C(n_3206),
.Y(n_3612)
);

AOI221xp5_ASAP7_75t_L g3613 ( 
.A1(n_3546),
.A2(n_3540),
.B1(n_3539),
.B2(n_3561),
.C(n_3560),
.Y(n_3613)
);

AO21x2_ASAP7_75t_L g3614 ( 
.A1(n_3525),
.A2(n_3287),
.B(n_3156),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3461),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3461),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3557),
.A2(n_3409),
.B1(n_3159),
.B2(n_3156),
.Y(n_3617)
);

BUFx3_ASAP7_75t_L g3618 ( 
.A(n_3503),
.Y(n_3618)
);

AO21x1_ASAP7_75t_SL g3619 ( 
.A1(n_3563),
.A2(n_3275),
.B(n_3272),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3499),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3519),
.Y(n_3621)
);

NAND3xp33_ASAP7_75t_L g3622 ( 
.A(n_3568),
.B(n_3444),
.C(n_3173),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3528),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3466),
.B(n_3209),
.Y(n_3624)
);

INVxp67_ASAP7_75t_L g3625 ( 
.A(n_3505),
.Y(n_3625)
);

NOR2x1_ASAP7_75t_SL g3626 ( 
.A(n_3563),
.B(n_3234),
.Y(n_3626)
);

AO21x2_ASAP7_75t_L g3627 ( 
.A1(n_3529),
.A2(n_3287),
.B(n_3156),
.Y(n_3627)
);

INVx8_ASAP7_75t_L g3628 ( 
.A(n_3469),
.Y(n_3628)
);

NOR2x1_ASAP7_75t_L g3629 ( 
.A(n_3502),
.B(n_3189),
.Y(n_3629)
);

BUFx2_ASAP7_75t_L g3630 ( 
.A(n_3469),
.Y(n_3630)
);

NAND3xp33_ASAP7_75t_L g3631 ( 
.A(n_3565),
.B(n_3173),
.C(n_3438),
.Y(n_3631)
);

OAI221xp5_ASAP7_75t_L g3632 ( 
.A1(n_3493),
.A2(n_3173),
.B1(n_3164),
.B2(n_3287),
.C(n_3273),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3549),
.B(n_3206),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3448),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3450),
.Y(n_3635)
);

CKINVDCx20_ASAP7_75t_R g3636 ( 
.A(n_3574),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3457),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_SL g3638 ( 
.A1(n_3494),
.A2(n_3216),
.B1(n_3159),
.B2(n_3156),
.Y(n_3638)
);

BUFx2_ASAP7_75t_L g3639 ( 
.A(n_3469),
.Y(n_3639)
);

NAND3xp33_ASAP7_75t_L g3640 ( 
.A(n_3538),
.B(n_3216),
.C(n_3383),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_SL g3641 ( 
.A(n_3509),
.B(n_3216),
.Y(n_3641)
);

NOR4xp25_ASAP7_75t_SL g3642 ( 
.A(n_3481),
.B(n_3169),
.C(n_3216),
.D(n_3215),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3466),
.B(n_3191),
.Y(n_3643)
);

OR2x2_ASAP7_75t_L g3644 ( 
.A(n_3489),
.B(n_3277),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_L g3645 ( 
.A1(n_3553),
.A2(n_3159),
.B1(n_3203),
.B2(n_3167),
.Y(n_3645)
);

OAI332xp33_ASAP7_75t_L g3646 ( 
.A1(n_3526),
.A2(n_3566),
.A3(n_3467),
.B1(n_3537),
.B2(n_3541),
.B3(n_3528),
.C1(n_3543),
.C2(n_3482),
.Y(n_3646)
);

NOR2xp67_ASAP7_75t_L g3647 ( 
.A(n_3462),
.B(n_3471),
.Y(n_3647)
);

OAI21xp33_ASAP7_75t_L g3648 ( 
.A1(n_3548),
.A2(n_3236),
.B(n_3243),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3534),
.Y(n_3649)
);

OAI221xp5_ASAP7_75t_L g3650 ( 
.A1(n_3521),
.A2(n_3273),
.B1(n_3294),
.B2(n_3221),
.C(n_3228),
.Y(n_3650)
);

OAI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3456),
.A2(n_3238),
.B1(n_3241),
.B2(n_3169),
.Y(n_3651)
);

AOI31xp33_ASAP7_75t_L g3652 ( 
.A1(n_3463),
.A2(n_3310),
.A3(n_3291),
.B(n_3191),
.Y(n_3652)
);

AOI221xp5_ASAP7_75t_L g3653 ( 
.A1(n_3570),
.A2(n_3464),
.B1(n_3550),
.B2(n_3548),
.C(n_3471),
.Y(n_3653)
);

NAND3xp33_ASAP7_75t_L g3654 ( 
.A(n_3474),
.B(n_3241),
.C(n_3238),
.Y(n_3654)
);

OAI221xp5_ASAP7_75t_L g3655 ( 
.A1(n_3456),
.A2(n_3224),
.B1(n_3228),
.B2(n_3282),
.C(n_3158),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3488),
.B(n_3282),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3506),
.B(n_3224),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3459),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3472),
.Y(n_3659)
);

INVx1_ASAP7_75t_SL g3660 ( 
.A(n_3502),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3468),
.B(n_3291),
.Y(n_3661)
);

OAI211xp5_ASAP7_75t_L g3662 ( 
.A1(n_3550),
.A2(n_3241),
.B(n_3175),
.C(n_3298),
.Y(n_3662)
);

INVx3_ASAP7_75t_L g3663 ( 
.A(n_3451),
.Y(n_3663)
);

NOR2xp67_ASAP7_75t_SL g3664 ( 
.A(n_3488),
.B(n_3299),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3468),
.B(n_3230),
.Y(n_3665)
);

INVxp67_ASAP7_75t_SL g3666 ( 
.A(n_3526),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3476),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3501),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_3480),
.Y(n_3669)
);

BUFx3_ASAP7_75t_L g3670 ( 
.A(n_3507),
.Y(n_3670)
);

HB1xp67_ASAP7_75t_L g3671 ( 
.A(n_3480),
.Y(n_3671)
);

AOI221xp5_ASAP7_75t_L g3672 ( 
.A1(n_3570),
.A2(n_3558),
.B1(n_3479),
.B2(n_3474),
.C(n_3478),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3534),
.Y(n_3673)
);

OA21x2_ASAP7_75t_L g3674 ( 
.A1(n_3542),
.A2(n_3551),
.B(n_3554),
.Y(n_3674)
);

INVx1_ASAP7_75t_SL g3675 ( 
.A(n_3507),
.Y(n_3675)
);

INVx3_ASAP7_75t_L g3676 ( 
.A(n_3451),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3470),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3486),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3470),
.B(n_3243),
.Y(n_3679)
);

INVx1_ASAP7_75t_SL g3680 ( 
.A(n_3552),
.Y(n_3680)
);

AO21x2_ASAP7_75t_L g3681 ( 
.A1(n_3494),
.A2(n_3159),
.B(n_3379),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3545),
.B(n_3230),
.Y(n_3682)
);

AOI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3558),
.A2(n_3158),
.B1(n_3162),
.B2(n_3168),
.C(n_3230),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3486),
.Y(n_3684)
);

AOI221xp5_ASAP7_75t_L g3685 ( 
.A1(n_3479),
.A2(n_3162),
.B1(n_3168),
.B2(n_3230),
.C(n_3236),
.Y(n_3685)
);

AOI221xp5_ASAP7_75t_L g3686 ( 
.A1(n_3566),
.A2(n_3179),
.B1(n_3172),
.B2(n_3177),
.C(n_3222),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3487),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3552),
.B(n_3193),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3522),
.B(n_3193),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_L g3690 ( 
.A1(n_3577),
.A2(n_3522),
.B1(n_3545),
.B2(n_3567),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3583),
.Y(n_3691)
);

OR2x2_ASAP7_75t_L g3692 ( 
.A(n_3680),
.B(n_3495),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3605),
.B(n_3531),
.Y(n_3693)
);

AO21x2_ASAP7_75t_L g3694 ( 
.A1(n_3666),
.A2(n_3524),
.B(n_3536),
.Y(n_3694)
);

NOR3xp33_ASAP7_75t_L g3695 ( 
.A(n_3646),
.B(n_3577),
.C(n_3576),
.Y(n_3695)
);

NAND3xp33_ASAP7_75t_L g3696 ( 
.A(n_3588),
.B(n_3593),
.C(n_3604),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3583),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3597),
.B(n_3517),
.Y(n_3698)
);

NAND3xp33_ASAP7_75t_L g3699 ( 
.A(n_3593),
.B(n_3524),
.C(n_3537),
.Y(n_3699)
);

INVxp67_ASAP7_75t_L g3700 ( 
.A(n_3608),
.Y(n_3700)
);

NAND3xp33_ASAP7_75t_L g3701 ( 
.A(n_3591),
.B(n_3530),
.C(n_3567),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3636),
.A2(n_3531),
.B1(n_3520),
.B2(n_3497),
.Y(n_3702)
);

OR2x2_ASAP7_75t_L g3703 ( 
.A(n_3609),
.B(n_3513),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_3618),
.B(n_3520),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3669),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3608),
.B(n_3490),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3587),
.B(n_3490),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3596),
.B(n_3518),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_L g3709 ( 
.A1(n_3594),
.A2(n_3595),
.B1(n_3592),
.B2(n_3575),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_L g3710 ( 
.A(n_3653),
.B(n_3513),
.C(n_3511),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3601),
.B(n_3518),
.Y(n_3711)
);

NAND4xp75_ASAP7_75t_L g3712 ( 
.A(n_3594),
.B(n_3475),
.C(n_3497),
.D(n_3491),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3597),
.B(n_3455),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_3630),
.B(n_3491),
.Y(n_3714)
);

NOR3xp33_ASAP7_75t_SL g3715 ( 
.A(n_3641),
.B(n_3511),
.C(n_3487),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3598),
.B(n_3455),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3607),
.B(n_3508),
.Y(n_3717)
);

AOI211xp5_ASAP7_75t_L g3718 ( 
.A1(n_3672),
.A2(n_3572),
.B(n_3551),
.C(n_3536),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3682),
.B(n_3508),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3618),
.B(n_3636),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3663),
.B(n_3510),
.Y(n_3721)
);

NOR3xp33_ASAP7_75t_SL g3722 ( 
.A(n_3641),
.B(n_3443),
.C(n_3177),
.Y(n_3722)
);

NAND3xp33_ASAP7_75t_L g3723 ( 
.A(n_3617),
.B(n_3465),
.C(n_3460),
.Y(n_3723)
);

INVx2_ASAP7_75t_SL g3724 ( 
.A(n_3628),
.Y(n_3724)
);

NAND4xp75_ASAP7_75t_L g3725 ( 
.A(n_3647),
.B(n_3516),
.C(n_3510),
.D(n_3572),
.Y(n_3725)
);

OR2x2_ASAP7_75t_L g3726 ( 
.A(n_3600),
.B(n_3460),
.Y(n_3726)
);

NOR3xp33_ASAP7_75t_L g3727 ( 
.A(n_3602),
.B(n_3569),
.C(n_3554),
.Y(n_3727)
);

INVx2_ASAP7_75t_SL g3728 ( 
.A(n_3628),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3663),
.B(n_3516),
.Y(n_3729)
);

OAI211xp5_ASAP7_75t_SL g3730 ( 
.A1(n_3580),
.A2(n_3569),
.B(n_3465),
.C(n_3500),
.Y(n_3730)
);

NAND4xp75_ASAP7_75t_L g3731 ( 
.A(n_3599),
.B(n_3492),
.C(n_3504),
.D(n_3500),
.Y(n_3731)
);

BUFx3_ASAP7_75t_L g3732 ( 
.A(n_3628),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3598),
.B(n_3492),
.Y(n_3733)
);

OAI211xp5_ASAP7_75t_L g3734 ( 
.A1(n_3580),
.A2(n_3175),
.B(n_3515),
.C(n_3512),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3575),
.A2(n_3512),
.B1(n_3504),
.B2(n_3167),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3676),
.B(n_3515),
.Y(n_3736)
);

OR2x2_ASAP7_75t_L g3737 ( 
.A(n_3579),
.B(n_3193),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3676),
.B(n_3304),
.Y(n_3738)
);

AOI211xp5_ASAP7_75t_L g3739 ( 
.A1(n_3622),
.A2(n_3437),
.B(n_3281),
.C(n_3286),
.Y(n_3739)
);

AND2x4_ASAP7_75t_L g3740 ( 
.A(n_3639),
.B(n_3201),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3625),
.B(n_3181),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3625),
.B(n_3181),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3586),
.B(n_3201),
.Y(n_3743)
);

NOR3xp33_ASAP7_75t_L g3744 ( 
.A(n_3602),
.B(n_3281),
.C(n_140),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3584),
.B(n_3201),
.Y(n_3745)
);

NAND3xp33_ASAP7_75t_L g3746 ( 
.A(n_3617),
.B(n_3175),
.C(n_3207),
.Y(n_3746)
);

NOR3xp33_ASAP7_75t_L g3747 ( 
.A(n_3613),
.B(n_140),
.C(n_141),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3612),
.B(n_3175),
.C(n_3207),
.Y(n_3748)
);

NAND3xp33_ASAP7_75t_L g3749 ( 
.A(n_3645),
.B(n_3207),
.C(n_3179),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_SL g3750 ( 
.A1(n_3626),
.A2(n_3167),
.B1(n_3203),
.B2(n_3207),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3585),
.B(n_3211),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3677),
.B(n_3211),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3669),
.Y(n_3753)
);

NAND3xp33_ASAP7_75t_L g3754 ( 
.A(n_3645),
.B(n_3172),
.C(n_3227),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_3660),
.B(n_3227),
.Y(n_3755)
);

NOR2x1_ASAP7_75t_L g3756 ( 
.A(n_3670),
.B(n_3599),
.Y(n_3756)
);

NOR3xp33_ASAP7_75t_L g3757 ( 
.A(n_3650),
.B(n_142),
.C(n_143),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3670),
.Y(n_3758)
);

AOI22xp33_ASAP7_75t_L g3759 ( 
.A1(n_3632),
.A2(n_3167),
.B1(n_3203),
.B2(n_3211),
.Y(n_3759)
);

OR2x2_ASAP7_75t_L g3760 ( 
.A(n_3589),
.B(n_3620),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3590),
.B(n_3222),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3624),
.B(n_3222),
.Y(n_3762)
);

NAND3xp33_ASAP7_75t_L g3763 ( 
.A(n_3631),
.B(n_3227),
.C(n_3185),
.Y(n_3763)
);

OR2x2_ASAP7_75t_L g3764 ( 
.A(n_3688),
.B(n_3181),
.Y(n_3764)
);

AND2x4_ASAP7_75t_L g3765 ( 
.A(n_3675),
.B(n_3166),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3668),
.B(n_3185),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3671),
.B(n_3185),
.Y(n_3767)
);

OAI211xp5_ASAP7_75t_SL g3768 ( 
.A1(n_3638),
.A2(n_3166),
.B(n_3190),
.C(n_3176),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3638),
.A2(n_3203),
.B1(n_3286),
.B2(n_3166),
.Y(n_3769)
);

INVx4_ASAP7_75t_L g3770 ( 
.A(n_3611),
.Y(n_3770)
);

AOI22xp33_ASAP7_75t_L g3771 ( 
.A1(n_3640),
.A2(n_3190),
.B1(n_3176),
.B2(n_3171),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3671),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3661),
.B(n_3171),
.Y(n_3773)
);

AND2x4_ASAP7_75t_L g3774 ( 
.A(n_3629),
.B(n_3171),
.Y(n_3774)
);

NAND3xp33_ASAP7_75t_L g3775 ( 
.A(n_3581),
.B(n_3190),
.C(n_3176),
.Y(n_3775)
);

NAND3xp33_ASAP7_75t_L g3776 ( 
.A(n_3581),
.B(n_142),
.C(n_144),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_SL g3777 ( 
.A(n_3652),
.B(n_2895),
.Y(n_3777)
);

NAND3xp33_ASAP7_75t_L g3778 ( 
.A(n_3581),
.B(n_145),
.C(n_146),
.Y(n_3778)
);

BUFx2_ASAP7_75t_L g3779 ( 
.A(n_3611),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3643),
.B(n_145),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3644),
.B(n_146),
.Y(n_3781)
);

HB1xp67_ASAP7_75t_L g3782 ( 
.A(n_3694),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3695),
.B(n_3633),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_L g3784 ( 
.A(n_3700),
.B(n_3633),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3705),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3695),
.B(n_3634),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3753),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3772),
.Y(n_3788)
);

AOI221xp5_ASAP7_75t_L g3789 ( 
.A1(n_3709),
.A2(n_3662),
.B1(n_3654),
.B2(n_3666),
.C(n_3685),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3694),
.Y(n_3790)
);

HB1xp67_ASAP7_75t_L g3791 ( 
.A(n_3776),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3779),
.Y(n_3792)
);

OAI31xp33_ASAP7_75t_L g3793 ( 
.A1(n_3696),
.A2(n_3651),
.A3(n_3648),
.B(n_3655),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3756),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3713),
.Y(n_3795)
);

INVx3_ASAP7_75t_L g3796 ( 
.A(n_3770),
.Y(n_3796)
);

NOR2xp67_ASAP7_75t_L g3797 ( 
.A(n_3770),
.B(n_3610),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3713),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3747),
.B(n_3635),
.Y(n_3799)
);

OAI21xp33_ASAP7_75t_L g3800 ( 
.A1(n_3747),
.A2(n_3689),
.B(n_3658),
.Y(n_3800)
);

OAI33xp33_ASAP7_75t_L g3801 ( 
.A1(n_3730),
.A2(n_3616),
.A3(n_3582),
.B1(n_3603),
.B2(n_3615),
.B3(n_3659),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3716),
.Y(n_3802)
);

INVxp67_ASAP7_75t_SL g3803 ( 
.A(n_3778),
.Y(n_3803)
);

OR2x2_ASAP7_75t_L g3804 ( 
.A(n_3692),
.B(n_3657),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3727),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_L g3806 ( 
.A(n_3700),
.B(n_3720),
.Y(n_3806)
);

INVx3_ASAP7_75t_L g3807 ( 
.A(n_3714),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3730),
.A2(n_3578),
.B1(n_3619),
.B2(n_3637),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3693),
.B(n_3665),
.Y(n_3809)
);

INVx2_ASAP7_75t_SL g3810 ( 
.A(n_3714),
.Y(n_3810)
);

INVx3_ASAP7_75t_L g3811 ( 
.A(n_3732),
.Y(n_3811)
);

INVx1_ASAP7_75t_SL g3812 ( 
.A(n_3706),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3716),
.Y(n_3813)
);

AOI22xp33_ASAP7_75t_L g3814 ( 
.A1(n_3757),
.A2(n_3578),
.B1(n_3667),
.B2(n_3683),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3691),
.B(n_3664),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3758),
.Y(n_3816)
);

BUFx2_ASAP7_75t_L g3817 ( 
.A(n_3697),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3690),
.B(n_3610),
.Y(n_3818)
);

OAI221xp5_ASAP7_75t_SL g3819 ( 
.A1(n_3734),
.A2(n_3651),
.B1(n_3686),
.B2(n_3621),
.C(n_3642),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3733),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3733),
.Y(n_3821)
);

AND2x4_ASAP7_75t_SL g3822 ( 
.A(n_3724),
.B(n_3621),
.Y(n_3822)
);

INVx3_ASAP7_75t_L g3823 ( 
.A(n_3774),
.Y(n_3823)
);

BUFx2_ASAP7_75t_L g3824 ( 
.A(n_3728),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3704),
.B(n_3679),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3698),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3760),
.B(n_3656),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3757),
.A2(n_3649),
.B1(n_3673),
.B2(n_3678),
.Y(n_3828)
);

OAI31xp33_ASAP7_75t_L g3829 ( 
.A1(n_3734),
.A2(n_3699),
.A3(n_3744),
.B(n_3701),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3717),
.B(n_3679),
.Y(n_3830)
);

INVx3_ASAP7_75t_L g3831 ( 
.A(n_3774),
.Y(n_3831)
);

INVx2_ASAP7_75t_SL g3832 ( 
.A(n_3721),
.Y(n_3832)
);

BUFx3_ASAP7_75t_L g3833 ( 
.A(n_3780),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3698),
.Y(n_3834)
);

AOI33xp33_ASAP7_75t_L g3835 ( 
.A1(n_3735),
.A2(n_3687),
.A3(n_3684),
.B1(n_3649),
.B2(n_3673),
.B3(n_3623),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3781),
.Y(n_3836)
);

OAI33xp33_ASAP7_75t_L g3837 ( 
.A1(n_3710),
.A2(n_3623),
.A3(n_3674),
.B1(n_3627),
.B2(n_3614),
.B3(n_3606),
.Y(n_3837)
);

OAI222xp33_ASAP7_75t_L g3838 ( 
.A1(n_3759),
.A2(n_3681),
.B1(n_3627),
.B2(n_3614),
.C1(n_3606),
.C2(n_3674),
.Y(n_3838)
);

OAI31xp33_ASAP7_75t_SL g3839 ( 
.A1(n_3746),
.A2(n_3681),
.A3(n_3606),
.B(n_3674),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3744),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3741),
.Y(n_3841)
);

XNOR2xp5_ASAP7_75t_L g3842 ( 
.A(n_3712),
.B(n_147),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3702),
.B(n_149),
.Y(n_3843)
);

OR2x2_ASAP7_75t_L g3844 ( 
.A(n_3726),
.B(n_150),
.Y(n_3844)
);

OAI33xp33_ASAP7_75t_L g3845 ( 
.A1(n_3723),
.A2(n_150),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.B3(n_154),
.Y(n_3845)
);

NAND3xp33_ASAP7_75t_SL g3846 ( 
.A(n_3715),
.B(n_151),
.C(n_153),
.Y(n_3846)
);

INVx1_ASAP7_75t_SL g3847 ( 
.A(n_3725),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3741),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3740),
.Y(n_3849)
);

INVx1_ASAP7_75t_SL g3850 ( 
.A(n_3731),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3718),
.B(n_155),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3719),
.B(n_155),
.Y(n_3852)
);

HB1xp67_ASAP7_75t_L g3853 ( 
.A(n_3727),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3755),
.B(n_3708),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3703),
.B(n_156),
.Y(n_3855)
);

NAND3xp33_ASAP7_75t_L g3856 ( 
.A(n_3722),
.B(n_157),
.C(n_158),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3707),
.B(n_157),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3742),
.Y(n_3858)
);

INVx1_ASAP7_75t_SL g3859 ( 
.A(n_3729),
.Y(n_3859)
);

OAI33xp33_ASAP7_75t_L g3860 ( 
.A1(n_3742),
.A2(n_3749),
.A3(n_3754),
.B1(n_3748),
.B2(n_3768),
.B3(n_3767),
.Y(n_3860)
);

NOR2x1_ASAP7_75t_L g3861 ( 
.A(n_3763),
.B(n_158),
.Y(n_3861)
);

OAI211xp5_ASAP7_75t_SL g3862 ( 
.A1(n_3739),
.A2(n_159),
.B(n_160),
.C(n_161),
.Y(n_3862)
);

AOI221x1_ASAP7_75t_L g3863 ( 
.A1(n_3768),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.C(n_163),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3711),
.B(n_162),
.Y(n_3864)
);

INVx5_ASAP7_75t_L g3865 ( 
.A(n_3740),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3736),
.B(n_164),
.Y(n_3866)
);

BUFx2_ASAP7_75t_L g3867 ( 
.A(n_3765),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3767),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3766),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3738),
.B(n_164),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3737),
.Y(n_3871)
);

BUFx3_ASAP7_75t_L g3872 ( 
.A(n_3765),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3743),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3805),
.B(n_3752),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3782),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3792),
.B(n_3764),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3809),
.B(n_3745),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3811),
.B(n_3777),
.Y(n_3878)
);

AOI32xp33_ASAP7_75t_L g3879 ( 
.A1(n_3862),
.A2(n_3769),
.A3(n_3750),
.B1(n_3771),
.B2(n_3751),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3805),
.B(n_3762),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3865),
.Y(n_3881)
);

OAI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3840),
.A2(n_3750),
.B1(n_3775),
.B2(n_3773),
.Y(n_3882)
);

OR2x2_ASAP7_75t_L g3883 ( 
.A(n_3792),
.B(n_3761),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3782),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3824),
.B(n_3811),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3865),
.Y(n_3886)
);

INVx2_ASAP7_75t_SL g3887 ( 
.A(n_3865),
.Y(n_3887)
);

AOI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_3846),
.A2(n_165),
.B1(n_170),
.B2(n_171),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3867),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3825),
.B(n_165),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3810),
.B(n_170),
.Y(n_3891)
);

AOI32xp33_ASAP7_75t_L g3892 ( 
.A1(n_3847),
.A2(n_171),
.A3(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3790),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3810),
.B(n_172),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3865),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3790),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3872),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3807),
.Y(n_3898)
);

INVxp67_ASAP7_75t_SL g3899 ( 
.A(n_3853),
.Y(n_3899)
);

NOR2x1_ASAP7_75t_L g3900 ( 
.A(n_3796),
.B(n_174),
.Y(n_3900)
);

XOR2x2_ASAP7_75t_L g3901 ( 
.A(n_3842),
.B(n_175),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3872),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3844),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3829),
.A2(n_175),
.B(n_176),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3812),
.B(n_176),
.Y(n_3905)
);

NAND2x2_ASAP7_75t_L g3906 ( 
.A(n_3833),
.B(n_177),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3804),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3797),
.B(n_177),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3783),
.B(n_178),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3807),
.Y(n_3910)
);

INVxp67_ASAP7_75t_L g3911 ( 
.A(n_3806),
.Y(n_3911)
);

OR2x2_ASAP7_75t_L g3912 ( 
.A(n_3816),
.B(n_178),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3796),
.Y(n_3913)
);

INVx1_ASAP7_75t_SL g3914 ( 
.A(n_3853),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3866),
.Y(n_3915)
);

NAND2x1p5_ASAP7_75t_L g3916 ( 
.A(n_3796),
.B(n_179),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3836),
.Y(n_3917)
);

OAI322xp33_ASAP7_75t_L g3918 ( 
.A1(n_3786),
.A2(n_180),
.A3(n_181),
.B1(n_182),
.B2(n_184),
.C1(n_185),
.C2(n_186),
.Y(n_3918)
);

NAND3xp33_ASAP7_75t_L g3919 ( 
.A(n_3851),
.B(n_181),
.C(n_182),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3855),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3803),
.B(n_186),
.Y(n_3921)
);

AND2x4_ASAP7_75t_L g3922 ( 
.A(n_3849),
.B(n_187),
.Y(n_3922)
);

OR2x2_ASAP7_75t_L g3923 ( 
.A(n_3816),
.B(n_187),
.Y(n_3923)
);

AOI32xp33_ASAP7_75t_L g3924 ( 
.A1(n_3803),
.A2(n_188),
.A3(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3864),
.Y(n_3925)
);

OA21x2_ASAP7_75t_L g3926 ( 
.A1(n_3838),
.A2(n_188),
.B(n_189),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3859),
.B(n_192),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3791),
.B(n_192),
.Y(n_3928)
);

XOR2x2_ASAP7_75t_L g3929 ( 
.A(n_3806),
.B(n_193),
.Y(n_3929)
);

NAND3xp33_ASAP7_75t_L g3930 ( 
.A(n_3791),
.B(n_193),
.C(n_194),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3831),
.Y(n_3931)
);

NAND5xp2_ASAP7_75t_L g3932 ( 
.A(n_3818),
.B(n_195),
.C(n_196),
.D(n_198),
.E(n_199),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3832),
.B(n_195),
.Y(n_3933)
);

OAI311xp33_ASAP7_75t_L g3934 ( 
.A1(n_3814),
.A2(n_196),
.A3(n_200),
.B1(n_201),
.C1(n_202),
.Y(n_3934)
);

HB1xp67_ASAP7_75t_L g3935 ( 
.A(n_3831),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3830),
.B(n_201),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3817),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3799),
.B(n_3832),
.Y(n_3938)
);

NAND4xp75_ASAP7_75t_L g3939 ( 
.A(n_3789),
.B(n_202),
.C(n_203),
.D(n_204),
.Y(n_3939)
);

OAI322xp33_ASAP7_75t_L g3940 ( 
.A1(n_3784),
.A2(n_203),
.A3(n_205),
.B1(n_207),
.B2(n_208),
.C1(n_209),
.C2(n_210),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3833),
.B(n_207),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3785),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3850),
.B(n_209),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3787),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3860),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_3945)
);

AOI211xp5_ASAP7_75t_L g3946 ( 
.A1(n_3819),
.A2(n_211),
.B(n_212),
.C(n_214),
.Y(n_3946)
);

OR2x2_ASAP7_75t_L g3947 ( 
.A(n_3827),
.B(n_215),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3788),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3857),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3831),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3849),
.Y(n_3951)
);

AND2x4_ASAP7_75t_L g3952 ( 
.A(n_3822),
.B(n_215),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3822),
.B(n_216),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3852),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3784),
.B(n_218),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3823),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3828),
.B(n_218),
.Y(n_3957)
);

INVx2_ASAP7_75t_SL g3958 ( 
.A(n_3823),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3794),
.Y(n_3959)
);

CKINVDCx16_ASAP7_75t_R g3960 ( 
.A(n_3843),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3870),
.Y(n_3961)
);

OR2x2_ASAP7_75t_L g3962 ( 
.A(n_3854),
.B(n_219),
.Y(n_3962)
);

INVx3_ASAP7_75t_L g3963 ( 
.A(n_3794),
.Y(n_3963)
);

AOI33xp33_ASAP7_75t_L g3964 ( 
.A1(n_3945),
.A2(n_3814),
.A3(n_3808),
.B1(n_3828),
.B2(n_3840),
.B3(n_3869),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3935),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3952),
.Y(n_3966)
);

INVxp67_ASAP7_75t_L g3967 ( 
.A(n_3900),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3885),
.B(n_3815),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3898),
.B(n_3815),
.Y(n_3969)
);

OR2x2_ASAP7_75t_L g3970 ( 
.A(n_3960),
.B(n_3871),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3931),
.Y(n_3971)
);

NAND3xp33_ASAP7_75t_L g3972 ( 
.A(n_3946),
.B(n_3839),
.C(n_3835),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3910),
.B(n_3861),
.Y(n_3973)
);

NAND3xp33_ASAP7_75t_SL g3974 ( 
.A(n_3946),
.B(n_3793),
.C(n_3856),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3950),
.Y(n_3975)
);

HB1xp67_ASAP7_75t_L g3976 ( 
.A(n_3887),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3939),
.A2(n_3800),
.B1(n_3845),
.B2(n_3808),
.Y(n_3977)
);

OR2x2_ASAP7_75t_L g3978 ( 
.A(n_3938),
.B(n_3873),
.Y(n_3978)
);

OR2x2_ASAP7_75t_L g3979 ( 
.A(n_3937),
.B(n_3795),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3890),
.B(n_3877),
.Y(n_3980)
);

OR2x2_ASAP7_75t_L g3981 ( 
.A(n_3889),
.B(n_3798),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3941),
.Y(n_3982)
);

INVx2_ASAP7_75t_SL g3983 ( 
.A(n_3952),
.Y(n_3983)
);

BUFx2_ASAP7_75t_L g3984 ( 
.A(n_3908),
.Y(n_3984)
);

NOR2xp33_ASAP7_75t_R g3985 ( 
.A(n_3897),
.B(n_3902),
.Y(n_3985)
);

BUFx2_ASAP7_75t_L g3986 ( 
.A(n_3908),
.Y(n_3986)
);

AOI222xp33_ASAP7_75t_L g3987 ( 
.A1(n_3914),
.A2(n_3801),
.B1(n_3834),
.B2(n_3826),
.C1(n_3837),
.C2(n_3813),
.Y(n_3987)
);

NOR3xp33_ASAP7_75t_L g3988 ( 
.A(n_3904),
.B(n_3820),
.C(n_3802),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3914),
.B(n_3821),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3881),
.Y(n_3990)
);

AND2x4_ASAP7_75t_SL g3991 ( 
.A(n_3936),
.B(n_3841),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3893),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3896),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3875),
.Y(n_3994)
);

INVx1_ASAP7_75t_SL g3995 ( 
.A(n_3953),
.Y(n_3995)
);

OAI221xp5_ASAP7_75t_L g3996 ( 
.A1(n_3879),
.A2(n_3858),
.B1(n_3848),
.B2(n_3868),
.C(n_3835),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3958),
.B(n_3863),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3951),
.B(n_220),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3916),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3899),
.B(n_220),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3957),
.B(n_222),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3911),
.B(n_223),
.Y(n_4002)
);

AND2x4_ASAP7_75t_L g4003 ( 
.A(n_3913),
.B(n_224),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3884),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3891),
.Y(n_4005)
);

AND2x4_ASAP7_75t_L g4006 ( 
.A(n_3886),
.B(n_225),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3915),
.B(n_225),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3883),
.B(n_226),
.Y(n_4008)
);

NOR2xp67_ASAP7_75t_SL g4009 ( 
.A(n_3905),
.B(n_226),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3895),
.Y(n_4010)
);

HB1xp67_ASAP7_75t_L g4011 ( 
.A(n_3963),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3894),
.Y(n_4012)
);

AND2x2_ASAP7_75t_SL g4013 ( 
.A(n_3907),
.B(n_227),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3927),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3925),
.B(n_228),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3912),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3957),
.B(n_228),
.Y(n_4017)
);

NOR2xp33_ASAP7_75t_L g4018 ( 
.A(n_3949),
.B(n_229),
.Y(n_4018)
);

NOR3xp33_ASAP7_75t_L g4019 ( 
.A(n_3961),
.B(n_229),
.C(n_230),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3923),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3963),
.Y(n_4021)
);

OAI21xp5_ASAP7_75t_SL g4022 ( 
.A1(n_3888),
.A2(n_230),
.B(n_231),
.Y(n_4022)
);

NOR3xp33_ASAP7_75t_SL g4023 ( 
.A(n_3934),
.B(n_231),
.C(n_232),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_3882),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3876),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3933),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3880),
.B(n_236),
.Y(n_4027)
);

OR2x4_ASAP7_75t_L g4028 ( 
.A(n_3920),
.B(n_237),
.Y(n_4028)
);

INVx1_ASAP7_75t_SL g4029 ( 
.A(n_3926),
.Y(n_4029)
);

OR2x2_ASAP7_75t_L g4030 ( 
.A(n_3880),
.B(n_238),
.Y(n_4030)
);

HB1xp67_ASAP7_75t_L g4031 ( 
.A(n_3956),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3954),
.B(n_241),
.Y(n_4032)
);

CKINVDCx5p33_ASAP7_75t_R g4033 ( 
.A(n_3929),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3874),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3930),
.B(n_242),
.Y(n_4035)
);

AND2x2_ASAP7_75t_SL g4036 ( 
.A(n_3962),
.B(n_242),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3922),
.Y(n_4037)
);

OR2x2_ASAP7_75t_L g4038 ( 
.A(n_3943),
.B(n_244),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3903),
.B(n_244),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3878),
.B(n_245),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3959),
.B(n_245),
.Y(n_4041)
);

OAI321xp33_ASAP7_75t_L g4042 ( 
.A1(n_3882),
.A2(n_246),
.A3(n_247),
.B1(n_248),
.B2(n_249),
.C(n_250),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3874),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3930),
.B(n_247),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3917),
.B(n_248),
.Y(n_4045)
);

OAI221xp5_ASAP7_75t_L g4046 ( 
.A1(n_3888),
.A2(n_3892),
.B1(n_3924),
.B2(n_3921),
.C(n_3919),
.Y(n_4046)
);

OAI31xp33_ASAP7_75t_L g4047 ( 
.A1(n_3934),
.A2(n_251),
.A3(n_252),
.B(n_253),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3984),
.B(n_3942),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3968),
.B(n_3909),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_4011),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3986),
.B(n_3944),
.Y(n_4051)
);

AND2x4_ASAP7_75t_L g4052 ( 
.A(n_3966),
.B(n_3948),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3966),
.B(n_3901),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3983),
.B(n_4029),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3990),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3970),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_4031),
.Y(n_4057)
);

NOR4xp25_ASAP7_75t_L g4058 ( 
.A(n_4029),
.B(n_3918),
.C(n_3919),
.D(n_3928),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3968),
.B(n_3922),
.Y(n_4059)
);

OR2x2_ASAP7_75t_L g4060 ( 
.A(n_3995),
.B(n_3947),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_4037),
.B(n_3955),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3976),
.Y(n_4062)
);

NOR2xp33_ASAP7_75t_L g4063 ( 
.A(n_3967),
.B(n_3932),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3965),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3997),
.B(n_3926),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3980),
.B(n_3906),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4021),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4006),
.Y(n_4068)
);

OAI31xp33_ASAP7_75t_L g4069 ( 
.A1(n_3972),
.A2(n_3932),
.A3(n_3918),
.B(n_3940),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3969),
.B(n_3940),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4006),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3997),
.B(n_251),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_4047),
.B(n_253),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_4010),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_3995),
.B(n_254),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_4047),
.B(n_254),
.Y(n_4076)
);

HB1xp67_ASAP7_75t_L g4077 ( 
.A(n_4028),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4003),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3973),
.B(n_3999),
.Y(n_4079)
);

CKINVDCx16_ASAP7_75t_R g4080 ( 
.A(n_3985),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4003),
.Y(n_4081)
);

INVx1_ASAP7_75t_SL g4082 ( 
.A(n_4013),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3998),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3991),
.B(n_255),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4028),
.Y(n_4085)
);

HB1xp67_ASAP7_75t_L g4086 ( 
.A(n_4000),
.Y(n_4086)
);

AND2x4_ASAP7_75t_L g4087 ( 
.A(n_4025),
.B(n_255),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3978),
.B(n_256),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_4040),
.B(n_3982),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4033),
.B(n_256),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4008),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4039),
.Y(n_4092)
);

HB1xp67_ASAP7_75t_L g4093 ( 
.A(n_4000),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_3981),
.B(n_257),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3971),
.B(n_258),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4007),
.Y(n_4096)
);

O2A1O1Ixp33_ASAP7_75t_L g4097 ( 
.A1(n_4042),
.A2(n_259),
.B(n_261),
.C(n_262),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4036),
.B(n_259),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3964),
.B(n_4023),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4032),
.Y(n_4100)
);

AND2x2_ASAP7_75t_L g4101 ( 
.A(n_3975),
.B(n_261),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4041),
.Y(n_4102)
);

NOR2xp33_ASAP7_75t_L g4103 ( 
.A(n_4046),
.B(n_263),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_3979),
.B(n_4027),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4002),
.Y(n_4105)
);

NAND4xp75_ASAP7_75t_L g4106 ( 
.A(n_3989),
.B(n_264),
.C(n_265),
.D(n_266),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4045),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_4038),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_4030),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3989),
.Y(n_4110)
);

NOR2xp67_ASAP7_75t_L g4111 ( 
.A(n_4042),
.B(n_4014),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4009),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_4035),
.Y(n_4113)
);

CKINVDCx16_ASAP7_75t_R g4114 ( 
.A(n_3974),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4080),
.B(n_3977),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_4054),
.Y(n_4116)
);

NAND2x1_ASAP7_75t_L g4117 ( 
.A(n_4052),
.B(n_3994),
.Y(n_4117)
);

NOR2xp33_ASAP7_75t_L g4118 ( 
.A(n_4076),
.B(n_4046),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_4076),
.A2(n_3972),
.B(n_4024),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_4114),
.A2(n_3996),
.B1(n_4044),
.B2(n_4035),
.Y(n_4120)
);

INVx3_ASAP7_75t_L g4121 ( 
.A(n_4052),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4077),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_4065),
.A2(n_3987),
.B(n_4044),
.Y(n_4123)
);

OAI21xp33_ASAP7_75t_L g4124 ( 
.A1(n_4063),
.A2(n_3987),
.B(n_4034),
.Y(n_4124)
);

AOI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_4073),
.A2(n_4001),
.B(n_4017),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_4059),
.B(n_4022),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_4082),
.B(n_4022),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_4052),
.Y(n_4128)
);

OAI32xp33_ASAP7_75t_L g4129 ( 
.A1(n_4099),
.A2(n_3988),
.A3(n_4043),
.B1(n_4004),
.B2(n_3992),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_4069),
.A2(n_4072),
.B(n_4097),
.Y(n_4130)
);

AOI32xp33_ASAP7_75t_L g4131 ( 
.A1(n_4063),
.A2(n_4019),
.A3(n_4001),
.B1(n_4017),
.B2(n_3993),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4077),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_4070),
.B(n_4016),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4048),
.Y(n_4134)
);

AOI22x1_ASAP7_75t_L g4135 ( 
.A1(n_4049),
.A2(n_4020),
.B1(n_4012),
.B2(n_4005),
.Y(n_4135)
);

BUFx2_ASAP7_75t_L g4136 ( 
.A(n_4048),
.Y(n_4136)
);

AO32x1_ASAP7_75t_L g4137 ( 
.A1(n_4062),
.A2(n_4026),
.A3(n_4018),
.B1(n_4015),
.B2(n_267),
.Y(n_4137)
);

OAI221xp5_ASAP7_75t_SL g4138 ( 
.A1(n_4058),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4066),
.B(n_270),
.Y(n_4139)
);

AOI321xp33_ASAP7_75t_L g4140 ( 
.A1(n_4056),
.A2(n_272),
.A3(n_273),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_4051),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4051),
.B(n_272),
.Y(n_4142)
);

AND2x4_ASAP7_75t_L g4143 ( 
.A(n_4084),
.B(n_273),
.Y(n_4143)
);

AOI21xp33_ASAP7_75t_L g4144 ( 
.A1(n_4060),
.A2(n_274),
.B(n_278),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4068),
.Y(n_4145)
);

OAI31xp33_ASAP7_75t_L g4146 ( 
.A1(n_4103),
.A2(n_278),
.A3(n_279),
.B(n_280),
.Y(n_4146)
);

BUFx3_ASAP7_75t_L g4147 ( 
.A(n_4071),
.Y(n_4147)
);

AOI32xp33_ASAP7_75t_L g4148 ( 
.A1(n_4103),
.A2(n_279),
.A3(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_4053),
.B(n_4078),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_4081),
.B(n_283),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_4084),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4075),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4089),
.Y(n_4153)
);

NAND2xp33_ASAP7_75t_R g4154 ( 
.A(n_4089),
.B(n_283),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4087),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4085),
.B(n_285),
.Y(n_4156)
);

AOI221xp5_ASAP7_75t_L g4157 ( 
.A1(n_4110),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.C(n_288),
.Y(n_4157)
);

OAI22x1_ASAP7_75t_L g4158 ( 
.A1(n_4112),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_4158)
);

OAI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_4111),
.A2(n_292),
.B(n_293),
.Y(n_4159)
);

NAND2x1p5_ASAP7_75t_L g4160 ( 
.A(n_4091),
.B(n_292),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4057),
.B(n_294),
.Y(n_4161)
);

AOI32xp33_ASAP7_75t_L g4162 ( 
.A1(n_4055),
.A2(n_294),
.A3(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4061),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4061),
.Y(n_4164)
);

AOI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_4079),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4050),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4079),
.B(n_300),
.Y(n_4167)
);

OAI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_4064),
.A2(n_301),
.B(n_302),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4092),
.B(n_305),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4096),
.A2(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_4170)
);

INVxp67_ASAP7_75t_L g4171 ( 
.A(n_4086),
.Y(n_4171)
);

OAI211xp5_ASAP7_75t_L g4172 ( 
.A1(n_4074),
.A2(n_4067),
.B(n_4086),
.C(n_4093),
.Y(n_4172)
);

AOI221xp5_ASAP7_75t_L g4173 ( 
.A1(n_4113),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4087),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_4100),
.B(n_309),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4088),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4095),
.Y(n_4177)
);

OAI21xp5_ASAP7_75t_SL g4178 ( 
.A1(n_4083),
.A2(n_310),
.B(n_313),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4087),
.B(n_4095),
.Y(n_4179)
);

INVx1_ASAP7_75t_SL g4180 ( 
.A(n_4136),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4121),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4128),
.B(n_4101),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4123),
.A2(n_4090),
.B1(n_4104),
.B2(n_4107),
.Y(n_4183)
);

OR2x2_ASAP7_75t_L g4184 ( 
.A(n_4121),
.B(n_4109),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4134),
.B(n_4101),
.Y(n_4185)
);

AOI211xp5_ASAP7_75t_SL g4186 ( 
.A1(n_4124),
.A2(n_4093),
.B(n_4094),
.C(n_4105),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4117),
.Y(n_4187)
);

INVxp67_ASAP7_75t_L g4188 ( 
.A(n_4154),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4179),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4155),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4174),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_4141),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4153),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4147),
.B(n_4102),
.Y(n_4194)
);

XNOR2x2_ASAP7_75t_L g4195 ( 
.A(n_4118),
.B(n_4106),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4126),
.Y(n_4196)
);

OAI211xp5_ASAP7_75t_L g4197 ( 
.A1(n_4119),
.A2(n_4113),
.B(n_4109),
.C(n_4108),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4160),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4151),
.Y(n_4199)
);

XNOR2x2_ASAP7_75t_L g4200 ( 
.A(n_4120),
.B(n_4098),
.Y(n_4200)
);

AO22x1_ASAP7_75t_L g4201 ( 
.A1(n_4163),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_4138),
.B(n_4177),
.Y(n_4202)
);

NAND2x1_ASAP7_75t_L g4203 ( 
.A(n_4164),
.B(n_314),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4139),
.B(n_315),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4122),
.B(n_317),
.Y(n_4205)
);

INVx2_ASAP7_75t_SL g4206 ( 
.A(n_4143),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_4132),
.B(n_317),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4143),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4159),
.B(n_318),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4152),
.B(n_318),
.Y(n_4210)
);

NAND4xp25_ASAP7_75t_L g4211 ( 
.A(n_4130),
.B(n_4115),
.C(n_4127),
.D(n_4133),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4142),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_L g4213 ( 
.A(n_4116),
.B(n_319),
.Y(n_4213)
);

INVx1_ASAP7_75t_SL g4214 ( 
.A(n_4158),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4145),
.B(n_319),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4148),
.B(n_4162),
.Y(n_4216)
);

XNOR2xp5_ASAP7_75t_L g4217 ( 
.A(n_4135),
.B(n_320),
.Y(n_4217)
);

INVxp67_ASAP7_75t_L g4218 ( 
.A(n_4167),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_4148),
.B(n_322),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4149),
.Y(n_4220)
);

AOI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_4137),
.A2(n_322),
.B(n_324),
.Y(n_4221)
);

AOI221xp5_ASAP7_75t_L g4222 ( 
.A1(n_4129),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_4222)
);

INVx1_ASAP7_75t_SL g4223 ( 
.A(n_4169),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4175),
.B(n_325),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4162),
.B(n_326),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4150),
.Y(n_4226)
);

CKINVDCx16_ASAP7_75t_R g4227 ( 
.A(n_4176),
.Y(n_4227)
);

NAND3xp33_ASAP7_75t_SL g4228 ( 
.A(n_4131),
.B(n_327),
.C(n_328),
.Y(n_4228)
);

AOI211xp5_ASAP7_75t_L g4229 ( 
.A1(n_4172),
.A2(n_329),
.B(n_330),
.C(n_331),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4156),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4166),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4171),
.B(n_329),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_4125),
.B(n_330),
.Y(n_4233)
);

OR2x2_ASAP7_75t_L g4234 ( 
.A(n_4161),
.B(n_4178),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4184),
.Y(n_4235)
);

O2A1O1Ixp5_ASAP7_75t_L g4236 ( 
.A1(n_4187),
.A2(n_4144),
.B(n_4168),
.C(n_4137),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_4206),
.Y(n_4237)
);

INVx2_ASAP7_75t_SL g4238 ( 
.A(n_4203),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4181),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_L g4240 ( 
.A(n_4180),
.B(n_4165),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4182),
.Y(n_4241)
);

OAI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_4221),
.A2(n_4146),
.B(n_4157),
.Y(n_4242)
);

INVxp67_ASAP7_75t_L g4243 ( 
.A(n_4202),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4208),
.Y(n_4244)
);

OAI211xp5_ASAP7_75t_SL g4245 ( 
.A1(n_4186),
.A2(n_4131),
.B(n_4188),
.C(n_4197),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_4180),
.B(n_4170),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4190),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4192),
.B(n_4173),
.Y(n_4248)
);

OAI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_4217),
.A2(n_4137),
.B(n_4140),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4192),
.B(n_331),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4194),
.B(n_332),
.Y(n_4251)
);

INVxp67_ASAP7_75t_SL g4252 ( 
.A(n_4185),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4191),
.Y(n_4253)
);

INVxp67_ASAP7_75t_SL g4254 ( 
.A(n_4195),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_4227),
.B(n_333),
.Y(n_4255)
);

AND3x2_ASAP7_75t_L g4256 ( 
.A(n_4229),
.B(n_334),
.C(n_335),
.Y(n_4256)
);

AOI21xp33_ASAP7_75t_L g4257 ( 
.A1(n_4198),
.A2(n_336),
.B(n_337),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4204),
.Y(n_4258)
);

NAND2xp33_ASAP7_75t_R g4259 ( 
.A(n_4220),
.B(n_337),
.Y(n_4259)
);

INVxp33_ASAP7_75t_L g4260 ( 
.A(n_4216),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_4201),
.B(n_338),
.Y(n_4261)
);

XOR2x2_ASAP7_75t_L g4262 ( 
.A(n_4200),
.B(n_338),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4224),
.Y(n_4263)
);

OR2x2_ASAP7_75t_L g4264 ( 
.A(n_4214),
.B(n_4228),
.Y(n_4264)
);

AOI32xp33_ASAP7_75t_L g4265 ( 
.A1(n_4214),
.A2(n_339),
.A3(n_340),
.B1(n_341),
.B2(n_344),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4215),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_4223),
.B(n_339),
.Y(n_4267)
);

NAND2x1p5_ASAP7_75t_L g4268 ( 
.A(n_4223),
.B(n_4210),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4199),
.Y(n_4269)
);

CKINVDCx14_ASAP7_75t_R g4270 ( 
.A(n_4183),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4209),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4186),
.B(n_340),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_4211),
.B(n_459),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4193),
.B(n_461),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4234),
.Y(n_4275)
);

OAI222xp33_ASAP7_75t_L g4276 ( 
.A1(n_4254),
.A2(n_4189),
.B1(n_4196),
.B2(n_4231),
.C1(n_4218),
.C2(n_4212),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4238),
.B(n_4222),
.Y(n_4277)
);

NOR3xp33_ASAP7_75t_L g4278 ( 
.A(n_4245),
.B(n_4211),
.C(n_4233),
.Y(n_4278)
);

AOI21xp5_ASAP7_75t_L g4279 ( 
.A1(n_4272),
.A2(n_4225),
.B(n_4219),
.Y(n_4279)
);

AOI22xp5_ASAP7_75t_L g4280 ( 
.A1(n_4270),
.A2(n_4230),
.B1(n_4213),
.B2(n_4226),
.Y(n_4280)
);

OAI22xp5_ASAP7_75t_L g4281 ( 
.A1(n_4243),
.A2(n_4207),
.B1(n_4205),
.B2(n_4232),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_L g4282 ( 
.A(n_4260),
.B(n_462),
.Y(n_4282)
);

AOI211x1_ASAP7_75t_L g4283 ( 
.A1(n_4249),
.A2(n_2895),
.B(n_1266),
.C(n_1254),
.Y(n_4283)
);

NOR2x1_ASAP7_75t_L g4284 ( 
.A(n_4264),
.B(n_955),
.Y(n_4284)
);

AOI21xp5_ASAP7_75t_L g4285 ( 
.A1(n_4255),
.A2(n_955),
.B(n_948),
.Y(n_4285)
);

AO22x2_ASAP7_75t_L g4286 ( 
.A1(n_4244),
.A2(n_1266),
.B1(n_1254),
.B2(n_1182),
.Y(n_4286)
);

AOI21xp5_ASAP7_75t_L g4287 ( 
.A1(n_4249),
.A2(n_955),
.B(n_948),
.Y(n_4287)
);

AO22x2_ASAP7_75t_L g4288 ( 
.A1(n_4235),
.A2(n_1266),
.B1(n_1254),
.B2(n_1182),
.Y(n_4288)
);

NOR3xp33_ASAP7_75t_L g4289 ( 
.A(n_4236),
.B(n_4275),
.C(n_4252),
.Y(n_4289)
);

NAND4xp75_ASAP7_75t_L g4290 ( 
.A(n_4240),
.B(n_955),
.C(n_948),
.D(n_943),
.Y(n_4290)
);

OA22x2_ASAP7_75t_L g4291 ( 
.A1(n_4256),
.A2(n_955),
.B1(n_948),
.B2(n_1266),
.Y(n_4291)
);

NOR3xp33_ASAP7_75t_L g4292 ( 
.A(n_4241),
.B(n_1167),
.C(n_1236),
.Y(n_4292)
);

XNOR2x1_ASAP7_75t_SL g4293 ( 
.A(n_4268),
.B(n_1266),
.Y(n_4293)
);

AOI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_4237),
.A2(n_948),
.B1(n_1254),
.B2(n_1237),
.Y(n_4294)
);

NOR3xp33_ASAP7_75t_L g4295 ( 
.A(n_4258),
.B(n_1254),
.C(n_1237),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4251),
.B(n_1237),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4268),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_4246),
.B(n_1237),
.Y(n_4298)
);

NOR3x1_ASAP7_75t_L g4299 ( 
.A(n_4242),
.B(n_1237),
.C(n_1232),
.Y(n_4299)
);

OAI211xp5_ASAP7_75t_SL g4300 ( 
.A1(n_4242),
.A2(n_1232),
.B(n_1207),
.C(n_930),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4297),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4277),
.Y(n_4302)
);

NOR3xp33_ASAP7_75t_L g4303 ( 
.A(n_4276),
.B(n_4289),
.C(n_4281),
.Y(n_4303)
);

OAI21xp33_ASAP7_75t_SL g4304 ( 
.A1(n_4293),
.A2(n_4248),
.B(n_4239),
.Y(n_4304)
);

OAI211xp5_ASAP7_75t_L g4305 ( 
.A1(n_4280),
.A2(n_4265),
.B(n_4250),
.C(n_4253),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4296),
.Y(n_4306)
);

AOI221xp5_ASAP7_75t_L g4307 ( 
.A1(n_4278),
.A2(n_4273),
.B1(n_4247),
.B2(n_4269),
.C(n_4246),
.Y(n_4307)
);

XNOR2xp5_ASAP7_75t_L g4308 ( 
.A(n_4279),
.B(n_4262),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4291),
.Y(n_4309)
);

AOI221x1_ASAP7_75t_L g4310 ( 
.A1(n_4282),
.A2(n_4263),
.B1(n_4266),
.B2(n_4271),
.C(n_4257),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4299),
.B(n_4261),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4284),
.B(n_4267),
.Y(n_4312)
);

AOI22xp5_ASAP7_75t_L g4313 ( 
.A1(n_4292),
.A2(n_4259),
.B1(n_4274),
.B2(n_4295),
.Y(n_4313)
);

HB1xp67_ASAP7_75t_L g4314 ( 
.A(n_4298),
.Y(n_4314)
);

NOR3xp33_ASAP7_75t_L g4315 ( 
.A(n_4300),
.B(n_1232),
.C(n_1207),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4288),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4301),
.B(n_4287),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_4302),
.Y(n_4318)
);

OA22x2_ASAP7_75t_L g4319 ( 
.A1(n_4308),
.A2(n_4310),
.B1(n_4305),
.B2(n_4313),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4311),
.Y(n_4320)
);

AO22x2_ASAP7_75t_L g4321 ( 
.A1(n_4303),
.A2(n_4290),
.B1(n_4283),
.B2(n_4285),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4312),
.Y(n_4322)
);

NOR2x1_ASAP7_75t_L g4323 ( 
.A(n_4316),
.B(n_4309),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4314),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4304),
.Y(n_4325)
);

OAI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4307),
.A2(n_4294),
.B1(n_4286),
.B2(n_1232),
.Y(n_4326)
);

AOI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4306),
.A2(n_4286),
.B1(n_1232),
.B2(n_1207),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4325),
.B(n_4315),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_4319),
.A2(n_4324),
.B(n_4318),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4323),
.B(n_1207),
.Y(n_4330)
);

OAI221xp5_ASAP7_75t_SL g4331 ( 
.A1(n_4320),
.A2(n_930),
.B1(n_942),
.B2(n_963),
.C(n_979),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4322),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4321),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4317),
.Y(n_4334)
);

OAI22xp5_ASAP7_75t_L g4335 ( 
.A1(n_4332),
.A2(n_4327),
.B1(n_4326),
.B2(n_930),
.Y(n_4335)
);

XOR2xp5_ASAP7_75t_L g4336 ( 
.A(n_4329),
.B(n_930),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4330),
.Y(n_4337)
);

INVx3_ASAP7_75t_L g4338 ( 
.A(n_4333),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4328),
.B(n_930),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4338),
.A2(n_4334),
.B(n_4331),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4336),
.A2(n_4335),
.B(n_4339),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4340),
.Y(n_4342)
);

AND2x4_ASAP7_75t_L g4343 ( 
.A(n_4341),
.B(n_4337),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4343),
.Y(n_4344)
);

NAND4xp75_ASAP7_75t_L g4345 ( 
.A(n_4344),
.B(n_4342),
.C(n_942),
.D(n_930),
.Y(n_4345)
);

OR3x1_ASAP7_75t_L g4346 ( 
.A(n_4345),
.B(n_942),
.C(n_963),
.Y(n_4346)
);

OAI21xp5_ASAP7_75t_SL g4347 ( 
.A1(n_4346),
.A2(n_942),
.B(n_963),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4347),
.Y(n_4348)
);

OAI22x1_ASAP7_75t_L g4349 ( 
.A1(n_4348),
.A2(n_942),
.B1(n_963),
.B2(n_979),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4349),
.Y(n_4350)
);

INVxp67_ASAP7_75t_SL g4351 ( 
.A(n_4350),
.Y(n_4351)
);

HB1xp67_ASAP7_75t_L g4352 ( 
.A(n_4351),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_4352),
.A2(n_942),
.B(n_979),
.Y(n_4353)
);

AOI221xp5_ASAP7_75t_L g4354 ( 
.A1(n_4353),
.A2(n_979),
.B1(n_1060),
.B2(n_1061),
.C(n_4325),
.Y(n_4354)
);

AOI211xp5_ASAP7_75t_L g4355 ( 
.A1(n_4354),
.A2(n_979),
.B(n_1061),
.C(n_4332),
.Y(n_4355)
);


endmodule