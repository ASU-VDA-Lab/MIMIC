module fake_aes_1021_n_681 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_681);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g78 ( .A(n_68), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_70), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_11), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_77), .B(n_58), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_6), .Y(n_82) );
INVx3_ASAP7_75t_L g83 ( .A(n_39), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_20), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_41), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_38), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_9), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_26), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_3), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_SL g93 ( .A(n_30), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_55), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_33), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_63), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_21), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_24), .Y(n_100) );
XNOR2x2_ASAP7_75t_L g101 ( .A(n_12), .B(n_61), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_23), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_67), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_29), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_15), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_34), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_53), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_11), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_20), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_50), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_28), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_86), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_79), .B(n_0), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_120), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_124), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_78), .B(n_1), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_80), .B(n_1), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_91), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_108), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_84), .B(n_2), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_87), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_84), .B(n_3), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_89), .B(n_4), .Y(n_152) );
NAND3xp33_ASAP7_75t_L g153 ( .A(n_89), .B(n_37), .C(n_74), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_101), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_119), .A2(n_32), .B(n_73), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_101), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_92), .B(n_4), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_90), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_92), .Y(n_161) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_95), .A2(n_40), .B(n_71), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_113), .B(n_5), .Y(n_163) );
INVxp33_ASAP7_75t_SL g164 ( .A(n_102), .Y(n_164) );
BUFx8_ASAP7_75t_L g165 ( .A(n_81), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_115), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_129), .B(n_110), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_129), .B(n_122), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_132), .B(n_122), .Y(n_170) );
NAND3x1_ASAP7_75t_L g171 ( .A(n_132), .B(n_113), .C(n_116), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_132), .B(n_151), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_135), .B(n_105), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_135), .B(n_106), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_127), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_125), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_141), .B(n_116), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_141), .B(n_107), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVxp67_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_126), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_148), .B(n_103), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_126), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_165), .B(n_111), .C(n_118), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_130), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
BUFx4_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_157), .A2(n_118), .B1(n_117), .B2(n_114), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
OR2x6_ASAP7_75t_L g199 ( .A(n_137), .B(n_81), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_161), .B(n_117), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_128), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_164), .B(n_100), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_128), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_128), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_161), .B(n_114), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_144), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_148), .B(n_99), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_145), .B(n_104), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_127), .B(n_109), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_131), .B(n_111), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_146), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_131), .B(n_96), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
AO22x2_ASAP7_75t_L g225 ( .A1(n_154), .A2(n_96), .B1(n_95), .B2(n_94), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_172), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_204), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_200), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_186), .B(n_165), .C(n_149), .Y(n_230) );
BUFx12f_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_172), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_204), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_139), .B1(n_143), .B2(n_134), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_175), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_200), .B(n_166), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_212), .B(n_165), .Y(n_239) );
NOR3xp33_ASAP7_75t_SL g240 ( .A(n_203), .B(n_156), .C(n_147), .Y(n_240) );
NOR3xp33_ASAP7_75t_SL g241 ( .A(n_215), .B(n_163), .C(n_138), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_181), .A2(n_134), .B(n_139), .C(n_143), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_212), .B(n_163), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_207), .B(n_158), .Y(n_245) );
OR2x6_ASAP7_75t_L g246 ( .A(n_199), .B(n_152), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_212), .B(n_158), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_183), .B(n_147), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_167), .B(n_138), .C(n_152), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_170), .B(n_162), .Y(n_252) );
INVxp33_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_170), .B(n_150), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_179), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_168), .B(n_144), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_170), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_179), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_179), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_197), .A2(n_150), .B1(n_160), .B2(n_159), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_199), .A2(n_121), .B1(n_160), .B2(n_159), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_199), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_189), .B(n_153), .C(n_6), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_199), .B(n_162), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_192), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_183), .B(n_160), .Y(n_271) );
AOI211xp5_ASAP7_75t_L g272 ( .A1(n_168), .A2(n_153), .B(n_159), .C(n_162), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_184), .B(n_112), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_184), .B(n_93), .Y(n_274) );
NOR3xp33_ASAP7_75t_SL g275 ( .A(n_214), .B(n_5), .C(n_7), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_210), .B(n_211), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_187), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_220), .B(n_7), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_197), .A2(n_8), .B1(n_10), .B2(n_12), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_171), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_171), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_223), .B(n_16), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_223), .B(n_18), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_173), .B(n_18), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_188), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_244), .B(n_196), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_231), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_233), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_243), .A2(n_178), .B(n_225), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_252), .A2(n_191), .B(n_218), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_250), .B(n_225), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_259), .A2(n_225), .B1(n_198), .B2(n_205), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_259), .B(n_225), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_255), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_264), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_270), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_228), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_270), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_226), .B(n_202), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_232), .B(n_195), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_246), .A2(n_205), .B1(n_188), .B2(n_190), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_246), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_238), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_265), .A2(n_190), .B1(n_206), .B2(n_208), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_248), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_249), .B(n_206), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_265), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_229), .B(n_195), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_248), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_258), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
INVx3_ASAP7_75t_SL g327 ( .A(n_249), .Y(n_327) );
INVx3_ASAP7_75t_SL g328 ( .A(n_285), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_263), .A2(n_213), .B1(n_208), .B2(n_201), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_239), .A2(n_217), .B(n_216), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_227), .B(n_213), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_248), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_256), .Y(n_335) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_257), .B(n_217), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_268), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_295), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_297), .A2(n_235), .B1(n_285), .B2(n_262), .Y(n_340) );
BUFx4f_ASAP7_75t_L g341 ( .A(n_322), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_289), .Y(n_342) );
BUFx4_ASAP7_75t_SL g343 ( .A(n_322), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_297), .B(n_251), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_294), .A2(n_301), .B1(n_235), .B2(n_262), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_301), .A2(n_268), .B1(n_280), .B2(n_283), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_292), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_322), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_252), .B(n_272), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_293), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_293), .B(n_251), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_299), .Y(n_353) );
AOI21x1_ASAP7_75t_L g354 ( .A1(n_336), .A2(n_267), .B(n_335), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_298), .B(n_227), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_300), .A2(n_240), .B1(n_241), .B2(n_280), .C(n_282), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_295), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_303), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_284), .B1(n_267), .B2(n_279), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_289), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_307), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_296), .A2(n_267), .B(n_216), .Y(n_363) );
NOR3xp33_ASAP7_75t_SL g364 ( .A(n_329), .B(n_230), .C(n_287), .Y(n_364) );
CKINVDCx11_ASAP7_75t_R g365 ( .A(n_290), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_308), .A2(n_274), .B1(n_273), .B2(n_286), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_314), .A2(n_242), .B(n_276), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_303), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_363), .A2(n_309), .B(n_335), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_356), .A2(n_313), .B1(n_325), .B2(n_333), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_366), .A2(n_317), .B1(n_240), .B2(n_241), .C(n_328), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_356), .A2(n_313), .B1(n_333), .B2(n_328), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_349), .A2(n_363), .B(n_352), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_307), .B1(n_321), .B2(n_253), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_349), .A2(n_242), .B(n_304), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_355), .B(n_313), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_366), .A2(n_327), .B1(n_291), .B2(n_316), .C(n_290), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_360), .A2(n_273), .B1(n_274), .B2(n_253), .C(n_271), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_340), .A2(n_310), .B1(n_305), .B2(n_318), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_275), .B(n_254), .C(n_266), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_360), .A2(n_310), .B1(n_337), .B2(n_307), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_343), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_309), .B(n_326), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_367), .A2(n_336), .B(n_277), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_344), .A2(n_245), .B(n_320), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_341), .A2(n_321), .B1(n_234), .B2(n_245), .Y(n_389) );
AO31x2_ASAP7_75t_L g390 ( .A1(n_351), .A2(n_304), .A3(n_330), .B(n_298), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_342), .A2(n_361), .B1(n_341), .B2(n_344), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_341), .A2(n_337), .B1(n_311), .B2(n_306), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_357), .B(n_311), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_340), .A2(n_327), .B1(n_306), .B2(n_330), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_346), .A2(n_266), .B(n_275), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_390), .B(n_355), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_390), .B(n_345), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_373), .Y(n_398) );
OAI33xp33_ASAP7_75t_L g399 ( .A1(n_395), .A2(n_348), .A3(n_302), .B1(n_364), .B2(n_222), .B3(n_219), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_374), .A2(n_354), .B(n_367), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_372), .A2(n_346), .B1(n_357), .B2(n_345), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_384), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_390), .B(n_350), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_379), .A2(n_302), .B1(n_364), .B2(n_357), .C(n_312), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_395), .A2(n_219), .A3(n_222), .B1(n_224), .B2(n_343), .B3(n_347), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_393), .Y(n_409) );
INVx4_ASAP7_75t_L g410 ( .A(n_385), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_390), .B(n_338), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_393), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_382), .A2(n_357), .B1(n_350), .B2(n_338), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_385), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_390), .B(n_350), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_377), .B(n_347), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_362), .A3(n_339), .B(n_358), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_376), .B(n_347), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_385), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
AO21x1_ASAP7_75t_SL g424 ( .A1(n_376), .A2(n_362), .B(n_339), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_383), .A2(n_339), .B1(n_362), .B2(n_358), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_380), .Y(n_427) );
OAI332xp33_ASAP7_75t_L g428 ( .A1(n_371), .A2(n_224), .A3(n_365), .B1(n_353), .B2(n_19), .B3(n_247), .C1(n_185), .C2(n_180), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_370), .A2(n_339), .B1(n_362), .B2(n_358), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_416), .B(n_353), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_416), .B(n_353), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_403), .Y(n_432) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_423), .B(n_362), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_403), .B(n_391), .Y(n_434) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_406), .A2(n_378), .B1(n_381), .B2(n_388), .C1(n_392), .C2(n_312), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_416), .B(n_368), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_428), .B(n_312), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_404), .B(n_387), .Y(n_441) );
AOI31xp33_ASAP7_75t_L g442 ( .A1(n_426), .A2(n_389), .A3(n_19), .B(n_359), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_406), .B(n_194), .C(n_174), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_423), .B(n_339), .Y(n_445) );
AND2x4_ASAP7_75t_SL g446 ( .A(n_410), .B(n_358), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_401), .B(n_368), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
INVx5_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
AOI221x1_ASAP7_75t_L g452 ( .A1(n_413), .A2(n_368), .B1(n_359), .B2(n_217), .C(n_216), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_398), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_396), .A2(n_185), .A3(n_180), .B1(n_177), .B2(n_169), .B3(n_359), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_396), .B(n_209), .Y(n_457) );
NOR2xp67_ASAP7_75t_L g458 ( .A(n_428), .B(n_234), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_419), .B(n_174), .C(n_176), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_398), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_398), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_402), .B(n_209), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_409), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_419), .B(n_169), .C(n_177), .D(n_257), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_397), .B(n_217), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_415), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_397), .B(n_217), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
AOI222xp33_ASAP7_75t_L g473 ( .A1(n_399), .A2(n_209), .B1(n_216), .B2(n_234), .C1(n_332), .C2(n_323), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_415), .B(n_324), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_422), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_422), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_425), .B(n_216), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_427), .B(n_323), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_450), .B(n_425), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_438), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_460), .B(n_422), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_472), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_442), .B(n_399), .C(n_408), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_472), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_453), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_430), .B(n_424), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_444), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_430), .B(n_427), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_449), .B(n_427), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_418), .B(n_405), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_455), .B(n_421), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_451), .B(n_412), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_462), .Y(n_496) );
NAND2xp33_ASAP7_75t_SL g497 ( .A(n_460), .B(n_413), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_431), .B(n_420), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_456), .B(n_421), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_461), .B(n_412), .Y(n_502) );
NAND2xp33_ASAP7_75t_L g503 ( .A(n_451), .B(n_429), .Y(n_503) );
AOI33xp33_ASAP7_75t_L g504 ( .A1(n_465), .A2(n_426), .A3(n_418), .B1(n_405), .B2(n_414), .B3(n_408), .Y(n_504) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_451), .B(n_420), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_436), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_451), .B(n_405), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_451), .Y(n_509) );
NOR2xp33_ASAP7_75t_R g510 ( .A(n_437), .B(n_234), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_434), .B(n_400), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_471), .B(n_400), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_448), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_471), .B(n_400), .Y(n_516) );
NOR4xp25_ASAP7_75t_SL g517 ( .A(n_475), .B(n_400), .C(n_25), .D(n_27), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_437), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_445), .Y(n_520) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_435), .B(n_414), .C(n_260), .D(n_261), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_457), .B(n_400), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_414), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_439), .B(n_332), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_457), .B(n_441), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_441), .B(n_194), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_441), .B(n_194), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_469), .B(n_194), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_476), .B(n_174), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_476), .B(n_174), .Y(n_530) );
INVx4_ASAP7_75t_L g531 ( .A(n_437), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_439), .B(n_22), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_477), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_470), .B(n_174), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_440), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_479), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_479), .Y(n_537) );
INVx5_ASAP7_75t_L g538 ( .A(n_509), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_531), .A2(n_458), .B1(n_443), .B2(n_440), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_483), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_484), .A2(n_454), .B1(n_459), .B2(n_460), .Y(n_542) );
AOI22xp5_ASAP7_75t_SL g543 ( .A1(n_509), .A2(n_460), .B1(n_440), .B2(n_468), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_510), .Y(n_544) );
OAI211xp5_ASAP7_75t_SL g545 ( .A1(n_524), .A2(n_473), .B(n_464), .C(n_478), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_532), .A2(n_477), .B1(n_460), .B2(n_468), .C(n_467), .Y(n_546) );
OAI221xp5_ASAP7_75t_SL g547 ( .A1(n_522), .A2(n_468), .B1(n_446), .B2(n_452), .C(n_323), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_508), .B(n_446), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_509), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_489), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_487), .B(n_492), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_501), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_489), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_514), .B(n_474), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_496), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_496), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_501), .B(n_474), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_503), .A2(n_474), .B1(n_332), .B2(n_334), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_506), .B(n_194), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_500), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_509), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_531), .A2(n_334), .B1(n_315), .B2(n_324), .Y(n_564) );
NAND2x1_ASAP7_75t_SL g565 ( .A(n_531), .B(n_334), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_509), .B(n_324), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_176), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_502), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_176), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_480), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_513), .B(n_176), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_497), .A2(n_176), .B1(n_260), .B2(n_261), .C(n_315), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_483), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_491), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_485), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_503), .A2(n_495), .B(n_482), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_491), .Y(n_579) );
NOR4xp25_ASAP7_75t_L g580 ( .A(n_519), .B(n_326), .C(n_42), .D(n_43), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_487), .B(n_31), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_521), .A2(n_45), .B(n_46), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_498), .B(n_47), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_518), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_513), .B(n_48), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_505), .A2(n_324), .B1(n_319), .B2(n_315), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_543), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_544), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_576), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_536), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_574), .B(n_511), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_541), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_515), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_575), .B(n_515), .Y(n_596) );
OAI21xp33_ASAP7_75t_SL g597 ( .A1(n_549), .A2(n_525), .B(n_507), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_579), .B(n_498), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_563), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_538), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_540), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_552), .B(n_525), .Y(n_602) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_546), .B(n_522), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_553), .B(n_490), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_570), .A2(n_512), .B1(n_516), .B2(n_494), .C1(n_520), .C2(n_490), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_550), .B(n_516), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_539), .A2(n_535), .B(n_526), .C(n_527), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_538), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_578), .B(n_535), .Y(n_611) );
NOR4xp25_ASAP7_75t_SL g612 ( .A(n_547), .B(n_504), .C(n_517), .D(n_526), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_539), .B(n_530), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_557), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_560), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_583), .B(n_512), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_559), .A2(n_523), .B1(n_533), .B2(n_486), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_582), .A2(n_523), .B(n_527), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_585), .B(n_533), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_562), .B(n_488), .Y(n_621) );
O2A1O1Ixp5_ASAP7_75t_L g622 ( .A1(n_549), .A2(n_488), .B(n_485), .C(n_529), .Y(n_622) );
NOR4xp25_ASAP7_75t_SL g623 ( .A(n_572), .B(n_530), .C(n_529), .D(n_493), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_581), .A2(n_534), .B(n_528), .C(n_493), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_597), .A2(n_580), .B1(n_545), .B2(n_542), .C(n_548), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_617), .B(n_576), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g627 ( .A1(n_588), .A2(n_565), .B(n_559), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_588), .A2(n_542), .B(n_538), .Y(n_628) );
AOI322xp5_ASAP7_75t_L g629 ( .A1(n_589), .A2(n_555), .A3(n_584), .B1(n_538), .B2(n_577), .C1(n_573), .C2(n_540), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_591), .Y(n_631) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_608), .A2(n_555), .B(n_587), .C(n_558), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_599), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_611), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_611), .A2(n_566), .B(n_587), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_607), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_609), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_614), .A2(n_566), .B1(n_586), .B2(n_564), .C(n_569), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g641 ( .A(n_622), .B(n_567), .C(n_561), .Y(n_641) );
XNOR2x1_ASAP7_75t_L g642 ( .A(n_603), .B(n_577), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_613), .Y(n_643) );
OAI21xp33_ASAP7_75t_SL g644 ( .A1(n_605), .A2(n_573), .B(n_571), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_603), .A2(n_534), .B(n_528), .Y(n_645) );
XNOR2x1_ASAP7_75t_L g646 ( .A(n_602), .B(n_51), .Y(n_646) );
NOR2x1p5_ASAP7_75t_SL g647 ( .A(n_601), .B(n_493), .Y(n_647) );
AOI21xp5_ASAP7_75t_SL g648 ( .A1(n_628), .A2(n_624), .B(n_590), .Y(n_648) );
O2A1O1Ixp5_ASAP7_75t_L g649 ( .A1(n_628), .A2(n_600), .B(n_610), .C(n_622), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_631), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_646), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_634), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_627), .B(n_610), .C(n_600), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_644), .A2(n_610), .B(n_624), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_625), .A2(n_592), .B(n_619), .C(n_606), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_642), .A2(n_590), .B(n_623), .Y(n_656) );
AOI222xp33_ASAP7_75t_L g657 ( .A1(n_625), .A2(n_618), .B1(n_616), .B2(n_615), .C1(n_620), .C2(n_621), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_635), .A2(n_595), .B(n_596), .Y(n_658) );
OAI31xp33_ASAP7_75t_L g659 ( .A1(n_640), .A2(n_598), .A3(n_604), .B(n_601), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_630), .B(n_612), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_637), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_645), .B(n_493), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_633), .A2(n_324), .B1(n_319), .B2(n_315), .C(n_277), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_636), .A2(n_319), .B(n_315), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g665 ( .A(n_632), .B(n_52), .Y(n_665) );
OAI21x1_ASAP7_75t_SL g666 ( .A1(n_630), .A2(n_56), .B(n_57), .Y(n_666) );
AOI221x1_ASAP7_75t_L g667 ( .A1(n_641), .A2(n_319), .B1(n_277), .B2(n_69), .C(n_75), .Y(n_667) );
NOR4xp75_ASAP7_75t_L g668 ( .A(n_640), .B(n_59), .C(n_62), .D(n_319), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_638), .B(n_277), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_652), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_660), .A2(n_655), .B1(n_651), .B2(n_662), .C1(n_658), .C2(n_665), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_657), .B(n_656), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_659), .B(n_654), .Y(n_673) );
NOR2x2_ASAP7_75t_L g674 ( .A(n_671), .B(n_660), .Y(n_674) );
OR3x1_ASAP7_75t_L g675 ( .A(n_672), .B(n_648), .C(n_649), .Y(n_675) );
OR4x2_ASAP7_75t_L g676 ( .A(n_673), .B(n_653), .C(n_668), .D(n_629), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_675), .A2(n_670), .B1(n_650), .B2(n_661), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_674), .B(n_626), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_674), .B1(n_676), .B2(n_664), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_677), .A3(n_643), .B1(n_639), .B2(n_669), .C1(n_667), .C2(n_666), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_663), .B(n_647), .Y(n_681) );
endmodule