module fake_jpeg_29491_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_47),
.B1(n_41),
.B2(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_60),
.Y(n_65)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_52),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_41),
.B1(n_1),
.B2(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_13),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_7),
.B(n_8),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_5),
.CI(n_6),
.CON(n_79),
.SN(n_79)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_32),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_30),
.B(n_31),
.Y(n_91)
);

OA21x2_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_9),
.B(n_11),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_12),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_18),
.B(n_21),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_33),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_40),
.B1(n_93),
.B2(n_92),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_36),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_101),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_105),
.B1(n_104),
.B2(n_107),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_112),
.B(n_98),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_103),
.C(n_114),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_95),
.C(n_102),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_94),
.Y(n_119)
);


endmodule