module fake_aes_4333_n_533 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_533);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_533;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_70;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g69 ( .A(n_11), .Y(n_69) );
NOR2xp33_ASAP7_75t_L g70 ( .A(n_9), .B(n_47), .Y(n_70) );
INVx2_ASAP7_75t_L g71 ( .A(n_30), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_62), .Y(n_72) );
CKINVDCx20_ASAP7_75t_R g73 ( .A(n_66), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_11), .Y(n_74) );
NOR2xp33_ASAP7_75t_L g75 ( .A(n_28), .B(n_29), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_15), .Y(n_76) );
INVxp33_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_26), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_58), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_52), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_34), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_37), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_9), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_3), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_8), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_54), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_0), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_45), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_42), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_51), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_53), .Y(n_98) );
INVx3_ASAP7_75t_L g99 ( .A(n_2), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_35), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_59), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
BUFx5_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_56), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_43), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_99), .B(n_0), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_99), .B(n_1), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_99), .B(n_1), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_105), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_80), .B(n_2), .Y(n_112) );
NOR2x1_ASAP7_75t_L g113 ( .A(n_99), .B(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_89), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_89), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_69), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_105), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_78), .B(n_4), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_74), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_77), .B(n_5), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_105), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_78), .B(n_5), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_71), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_103), .B(n_6), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_72), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_72), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_73), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_104), .B(n_6), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_129), .Y(n_138) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_136), .A2(n_107), .B(n_106), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_134), .B(n_86), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_134), .B(n_87), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g145 ( .A1(n_135), .A2(n_90), .B1(n_88), .B2(n_96), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_134), .B(n_76), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_129), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_108), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_108), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_123), .A2(n_92), .B1(n_74), .B2(n_76), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_126), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_131), .B(n_93), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_116), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_116), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_126), .B(n_83), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_109), .B(n_107), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_123), .B(n_92), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_116), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_130), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_128), .B1(n_123), .B2(n_110), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_163), .B(n_130), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_170), .A2(n_130), .B1(n_125), .B2(n_136), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_164), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_154), .B(n_123), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_159), .B(n_125), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_164), .A2(n_128), .B1(n_123), .B2(n_109), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_146), .B(n_131), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_154), .B(n_128), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_146), .B(n_109), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_146), .B(n_164), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_146), .A2(n_128), .B1(n_110), .B2(n_132), .Y(n_203) );
AO22x1_ASAP7_75t_L g204 ( .A1(n_165), .A2(n_128), .B1(n_110), .B2(n_113), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
OR2x6_ASAP7_75t_L g206 ( .A(n_165), .B(n_113), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_140), .B(n_132), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx5_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_142), .B(n_137), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
OAI221xp5_ASAP7_75t_L g213 ( .A1(n_176), .A2(n_145), .B1(n_112), .B2(n_157), .C(n_102), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_177), .Y(n_214) );
BUFx10_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_183), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_198), .B(n_165), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_198), .B(n_139), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_172), .A2(n_139), .B(n_158), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_193), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_183), .B(n_139), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_205), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_172), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_188), .B(n_137), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_178), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_187), .B(n_137), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_189), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
AND2x2_ASAP7_75t_SL g235 ( .A(n_191), .B(n_117), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_175), .B(n_112), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_187), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
INVx6_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
INVx5_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_173), .A2(n_117), .B1(n_118), .B2(n_137), .Y(n_243) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_196), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_199), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_188), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_203), .B(n_117), .Y(n_247) );
INVx6_ASAP7_75t_L g248 ( .A(n_188), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_248), .A2(n_197), .B1(n_206), .B2(n_212), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_185), .B(n_181), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_181), .B(n_182), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_233), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g253 ( .A1(n_213), .A2(n_207), .B1(n_203), .B2(n_195), .C(n_173), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_228), .B(n_197), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_228), .B(n_197), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_226), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_218), .A2(n_190), .B1(n_197), .B2(n_185), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_225), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_204), .B1(n_211), .B2(n_212), .C(n_190), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g261 ( .A1(n_217), .A2(n_206), .B1(n_182), .B2(n_194), .C(n_179), .Y(n_261) );
AOI21xp33_ASAP7_75t_L g262 ( .A1(n_222), .A2(n_206), .B(n_194), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_248), .A2(n_206), .B1(n_186), .B2(n_179), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_248), .A2(n_206), .B1(n_186), .B2(n_179), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_231), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_242), .B(n_174), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_204), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_223), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_220), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_246), .B(n_174), .Y(n_272) );
OAI222xp33_ASAP7_75t_L g273 ( .A1(n_243), .A2(n_102), .B1(n_137), .B2(n_84), .C1(n_85), .C2(n_94), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_260), .A2(n_232), .B(n_241), .C(n_237), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_257), .A2(n_248), .B1(n_221), .B2(n_224), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_247), .B1(n_232), .B2(n_241), .C(n_237), .Y(n_277) );
AO22x1_ASAP7_75t_L g278 ( .A1(n_252), .A2(n_222), .B1(n_242), .B2(n_101), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_221), .B1(n_224), .B2(n_229), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_256), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_268), .A2(n_215), .B1(n_245), .B2(n_235), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_261), .A2(n_229), .B1(n_235), .B2(n_222), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_252), .A2(n_133), .B(n_117), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_254), .B(n_245), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_250), .A2(n_234), .B(n_227), .Y(n_285) );
AO22x1_ASAP7_75t_L g286 ( .A1(n_268), .A2(n_222), .B1(n_242), .B2(n_91), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_249), .A2(n_230), .B1(n_239), .B2(n_186), .C(n_179), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_215), .B1(n_235), .B2(n_231), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_230), .B1(n_239), .B2(n_186), .C(n_174), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_234), .B1(n_227), .B2(n_214), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_270), .Y(n_291) );
AOI21xp33_ASAP7_75t_L g292 ( .A1(n_258), .A2(n_216), .B(n_244), .Y(n_292) );
AOI222xp33_ASAP7_75t_L g293 ( .A1(n_254), .A2(n_215), .B1(n_231), .B2(n_114), .C1(n_115), .C2(n_119), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g294 ( .A1(n_269), .A2(n_215), .B1(n_242), .B2(n_238), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_256), .A2(n_274), .A3(n_263), .B(n_259), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_280), .B(n_259), .Y(n_297) );
AOI222xp33_ASAP7_75t_L g298 ( .A1(n_276), .A2(n_254), .B1(n_255), .B2(n_273), .C1(n_269), .C2(n_98), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_284), .B(n_269), .Y(n_299) );
AOI33xp33_ASAP7_75t_L g300 ( .A1(n_296), .A2(n_119), .A3(n_114), .B1(n_115), .B2(n_85), .B3(n_94), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_293), .A2(n_282), .B1(n_277), .B2(n_255), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_279), .A2(n_255), .B1(n_262), .B2(n_265), .C(n_124), .Y(n_302) );
AOI211xp5_ASAP7_75t_L g303 ( .A1(n_286), .A2(n_262), .B(n_255), .C(n_266), .Y(n_303) );
INVx4_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_272), .B1(n_266), .B2(n_259), .C1(n_274), .C2(n_263), .Y(n_305) );
AOI33xp33_ASAP7_75t_L g306 ( .A1(n_294), .A2(n_95), .A3(n_100), .B1(n_81), .B2(n_98), .B3(n_84), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_295), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_295), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_295), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_288), .A2(n_272), .B1(n_271), .B2(n_239), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_272), .B1(n_271), .B2(n_239), .Y(n_311) );
AO22x1_ASAP7_75t_L g312 ( .A1(n_291), .A2(n_274), .B1(n_263), .B2(n_272), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_289), .A2(n_231), .B1(n_238), .B2(n_214), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_275), .A2(n_251), .B(n_118), .C(n_117), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_278), .B(n_70), .C(n_100), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_285), .B(n_251), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_283), .A2(n_267), .B1(n_242), .B2(n_292), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_280), .B(n_124), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_304), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_297), .B(n_124), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_309), .B(n_118), .Y(n_326) );
AOI221x1_ASAP7_75t_L g327 ( .A1(n_317), .A2(n_97), .B1(n_106), .B2(n_95), .C(n_270), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_297), .B(n_97), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_308), .B(n_118), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_322), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_322), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_321), .B(n_105), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_299), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_301), .A2(n_267), .B1(n_270), .B2(n_242), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_320), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_317), .A2(n_267), .B1(n_270), .B2(n_220), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_321), .B(n_105), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_298), .A2(n_105), .B1(n_79), .B2(n_83), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_320), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_303), .B(n_71), .C(n_79), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_321), .B(n_118), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_307), .B(n_127), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_307), .B(n_127), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_307), .B(n_7), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_166), .B(n_158), .Y(n_349) );
OAI221xp5_ASAP7_75t_SL g350 ( .A1(n_306), .A2(n_122), .B1(n_111), .B2(n_120), .C(n_121), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_318), .B(n_127), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_302), .A2(n_133), .B1(n_75), .B2(n_120), .C(n_121), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_312), .B(n_270), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_318), .B(n_122), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_7), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_305), .B(n_122), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_305), .A2(n_216), .B1(n_240), .B2(n_192), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_300), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_348), .B(n_314), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_356), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_314), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_356), .B(n_304), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_330), .B(n_331), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_333), .B(n_303), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_324), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_324), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_326), .B(n_314), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_329), .B(n_316), .Y(n_376) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_324), .B(n_319), .Y(n_377) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_327), .B(n_310), .C(n_311), .D(n_313), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_352), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_353), .B(n_8), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_335), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_332), .B(n_10), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_332), .B(n_12), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_352), .Y(n_385) );
AOI211x1_ASAP7_75t_L g386 ( .A1(n_361), .A2(n_12), .B(n_13), .C(n_14), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_328), .B(n_13), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_14), .Y(n_388) );
AOI31xp33_ASAP7_75t_L g389 ( .A1(n_343), .A2(n_16), .A3(n_111), .B(n_120), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_352), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_325), .B(n_16), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_340), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_347), .B(n_111), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_350), .B(n_17), .Y(n_394) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_347), .B(n_270), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_357), .B(n_121), .Y(n_398) );
OAI33xp33_ASAP7_75t_L g399 ( .A1(n_351), .A2(n_162), .A3(n_166), .B1(n_167), .B2(n_192), .B3(n_200), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_357), .B(n_133), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g401 ( .A1(n_338), .A2(n_18), .B(n_20), .C(n_21), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_169), .B1(n_144), .B2(n_147), .C(n_149), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_351), .A2(n_167), .B(n_162), .C(n_201), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_355), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_359), .B(n_23), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_334), .B(n_24), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_359), .B(n_171), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_344), .B(n_171), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_369), .B(n_344), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_368), .B(n_346), .Y(n_410) );
INVx4_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_396), .B(n_346), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_327), .B(n_336), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
INVxp33_ASAP7_75t_L g415 ( .A(n_393), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_367), .B(n_355), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_392), .B(n_345), .Y(n_417) );
AOI32xp33_ASAP7_75t_L g418 ( .A1(n_380), .A2(n_345), .A3(n_354), .B1(n_355), .B2(n_360), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_386), .B(n_355), .C(n_138), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_364), .B(n_367), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_365), .B(n_349), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_401), .B(n_138), .C(n_144), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_401), .A2(n_349), .B(n_220), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_371), .B(n_349), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_371), .B(n_27), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_370), .B(n_138), .Y(n_427) );
OAI222xp33_ASAP7_75t_L g428 ( .A1(n_372), .A2(n_160), .B1(n_32), .B2(n_33), .C1(n_36), .C2(n_40), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_378), .B(n_31), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_372), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_404), .B(n_41), .Y(n_431) );
XOR2xp5_ASAP7_75t_L g432 ( .A(n_388), .B(n_44), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_379), .B(n_171), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_389), .B(n_387), .C(n_391), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_373), .B(n_169), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_379), .B(n_46), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_397), .B(n_169), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_395), .B(n_220), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_382), .B(n_48), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_366), .B(n_161), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_405), .A2(n_220), .B(n_161), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_407), .A2(n_169), .B1(n_161), .B2(n_171), .C(n_149), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_390), .B(n_169), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_390), .B(n_50), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_375), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_362), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
NAND2xp33_ASAP7_75t_L g450 ( .A(n_377), .B(n_161), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_383), .B(n_55), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_408), .B(n_406), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_57), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_448), .B(n_400), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g455 ( .A(n_411), .B(n_394), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_418), .A2(n_402), .B(n_403), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_430), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_432), .B(n_60), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_411), .B(n_399), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_434), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_449), .B(n_171), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_435), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_448), .B(n_161), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_414), .Y(n_464) );
XOR2x2_ASAP7_75t_L g465 ( .A(n_436), .B(n_416), .Y(n_465) );
XNOR2x1_ASAP7_75t_L g466 ( .A(n_421), .B(n_63), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_409), .B(n_64), .Y(n_467) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_431), .B(n_144), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_447), .B(n_68), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_410), .B(n_144), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_436), .B(n_147), .C(n_149), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_412), .B(n_147), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_423), .B(n_147), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_417), .B(n_160), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_429), .B(n_160), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_422), .B(n_160), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_430), .B(n_160), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_443), .A2(n_240), .B1(n_160), .B2(n_210), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_441), .A2(n_240), .B1(n_209), .B2(n_202), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g485 ( .A1(n_415), .A2(n_208), .B(n_210), .C(n_428), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_426), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_441), .A2(n_208), .A3(n_210), .B(n_451), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_452), .B(n_210), .Y(n_489) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_420), .A2(n_210), .B(n_208), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_413), .A2(n_450), .B1(n_451), .B2(n_438), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_452), .B(n_425), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_450), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_442), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_452), .B(n_440), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_453), .A2(n_446), .B1(n_440), .B2(n_444), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_424), .B(n_411), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g499 ( .A(n_432), .B(n_333), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_430), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_436), .A2(n_389), .B(n_429), .C(n_428), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_472), .B(n_459), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_501), .A2(n_472), .B(n_485), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_501), .A2(n_498), .B(n_488), .C(n_455), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_469), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_486), .B(n_495), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
OA22x2_ASAP7_75t_L g509 ( .A1(n_499), .A2(n_479), .B1(n_458), .B2(n_460), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_456), .B(n_478), .C(n_463), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_491), .A2(n_493), .B1(n_479), .B2(n_454), .Y(n_511) );
XNOR2x1_ASAP7_75t_L g512 ( .A(n_466), .B(n_462), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_491), .A2(n_494), .B1(n_476), .B2(n_475), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_474), .A2(n_493), .B(n_482), .Y(n_514) );
OAI211xp5_ASAP7_75t_SL g515 ( .A1(n_503), .A2(n_496), .B(n_490), .C(n_489), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_510), .B(n_464), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_507), .B(n_492), .Y(n_517) );
NAND4xp25_ASAP7_75t_L g518 ( .A(n_504), .B(n_467), .C(n_470), .D(n_484), .Y(n_518) );
AOI21xp33_ASAP7_75t_SL g519 ( .A1(n_509), .A2(n_457), .B(n_500), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_511), .A2(n_487), .B1(n_477), .B2(n_497), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_506), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_519), .B(n_505), .C(n_502), .Y(n_522) );
NAND5xp2_ASAP7_75t_L g523 ( .A(n_520), .B(n_514), .C(n_513), .D(n_473), .E(n_512), .Y(n_523) );
NAND2xp33_ASAP7_75t_SL g524 ( .A(n_516), .B(n_468), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_515), .A2(n_507), .B1(n_508), .B2(n_483), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_525), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_522), .A2(n_516), .B1(n_518), .B2(n_521), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_527), .A2(n_523), .B1(n_524), .B2(n_517), .C(n_481), .Y(n_528) );
XNOR2xp5_ASAP7_75t_L g529 ( .A(n_526), .B(n_471), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_529), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_530), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_531), .A2(n_528), .B(n_480), .C(n_461), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_532), .A2(n_461), .B(n_480), .Y(n_533) );
endmodule