module real_jpeg_30105_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_244;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_1),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_67),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_31),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_5),
.A2(n_47),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_47),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_51),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_54),
.B1(n_224),
.B2(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_32),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_6),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_135),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_135),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_135),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_10),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_183)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_25),
.B1(n_47),
.B2(n_48),
.Y(n_244)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_98),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_98),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_98),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_16),
.A2(n_56),
.B1(n_57),
.B2(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_76),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_21),
.B(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_22),
.B(n_77),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_22),
.Y(n_280)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.CI(n_52),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_38),
.C(n_52),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_26),
.A2(n_35),
.B(n_139),
.C(n_140),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_28),
.A2(n_31),
.B1(n_134),
.B2(n_163),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_31),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_32),
.A2(n_48),
.A3(n_241),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_33),
.B(n_139),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_36),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_41),
.B1(n_51),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_41),
.A2(n_51),
.B1(n_161),
.B2(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_42),
.A2(n_46),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_42),
.A2(n_46),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_42),
.A2(n_46),
.B1(n_144),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_42),
.A2(n_46),
.B1(n_181),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_48),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_47),
.A2(n_57),
.A3(n_72),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_47),
.B(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_68),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_53),
.B(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_66),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_61),
.B1(n_63),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_54),
.A2(n_63),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_54),
.A2(n_63),
.B1(n_218),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_54),
.A2(n_63),
.B1(n_213),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_55),
.A2(n_64),
.B1(n_92),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_55),
.A2(n_64),
.B1(n_142),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_55),
.A2(n_64),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_56),
.B(n_73),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_56),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_65),
.B(n_139),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_70),
.A2(n_71),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_70),
.A2(n_71),
.B1(n_199),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_70),
.A2(n_71),
.B1(n_166),
.B2(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_71),
.B(n_139),
.Y(n_225)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_81),
.A2(n_84),
.B1(n_95),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_81),
.A2(n_84),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_86),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_99),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_93),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_99),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_97),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_100),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_122),
.B2(n_123),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_110),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_108),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_118),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_149),
.B(n_278),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_147),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_128),
.B(n_147),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_146),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_146),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.C(n_143),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_186),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_169),
.B(n_185),
.Y(n_151)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_167),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.C(n_164),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_173),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_276),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_176),
.Y(n_276)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_179),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_182),
.B(n_184),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_183),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.C(n_189),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_272),
.B(n_277),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_258),
.B(n_271),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_234),
.B(n_257),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_214),
.B(n_233),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_209),
.C(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_212),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_221),
.B(n_232),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_220),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_231),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_225),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_246),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_253),
.Y(n_266)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_267),
.C(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);


endmodule