module fake_aes_6876_n_1134 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1134);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1134;
wire n_663;
wire n_791;
wire n_707;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1097;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_1078;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_950;
wire n_427;
wire n_910;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_570;
wire n_508;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_45), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_179), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_6), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_120), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_145), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_140), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_129), .B(n_63), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_241), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_245), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_11), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_190), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_185), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_98), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_77), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_160), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_133), .Y(n_279) );
CKINVDCx16_ASAP7_75t_R g280 ( .A(n_17), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_19), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_191), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_243), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_136), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_101), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_77), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_197), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_1), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_27), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_148), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_91), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_22), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_260), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_53), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_218), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_108), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_168), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_194), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_87), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_90), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_41), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_72), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_25), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_180), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_88), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_173), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_213), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_124), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_163), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_170), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_92), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g315 ( .A(n_144), .B(n_89), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_138), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_34), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_217), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_132), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_198), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_127), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_201), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_137), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_11), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_102), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_141), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_115), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_224), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_244), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_44), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_178), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_59), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_39), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_71), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_211), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_63), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_48), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_99), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_195), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_58), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_119), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_208), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_112), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_223), .B(n_236), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_186), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_86), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_155), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_20), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_84), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_205), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_222), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_238), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_12), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_82), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_15), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_13), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_82), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_106), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_182), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_85), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_258), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_183), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_103), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_162), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_151), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_6), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_2), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_228), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_35), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_193), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_154), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_126), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_196), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_212), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_50), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_189), .B(n_139), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_23), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_74), .Y(n_380) );
INVxp33_ASAP7_75t_L g381 ( .A(n_5), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_125), .B(n_109), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_158), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_27), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_184), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_79), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_105), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_225), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_131), .Y(n_389) );
CKINVDCx14_ASAP7_75t_R g390 ( .A(n_149), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_227), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_62), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_253), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_130), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_31), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_192), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_153), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_0), .Y(n_398) );
BUFx5_ASAP7_75t_L g399 ( .A(n_206), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_188), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_249), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_248), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_221), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_229), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_81), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_341), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_364), .B(n_0), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_341), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_381), .B(n_1), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_316), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_364), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_316), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_266), .B(n_2), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g414 ( .A(n_399), .B(n_93), .Y(n_414) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_296), .B(n_259), .Y(n_415) );
INVxp33_ASAP7_75t_SL g416 ( .A(n_262), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_267), .A2(n_95), .B(n_94), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_335), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_335), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_381), .B(n_3), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_316), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_265), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_399), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_267), .A2(n_97), .B(n_96), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_279), .B(n_3), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_268), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_262), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_299), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g432 ( .A1(n_305), .A2(n_7), .B1(n_4), .B2(n_5), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_271), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_273), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_264), .B(n_4), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_275), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_280), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_290), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_399), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_316), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_329), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_348), .B(n_8), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_272), .B(n_9), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_430), .B(n_290), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
BUFx4f_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_407), .B(n_263), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_414), .B(n_278), .C(n_276), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_430), .B(n_390), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_409), .A2(n_286), .B1(n_288), .B2(n_277), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_416), .B(n_347), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_422), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
BUFx10_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_415), .B(n_263), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_415), .B(n_274), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_411), .B(n_293), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_419), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_439), .B(n_349), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_439), .B(n_353), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_410), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
AND2x6_ASAP7_75t_L g472 ( .A(n_411), .B(n_428), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_426), .B(n_269), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_431), .Y(n_475) );
AND2x6_ASAP7_75t_L g476 ( .A(n_411), .B(n_299), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_390), .Y(n_477) );
INVx5_ASAP7_75t_L g478 ( .A(n_410), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_443), .A2(n_270), .B1(n_375), .B2(n_338), .Y(n_479) );
INVxp33_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
NOR2x1p5_ASAP7_75t_L g481 ( .A(n_428), .B(n_337), .Y(n_481) );
OR2x2_ASAP7_75t_SL g482 ( .A(n_432), .B(n_435), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_424), .B(n_360), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_429), .B(n_337), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_410), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_429), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_433), .B(n_338), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_419), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_425), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_433), .B(n_282), .Y(n_490) );
INVx5_ASAP7_75t_L g491 ( .A(n_410), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_434), .A2(n_333), .B1(n_334), .B2(n_325), .Y(n_492) );
INVx5_ASAP7_75t_L g493 ( .A(n_476), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_457), .B(n_434), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_465), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_486), .B(n_437), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_447), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_477), .B(n_437), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_472), .A2(n_427), .B1(n_436), .B2(n_425), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_471), .B(n_362), .Y(n_500) );
AO22x1_ASAP7_75t_L g501 ( .A1(n_480), .A2(n_438), .B1(n_369), .B2(n_392), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_447), .B(n_283), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_462), .A2(n_413), .B1(n_270), .B2(n_375), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_477), .B(n_420), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_479), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_452), .B(n_435), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_452), .B(n_350), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_471), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_479), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_484), .B(n_420), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_484), .B(n_421), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_448), .A2(n_418), .B(n_426), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_487), .B(n_421), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_460), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_454), .B(n_284), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_472), .A2(n_427), .B1(n_436), .B2(n_425), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_467), .B(n_284), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_463), .A2(n_432), .B1(n_392), .B2(n_369), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_468), .B(n_319), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_445), .B(n_444), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_472), .A2(n_436), .B1(n_440), .B2(n_427), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_481), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_465), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_483), .B(n_319), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_453), .A2(n_438), .B1(n_395), .B2(n_351), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g529 ( .A(n_472), .B(n_378), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_465), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_472), .A2(n_440), .B1(n_408), .B2(n_406), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_460), .B(n_406), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_464), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_473), .Y(n_534) );
AND2x6_ASAP7_75t_SL g535 ( .A(n_482), .B(n_355), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_459), .B(n_365), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_482), .A2(n_386), .B1(n_405), .B2(n_305), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_461), .A2(n_303), .B1(n_357), .B2(n_356), .Y(n_539) );
INVx5_ASAP7_75t_L g540 ( .A(n_476), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_459), .B(n_408), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_459), .B(n_370), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_461), .B(n_386), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_490), .B(n_403), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_476), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_473), .B(n_404), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_474), .A2(n_418), .B(n_426), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_473), .B(n_404), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_461), .A2(n_440), .B1(n_359), .B2(n_368), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_492), .B(n_295), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_449), .A2(n_418), .B(n_377), .C(n_379), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_475), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_475), .B(n_340), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_449), .B(n_304), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_476), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_474), .A2(n_426), .B(n_382), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_476), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_461), .A2(n_380), .B1(n_384), .B2(n_358), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_450), .A2(n_317), .B1(n_371), .B2(n_398), .Y(n_560) );
AO22x1_ASAP7_75t_L g561 ( .A1(n_476), .A2(n_330), .B1(n_310), .B2(n_405), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_451), .B(n_352), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_458), .A2(n_287), .B1(n_291), .B2(n_289), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_466), .A2(n_292), .B1(n_298), .B2(n_294), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_466), .B(n_354), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_469), .B(n_328), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_469), .B(n_344), .Y(n_568) );
AO22x1_ASAP7_75t_L g569 ( .A1(n_488), .A2(n_300), .B1(n_306), .B2(n_301), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_474), .B(n_488), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_489), .B(n_376), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_489), .A2(n_307), .B1(n_309), .B2(n_308), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_556), .A2(n_346), .B(n_455), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_513), .A2(n_456), .B(n_455), .Y(n_574) );
OR2x6_ASAP7_75t_L g575 ( .A(n_501), .B(n_281), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_507), .Y(n_576) );
NOR2xp33_ASAP7_75t_SL g577 ( .A(n_570), .B(n_315), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_506), .B(n_494), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_547), .A2(n_312), .B(n_311), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_536), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_515), .A2(n_456), .B(n_455), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_506), .B(n_402), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_535), .Y(n_583) );
OR2x4_ASAP7_75t_L g584 ( .A(n_550), .B(n_281), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_543), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_521), .A2(n_318), .B(n_320), .C(n_313), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_511), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_532), .A2(n_323), .B(n_324), .C(n_321), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_523), .B(n_326), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_498), .B(n_281), .Y(n_590) );
INVx3_ASAP7_75t_SL g591 ( .A(n_505), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_551), .B(n_331), .C(n_327), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_552), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_541), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_527), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_508), .B(n_332), .Y(n_596) );
NOR3xp33_ASAP7_75t_L g597 ( .A(n_538), .B(n_528), .C(n_509), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_533), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_510), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_500), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_538), .B(n_10), .Y(n_602) );
OAI22x1_ASAP7_75t_L g603 ( .A1(n_519), .A2(n_339), .B1(n_343), .B2(n_336), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_503), .B(n_331), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_546), .B(n_345), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_548), .B(n_361), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_549), .A2(n_366), .B1(n_367), .B2(n_363), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_515), .A2(n_470), .B(n_456), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_496), .B(n_10), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_512), .B(n_372), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_552), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_516), .B(n_373), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_529), .A2(n_554), .B1(n_549), .B2(n_559), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_514), .B(n_374), .Y(n_614) );
INVx5_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_493), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_504), .B(n_383), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_539), .B(n_385), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_554), .A2(n_388), .B1(n_389), .B2(n_387), .Y(n_619) );
NOR2xp67_ASAP7_75t_SL g620 ( .A(n_493), .B(n_322), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_571), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_561), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_559), .B(n_393), .C(n_391), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_569), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_524), .A2(n_520), .B(n_518), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_495), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_562), .A2(n_485), .B(n_470), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_544), .B(n_396), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_526), .B(n_397), .Y(n_630) );
AOI33xp33_ASAP7_75t_L g631 ( .A1(n_560), .A2(n_400), .A3(n_401), .B1(n_302), .B2(n_314), .B3(n_394), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_524), .A2(n_297), .B1(n_302), .B2(n_285), .Y(n_632) );
AND2x6_ASAP7_75t_L g633 ( .A(n_558), .B(n_322), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_567), .A2(n_297), .B(n_314), .C(n_285), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_563), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_525), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_545), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_531), .B(n_394), .C(n_342), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_530), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_565), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_566), .A2(n_485), .B(n_478), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_537), .A2(n_491), .B(n_478), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_540), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_534), .A2(n_491), .B(n_478), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_502), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_553), .B(n_14), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_499), .B(n_517), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_517), .A2(n_442), .B(n_441), .C(n_342), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_542), .A2(n_522), .B(n_557), .C(n_555), .Y(n_650) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_522), .A2(n_442), .B(n_342), .C(n_329), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_500), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_500), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_541), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_507), .B(n_16), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_521), .A2(n_342), .B1(n_423), .B2(n_412), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_500), .B(n_16), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_505), .B(n_18), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_541), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_494), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_494), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_500), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_521), .A2(n_412), .B(n_423), .C(n_491), .Y(n_664) );
BUFx4f_ASAP7_75t_L g665 ( .A(n_507), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_556), .A2(n_446), .B(n_412), .Y(n_666) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_519), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_667) );
BUFx4f_ASAP7_75t_L g668 ( .A(n_507), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_497), .A2(n_423), .B1(n_412), .B2(n_23), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_541), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_506), .B(n_21), .Y(n_671) );
AND2x2_ASAP7_75t_SL g672 ( .A(n_543), .B(n_21), .Y(n_672) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_538), .B(n_22), .C(n_24), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_552), .Y(n_674) );
INVx4_ASAP7_75t_L g675 ( .A(n_493), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_556), .A2(n_446), .B(n_412), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_507), .B(n_24), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_497), .A2(n_423), .B1(n_412), .B2(n_28), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_556), .A2(n_446), .B(n_412), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_661), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_635), .B(n_25), .Y(n_681) );
AOI22x1_ASAP7_75t_SL g682 ( .A1(n_583), .A2(n_26), .B1(n_28), .B2(n_29), .Y(n_682) );
AO31x2_ASAP7_75t_L g683 ( .A1(n_651), .A2(n_423), .A3(n_446), .B(n_30), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_662), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_665), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_665), .Y(n_686) );
OAI22xp33_ASAP7_75t_SL g687 ( .A1(n_602), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_597), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_591), .A2(n_32), .B(n_33), .C(n_34), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_SL g690 ( .A1(n_664), .A2(n_152), .B(n_256), .C(n_254), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_653), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_581), .A2(n_104), .B(n_100), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_608), .A2(n_110), .B(n_107), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_586), .A2(n_36), .B(n_37), .C(n_39), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_668), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_621), .A2(n_40), .B(n_41), .C(n_42), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_622), .A2(n_40), .B(n_42), .C(n_43), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_676), .A2(n_113), .B(n_111), .Y(n_698) );
AND2x6_ASAP7_75t_L g699 ( .A(n_613), .B(n_43), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_679), .A2(n_116), .B(n_114), .Y(n_700) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_668), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_625), .Y(n_702) );
AOI221x1_ASAP7_75t_L g703 ( .A1(n_592), .A2(n_44), .B1(n_45), .B2(n_46), .C(n_47), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_613), .A2(n_46), .B(n_47), .C(n_48), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_599), .B(n_49), .Y(n_705) );
AO31x2_ASAP7_75t_L g706 ( .A1(n_649), .A2(n_49), .A3(n_50), .B(n_51), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_672), .B(n_51), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_592), .A2(n_118), .B(n_117), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_630), .A2(n_52), .B(n_54), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_574), .A2(n_122), .B(n_121), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_653), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_626), .A2(n_128), .B(n_123), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
BUFx8_ASAP7_75t_SL g714 ( .A(n_575), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_575), .Y(n_715) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_593), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_642), .A2(n_172), .B(n_251), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_587), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_584), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_595), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_640), .B(n_52), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_600), .B(n_54), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_648), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_578), .A2(n_171), .B(n_250), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_641), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_598), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_652), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_638), .A2(n_175), .B(n_247), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_663), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_596), .A2(n_61), .B1(n_64), .B2(n_65), .C(n_66), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_650), .A2(n_176), .B(n_246), .Y(n_731) );
INVx4_ASAP7_75t_L g732 ( .A(n_615), .Y(n_732) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_673), .A2(n_64), .B(n_65), .C(n_66), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_659), .B(n_67), .Y(n_734) );
INVx8_ASAP7_75t_L g735 ( .A(n_615), .Y(n_735) );
BUFx8_ASAP7_75t_L g736 ( .A(n_623), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_628), .A2(n_174), .B(n_242), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_609), .Y(n_738) );
AO31x2_ASAP7_75t_L g739 ( .A1(n_588), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_582), .B(n_68), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_658), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_631), .B(n_69), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_585), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_627), .Y(n_744) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_618), .B(n_70), .C(n_73), .D(n_74), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_605), .A2(n_177), .B(n_237), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_660), .B(n_73), .Y(n_747) );
BUFx4f_ASAP7_75t_L g748 ( .A(n_589), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_619), .B(n_75), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_646), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_647), .A2(n_75), .B(n_76), .C(n_78), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_655), .A2(n_76), .B1(n_78), .B2(n_80), .C(n_81), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_607), .A2(n_80), .B(n_83), .C(n_84), .Y(n_753) );
AOI221x1_ASAP7_75t_L g754 ( .A1(n_669), .A2(n_83), .B1(n_85), .B2(n_86), .C(n_134), .Y(n_754) );
AO31x2_ASAP7_75t_L g755 ( .A1(n_678), .A2(n_135), .A3(n_142), .B(n_143), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_636), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_660), .B(n_257), .Y(n_757) );
AO31x2_ASAP7_75t_L g758 ( .A1(n_632), .A2(n_146), .A3(n_147), .B(n_150), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_677), .A2(n_156), .B1(n_157), .B2(n_159), .Y(n_759) );
AO31x2_ASAP7_75t_L g760 ( .A1(n_590), .A2(n_161), .A3(n_164), .B(n_165), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g761 ( .A1(n_671), .A2(n_166), .B(n_167), .C(n_169), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_589), .B(n_187), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_603), .A2(n_199), .A3(n_200), .B(n_202), .Y(n_763) );
AO21x1_ASAP7_75t_L g764 ( .A1(n_577), .A2(n_203), .B(n_204), .Y(n_764) );
HB1xp67_ASAP7_75t_SL g765 ( .A(n_667), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_593), .Y(n_766) );
AO32x2_ASAP7_75t_L g767 ( .A1(n_577), .A2(n_207), .A3(n_209), .B1(n_210), .B2(n_215), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_606), .A2(n_216), .B(n_219), .Y(n_768) );
INVx2_ASAP7_75t_SL g769 ( .A(n_594), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_639), .Y(n_770) );
OR2x6_ASAP7_75t_L g771 ( .A(n_616), .B(n_220), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_654), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_604), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_624), .A2(n_226), .B1(n_230), .B2(n_231), .C(n_232), .Y(n_774) );
OAI21x1_ASAP7_75t_SL g775 ( .A1(n_644), .A2(n_233), .B(n_234), .Y(n_775) );
OR2x6_ASAP7_75t_L g776 ( .A(n_580), .B(n_235), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_617), .Y(n_777) );
NOR2x1_ASAP7_75t_SL g778 ( .A(n_615), .B(n_675), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_610), .A2(n_614), .B1(n_637), .B2(n_629), .Y(n_779) );
AOI221x1_ASAP7_75t_L g780 ( .A1(n_612), .A2(n_674), .B1(n_611), .B2(n_656), .C(n_645), .Y(n_780) );
BUFx2_ASAP7_75t_SL g781 ( .A(n_670), .Y(n_781) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_634), .A2(n_643), .B(n_657), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_675), .A2(n_644), .A3(n_633), .B(n_674), .Y(n_783) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_611), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_620), .A2(n_622), .B(n_621), .C(n_613), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_633), .B(n_576), .Y(n_786) );
NAND2xp33_ASAP7_75t_L g787 ( .A(n_633), .B(n_661), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_573), .A2(n_556), .B(n_447), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g789 ( .A1(n_584), .A2(n_479), .B1(n_543), .B2(n_509), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_665), .Y(n_790) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_597), .A2(n_653), .B1(n_519), .B2(n_507), .C(n_479), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_661), .Y(n_792) );
BUFx10_ASAP7_75t_L g793 ( .A(n_584), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_573), .A2(n_556), .B(n_447), .Y(n_794) );
AO31x2_ASAP7_75t_L g795 ( .A1(n_651), .A2(n_551), .A3(n_513), .B(n_649), .Y(n_795) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_735), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_699), .A2(n_789), .B1(n_791), .B2(n_707), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_686), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_735), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_684), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_787), .A2(n_782), .B(n_731), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_777), .A2(n_773), .B(n_742), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_792), .B(n_718), .Y(n_803) );
AO31x2_ASAP7_75t_L g804 ( .A1(n_703), .A2(n_764), .A3(n_754), .B(n_704), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_681), .B(n_701), .Y(n_805) );
AO31x2_ASAP7_75t_L g806 ( .A1(n_712), .A2(n_710), .A3(n_700), .B(n_698), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_732), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_741), .B(n_705), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_720), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_699), .A2(n_722), .B1(n_740), .B2(n_745), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_726), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_L g812 ( .A1(n_733), .A2(n_687), .B(n_751), .C(n_752), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_713), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_744), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_685), .Y(n_815) );
NOR2xp33_ASAP7_75t_SL g816 ( .A(n_714), .B(n_699), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_721), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_756), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_719), .A2(n_747), .B1(n_738), .B2(n_734), .Y(n_819) );
AO21x2_ASAP7_75t_L g820 ( .A1(n_728), .A2(n_775), .B(n_690), .Y(n_820) );
INVx4_ASAP7_75t_L g821 ( .A(n_695), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_770), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_695), .B(n_790), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_749), .A2(n_694), .B(n_737), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_790), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_743), .A2(n_730), .B1(n_753), .B2(n_688), .C(n_723), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_709), .A2(n_697), .B(n_696), .C(n_725), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_781), .A2(n_682), .B1(n_736), .B2(n_793), .Y(n_828) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_692), .A2(n_693), .B(n_717), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_747), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_702), .A2(n_776), .B1(n_762), .B2(n_750), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_772), .B(n_786), .Y(n_832) );
A2O1A1Ixp33_ASAP7_75t_L g833 ( .A1(n_727), .A2(n_689), .B(n_761), .C(n_691), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_739), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_715), .A2(n_776), .B1(n_771), .B2(n_769), .Y(n_835) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_759), .A2(n_757), .B(n_724), .C(n_729), .Y(n_836) );
INVx3_ASAP7_75t_L g837 ( .A(n_771), .Y(n_837) );
OA21x2_ASAP7_75t_L g838 ( .A1(n_746), .A2(n_768), .B(n_774), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_706), .Y(n_839) );
INVx6_ASAP7_75t_L g840 ( .A(n_716), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_706), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_795), .B(n_778), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_763), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_783), .Y(n_844) );
BUFx6f_ASAP7_75t_SL g845 ( .A(n_766), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_767), .B(n_763), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_795), .B(n_784), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_767), .A2(n_755), .B1(n_758), .B2(n_763), .C(n_683), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_683), .B(n_760), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_680), .Y(n_850) );
INVx5_ASAP7_75t_L g851 ( .A(n_735), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_779), .A2(n_584), .B1(n_613), .B2(n_705), .Y(n_852) );
INVx1_ASAP7_75t_SL g853 ( .A(n_711), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_748), .B(n_672), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_684), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_707), .A2(n_699), .B1(n_672), .B2(n_543), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_711), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_788), .A2(n_676), .B(n_666), .Y(n_858) );
AOI21xp33_ASAP7_75t_L g859 ( .A1(n_779), .A2(n_789), .B(n_577), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_777), .B(n_680), .Y(n_860) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_735), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_680), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_684), .Y(n_863) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_788), .A2(n_794), .B(n_579), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_684), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_788), .A2(n_676), .B(n_666), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_680), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g868 ( .A1(n_788), .A2(n_794), .B(n_579), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_788), .A2(n_676), .B(n_666), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_777), .B(n_680), .Y(n_870) );
NOR2xp33_ASAP7_75t_SL g871 ( .A(n_714), .B(n_699), .Y(n_871) );
AO21x2_ASAP7_75t_L g872 ( .A1(n_708), .A2(n_579), .B(n_592), .Y(n_872) );
AOI21xp33_ASAP7_75t_L g873 ( .A1(n_779), .A2(n_789), .B(n_577), .Y(n_873) );
INVxp67_ASAP7_75t_L g874 ( .A(n_765), .Y(n_874) );
CKINVDCx11_ASAP7_75t_R g875 ( .A(n_685), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_735), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_788), .A2(n_676), .B(n_666), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_680), .Y(n_878) );
AO31x2_ASAP7_75t_L g879 ( .A1(n_780), .A2(n_551), .A3(n_703), .B(n_764), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_684), .Y(n_880) );
A2O1A1Ixp33_ASAP7_75t_L g881 ( .A1(n_785), .A2(n_647), .B(n_777), .C(n_613), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_777), .B(n_680), .Y(n_882) );
AO31x2_ASAP7_75t_L g883 ( .A1(n_780), .A2(n_551), .A3(n_703), .B(n_764), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_788), .A2(n_676), .B(n_666), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_684), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_777), .B(n_680), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_684), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_684), .Y(n_888) );
AO221x2_ASAP7_75t_L g889 ( .A1(n_789), .A2(n_432), .B1(n_538), .B2(n_438), .C(n_743), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_699), .A2(n_597), .B1(n_672), .B2(n_789), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_680), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_680), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g893 ( .A1(n_791), .A2(n_597), .B1(n_707), .B2(n_519), .C(n_602), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_834), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_860), .B(n_870), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_803), .B(n_852), .Y(n_896) );
OR2x6_ASAP7_75t_L g897 ( .A(n_852), .B(n_837), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_809), .B(n_811), .Y(n_898) );
AO21x2_ASAP7_75t_L g899 ( .A1(n_866), .A2(n_869), .B(n_849), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_870), .B(n_882), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_800), .B(n_855), .Y(n_901) );
AO21x2_ASAP7_75t_L g902 ( .A1(n_866), .A2(n_869), .B(n_801), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_863), .B(n_865), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_844), .Y(n_904) );
INVx3_ASAP7_75t_L g905 ( .A(n_851), .Y(n_905) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_832), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_839), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_880), .B(n_885), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_887), .B(n_888), .Y(n_909) );
OA21x2_ASAP7_75t_L g910 ( .A1(n_848), .A2(n_843), .B(n_841), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_842), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_813), .B(n_814), .Y(n_912) );
OA21x2_ASAP7_75t_L g913 ( .A1(n_848), .A2(n_868), .B(n_864), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_864), .A2(n_868), .B(n_877), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_818), .B(n_822), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_832), .B(n_882), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_842), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_875), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_886), .B(n_850), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_862), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_847), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_886), .B(n_867), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_878), .B(n_891), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_853), .B(n_857), .Y(n_924) );
INVx4_ASAP7_75t_L g925 ( .A(n_851), .Y(n_925) );
OA21x2_ASAP7_75t_L g926 ( .A1(n_858), .A2(n_884), .B(n_846), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_892), .B(n_802), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_802), .B(n_817), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_810), .A2(n_856), .B1(n_890), .B2(n_819), .C(n_893), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_816), .B(n_871), .Y(n_930) );
INVx2_ASAP7_75t_SL g931 ( .A(n_851), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_816), .B(n_871), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_808), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_889), .B(n_805), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_881), .A2(n_812), .B(n_833), .Y(n_935) );
OR2x6_ASAP7_75t_L g936 ( .A(n_854), .B(n_874), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_797), .B(n_830), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_827), .A2(n_893), .B(n_826), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_859), .B(n_873), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_835), .B(n_831), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_859), .B(n_807), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_829), .A2(n_836), .B(n_824), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_840), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_804), .B(n_826), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_879), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_883), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_828), .A2(n_876), .B1(n_799), .B2(n_796), .Y(n_947) );
INVx2_ASAP7_75t_SL g948 ( .A(n_861), .Y(n_948) );
BUFx5_ASAP7_75t_L g949 ( .A(n_845), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_804), .B(n_840), .Y(n_950) );
OR2x6_ASAP7_75t_L g951 ( .A(n_799), .B(n_876), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_883), .Y(n_952) );
INVxp33_ASAP7_75t_L g953 ( .A(n_823), .Y(n_953) );
INVx5_ASAP7_75t_L g954 ( .A(n_821), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_804), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_906), .B(n_821), .Y(n_956) );
AND2x2_ASAP7_75t_SL g957 ( .A(n_904), .B(n_798), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_944), .B(n_820), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_944), .B(n_872), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_894), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_919), .B(n_815), .Y(n_961) );
INVx5_ASAP7_75t_L g962 ( .A(n_925), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_911), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_894), .Y(n_964) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_924), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_924), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_919), .B(n_825), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_933), .Y(n_968) );
INVx5_ASAP7_75t_L g969 ( .A(n_925), .Y(n_969) );
OR2x2_ASAP7_75t_L g970 ( .A(n_896), .B(n_806), .Y(n_970) );
AND2x4_ASAP7_75t_L g971 ( .A(n_950), .B(n_806), .Y(n_971) );
INVxp33_ASAP7_75t_SL g972 ( .A(n_918), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_921), .B(n_927), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_921), .B(n_838), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_917), .B(n_913), .Y(n_975) );
OR2x2_ASAP7_75t_L g976 ( .A(n_896), .B(n_916), .Y(n_976) );
NAND2x1_ASAP7_75t_L g977 ( .A(n_897), .B(n_925), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_913), .B(n_922), .Y(n_978) );
AND2x4_ASAP7_75t_L g979 ( .A(n_950), .B(n_897), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_913), .B(n_922), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_907), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_916), .B(n_897), .Y(n_982) );
INVx4_ASAP7_75t_R g983 ( .A(n_931), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_928), .B(n_923), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_898), .B(n_901), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_903), .B(n_908), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_909), .B(n_912), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_895), .B(n_900), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_915), .B(n_897), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_940), .B(n_934), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_940), .B(n_937), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_910), .B(n_939), .Y(n_992) );
BUFx6f_ASAP7_75t_SL g993 ( .A(n_931), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_910), .B(n_939), .Y(n_994) );
INVx4_ASAP7_75t_L g995 ( .A(n_905), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_899), .B(n_941), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_978), .B(n_980), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_978), .B(n_899), .Y(n_998) );
NOR2xp33_ASAP7_75t_SL g999 ( .A(n_972), .B(n_918), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_980), .B(n_899), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_990), .B(n_929), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_996), .B(n_955), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_965), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_966), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_996), .B(n_914), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_984), .B(n_914), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_984), .B(n_914), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_985), .B(n_920), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_985), .B(n_938), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_992), .B(n_946), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_968), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_992), .B(n_946), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_976), .B(n_926), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_994), .B(n_926), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_994), .B(n_926), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_991), .B(n_902), .Y(n_1016) );
INVx2_ASAP7_75t_SL g1017 ( .A(n_983), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_960), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_983), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_960), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_964), .Y(n_1021) );
NOR2xp33_ASAP7_75t_R g1022 ( .A(n_962), .B(n_949), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_991), .B(n_902), .Y(n_1023) );
INVxp67_ASAP7_75t_SL g1024 ( .A(n_963), .Y(n_1024) );
NAND2x1p5_ASAP7_75t_L g1025 ( .A(n_962), .B(n_954), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_973), .B(n_952), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_990), .A2(n_932), .B1(n_930), .B2(n_935), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_995), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_975), .B(n_945), .Y(n_1029) );
AOI21xp33_ASAP7_75t_SL g1030 ( .A1(n_1017), .A2(n_957), .B(n_956), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_997), .B(n_959), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_997), .B(n_971), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1006), .B(n_971), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1006), .B(n_971), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1007), .B(n_971), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1007), .B(n_958), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_998), .B(n_975), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1000), .B(n_959), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1018), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1020), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1005), .B(n_979), .Y(n_1041) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_999), .B(n_947), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1021), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1009), .B(n_986), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1003), .B(n_987), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1016), .B(n_970), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1010), .B(n_981), .Y(n_1047) );
AND2x4_ASAP7_75t_L g1048 ( .A(n_1014), .B(n_1015), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1002), .B(n_989), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_1014), .B(n_974), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1012), .B(n_989), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1028), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1004), .B(n_987), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1015), .B(n_970), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_1001), .B(n_953), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_1022), .Y(n_1056) );
NAND2xp5_ASAP7_75t_SL g1057 ( .A(n_1030), .B(n_957), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1039), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1037), .B(n_1036), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1039), .Y(n_1060) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_1052), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1036), .B(n_1011), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1031), .B(n_1013), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_1031), .B(n_1013), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1040), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_1052), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1048), .B(n_1023), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_1048), .B(n_1023), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1048), .B(n_1029), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1038), .B(n_1027), .Y(n_1070) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_1055), .Y(n_1071) );
INVx1_ASAP7_75t_SL g1072 ( .A(n_1045), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1042), .B(n_1001), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1054), .B(n_1008), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1040), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1048), .B(n_1026), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1043), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1043), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1079 ( .A(n_1073), .B(n_1044), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1063), .Y(n_1080) );
OAI21xp5_ASAP7_75t_SL g1081 ( .A1(n_1057), .A2(n_1056), .B(n_1019), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1076), .B(n_1032), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1070), .B(n_1054), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1072), .B(n_1051), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1063), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1067), .B(n_1032), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1076), .B(n_1033), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1059), .B(n_1049), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1064), .B(n_1049), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_1057), .A2(n_1056), .B(n_1019), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1064), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1062), .B(n_1047), .Y(n_1092) );
INVx1_ASAP7_75t_SL g1093 ( .A(n_1061), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g1094 ( .A(n_1071), .B(n_1053), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1080), .Y(n_1095) );
NAND4xp25_ASAP7_75t_L g1096 ( .A(n_1090), .B(n_988), .C(n_937), .D(n_942), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_1093), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_1079), .A2(n_1074), .B1(n_1068), .B2(n_1075), .C(n_1077), .Y(n_1098) );
OAI211xp5_ASAP7_75t_SL g1099 ( .A1(n_1081), .A2(n_1066), .B(n_1069), .C(n_967), .Y(n_1099) );
OAI21xp5_ASAP7_75t_L g1100 ( .A1(n_1094), .A2(n_1069), .B(n_1025), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1083), .B(n_1050), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1085), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1087), .B(n_1041), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_1084), .A2(n_977), .B(n_1025), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1091), .Y(n_1105) );
A2O1A1Ixp33_ASAP7_75t_L g1106 ( .A1(n_1099), .A2(n_1082), .B(n_1092), .C(n_1089), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1098), .B(n_1088), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1100), .B(n_1086), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g1109 ( .A1(n_1096), .A2(n_969), .B(n_962), .Y(n_1109) );
INVx2_ASAP7_75t_SL g1110 ( .A(n_1097), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1095), .B(n_1105), .Y(n_1111) );
AOI32xp33_ASAP7_75t_L g1112 ( .A1(n_1103), .A2(n_1034), .A3(n_1033), .B1(n_1035), .B2(n_1041), .Y(n_1112) );
OAI211xp5_ASAP7_75t_L g1113 ( .A1(n_1104), .A2(n_1022), .B(n_962), .C(n_969), .Y(n_1113) );
A2O1A1O1Ixp25_ASAP7_75t_L g1114 ( .A1(n_1101), .A2(n_1024), .B(n_1065), .C(n_1060), .D(n_1058), .Y(n_1114) );
OR5x1_ASAP7_75t_L g1115 ( .A(n_1113), .B(n_1102), .C(n_936), .D(n_993), .E(n_949), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1110), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1107), .B(n_1046), .Y(n_1117) );
NAND4xp25_ASAP7_75t_L g1118 ( .A(n_1109), .B(n_961), .C(n_995), .D(n_982), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1106), .B(n_1078), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1117), .B(n_1111), .Y(n_1120) );
OR4x2_ASAP7_75t_L g1121 ( .A(n_1115), .B(n_1114), .C(n_1112), .D(n_1108), .Y(n_1121) );
OR2x2_ASAP7_75t_SL g1122 ( .A(n_1116), .B(n_1109), .Y(n_1122) );
NOR2x1_ASAP7_75t_L g1123 ( .A(n_1118), .B(n_951), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1122), .Y(n_1124) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1120), .Y(n_1125) );
XNOR2x1_ASAP7_75t_L g1126 ( .A(n_1123), .B(n_1119), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1121), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_1125), .Y(n_1128) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_1124), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_1128), .A2(n_1127), .B1(n_1126), .B2(n_1129), .Y(n_1130) );
OAI22xp5_ASAP7_75t_SL g1131 ( .A1(n_1130), .A2(n_951), .B1(n_954), .B2(n_948), .Y(n_1131) );
XNOR2xp5_ASAP7_75t_L g1132 ( .A(n_1131), .B(n_951), .Y(n_1132) );
XNOR2xp5_ASAP7_75t_L g1133 ( .A(n_1132), .B(n_951), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1134 ( .A1(n_1133), .A2(n_954), .B(n_943), .Y(n_1134) );
endmodule