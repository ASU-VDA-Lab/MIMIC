module fake_jpeg_31747_n_269 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_22),
.Y(n_82)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_28),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_27),
.C(n_22),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_61),
.B(n_70),
.Y(n_121)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_39),
.B1(n_38),
.B2(n_30),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_19),
.B1(n_25),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_38),
.B1(n_30),
.B2(n_34),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_73),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_13),
.Y(n_100)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_35),
.B1(n_25),
.B2(n_29),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_46),
.B1(n_52),
.B2(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_2),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_35),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_40),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_100),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_96),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_24),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_116),
.C(n_84),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_123),
.B1(n_85),
.B2(n_62),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_84),
.B1(n_79),
.B2(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_52),
.Y(n_110)
);

OR2x4_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_44),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_8),
.B(n_9),
.Y(n_151)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_44),
.B(n_56),
.C(n_43),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_87),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_47),
.C(n_1),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_15),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_124),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_75),
.B1(n_67),
.B2(n_86),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_59),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_7),
.CI(n_8),
.CON(n_125),
.SN(n_125)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_134),
.B1(n_118),
.B2(n_119),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_118),
.A2(n_75),
.B1(n_86),
.B2(n_67),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_153),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_60),
.B1(n_85),
.B2(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_141),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_96),
.B1(n_114),
.B2(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_16),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_87),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_149),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_7),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_95),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_125),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_110),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_124),
.C(n_116),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_135),
.B1(n_148),
.B2(n_128),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_157),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_122),
.B1(n_112),
.B2(n_107),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_154),
.B(n_166),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_150),
.C(n_136),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_175),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_124),
.B(n_125),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_135),
.B(n_128),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_180),
.B1(n_151),
.B2(n_132),
.C(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_100),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_177),
.C(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_102),
.B1(n_109),
.B2(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_134),
.Y(n_188)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_96),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_131),
.B(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_103),
.A3(n_115),
.B1(n_12),
.B2(n_10),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_186),
.C(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_145),
.B(n_144),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_195),
.B(n_162),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_200),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_201),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_147),
.B(n_148),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_166),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_129),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_129),
.C1(n_113),
.C2(n_99),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_207),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_212),
.Y(n_225)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_167),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_163),
.B(n_156),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_188),
.B(n_176),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_171),
.B1(n_194),
.B2(n_163),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_165),
.Y(n_219)
);

NOR4xp25_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_165),
.C(n_182),
.D(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_181),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_226),
.C(n_227),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_187),
.C(n_186),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_190),
.C(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_197),
.C(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_205),
.C(n_216),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_193),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_208),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_205),
.B1(n_172),
.B2(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_222),
.C(n_232),
.Y(n_239)
);

OAI22x1_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_215),
.B1(n_206),
.B2(n_208),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_240),
.A2(n_215),
.B1(n_180),
.B2(n_218),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_217),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_231),
.B(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_233),
.C(n_168),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_202),
.B1(n_238),
.B2(n_240),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_242),
.A3(n_207),
.B1(n_218),
.B2(n_233),
.C1(n_194),
.C2(n_174),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_159),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_256),
.A2(n_173),
.B1(n_129),
.B2(n_10),
.Y(n_261)
);

AOI31xp33_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_174),
.A3(n_178),
.B(n_159),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_173),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_254),
.A2(n_244),
.B(n_246),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.C(n_173),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_263),
.A2(n_259),
.B(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_266),
.B(n_267),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_263),
.Y(n_269)
);


endmodule