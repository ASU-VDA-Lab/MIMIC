module real_aes_215_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_246;
wire n_412;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_294;
wire n_393;
wire n_258;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_0), .A2(n_219), .B1(n_444), .B2(n_446), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_1), .A2(n_189), .B1(n_419), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_2), .A2(n_82), .B1(n_243), .B2(n_261), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_3), .A2(n_187), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_4), .A2(n_117), .B1(n_329), .B2(n_330), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_5), .A2(n_72), .B1(n_220), .B2(n_365), .C1(n_366), .C2(n_367), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_6), .A2(n_77), .B1(n_486), .B2(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_7), .A2(n_58), .B1(n_326), .B2(n_327), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_8), .A2(n_137), .B1(n_341), .B2(n_342), .Y(n_358) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_9), .A2(n_170), .B1(n_248), .B2(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g581 ( .A(n_9), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_10), .A2(n_142), .B1(n_261), .B2(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_11), .A2(n_66), .B1(n_386), .B2(n_531), .Y(n_594) );
XOR2x2_ASAP7_75t_L g401 ( .A(n_12), .B(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_13), .A2(n_99), .B1(n_348), .B2(n_362), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_14), .A2(n_169), .B1(n_332), .B2(n_333), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_15), .A2(n_84), .B1(n_341), .B2(n_342), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_16), .A2(n_96), .B1(n_315), .B2(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_17), .A2(n_35), .B1(n_326), .B2(n_327), .Y(n_465) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_18), .A2(n_56), .B1(n_248), .B2(n_249), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_18), .B(n_580), .Y(n_579) );
OA22x2_ASAP7_75t_L g538 ( .A1(n_19), .A2(n_539), .B1(n_553), .B2(n_554), .Y(n_538) );
INVx1_ASAP7_75t_L g553 ( .A(n_19), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_20), .A2(n_54), .B1(n_276), .B2(n_496), .Y(n_495) );
AOI22xp5_ASAP7_75t_SL g491 ( .A1(n_21), .A2(n_203), .B1(n_266), .B2(n_420), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_22), .A2(n_129), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_23), .A2(n_112), .B1(n_398), .B2(n_399), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_24), .A2(n_111), .B1(n_326), .B2(n_327), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_25), .A2(n_125), .B1(n_292), .B2(n_296), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_26), .A2(n_37), .B1(n_345), .B2(n_360), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_27), .A2(n_223), .B(n_232), .C(n_583), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_28), .A2(n_164), .B1(n_300), .B2(n_303), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_29), .A2(n_198), .B1(n_305), .B2(n_531), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_30), .B(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_31), .A2(n_155), .B1(n_315), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_32), .A2(n_214), .B1(n_276), .B2(n_417), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_33), .A2(n_95), .B1(n_302), .B2(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_34), .A2(n_196), .B1(n_365), .B2(n_366), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_36), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_38), .A2(n_197), .B1(n_332), .B2(n_333), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_39), .B(n_285), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_40), .A2(n_182), .B1(n_276), .B2(n_280), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_41), .A2(n_45), .B1(n_261), .B2(n_395), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_42), .A2(n_156), .B1(n_341), .B2(n_342), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_43), .A2(n_181), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_44), .A2(n_216), .B1(n_341), .B2(n_342), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_46), .A2(n_151), .B1(n_548), .B2(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_47), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_48), .A2(n_148), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_49), .A2(n_136), .B1(n_329), .B2(n_330), .Y(n_566) );
OAI22x1_ASAP7_75t_SL g504 ( .A1(n_50), .A2(n_505), .B1(n_533), .B2(n_534), .Y(n_504) );
INVx1_ASAP7_75t_L g533 ( .A(n_50), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_51), .A2(n_85), .B1(n_338), .B2(n_339), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_52), .A2(n_186), .B1(n_524), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_53), .A2(n_179), .B1(n_510), .B2(n_512), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_55), .A2(n_57), .B1(n_411), .B2(n_412), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_59), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_60), .A2(n_175), .B1(n_329), .B2(n_330), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_61), .A2(n_128), .B1(n_190), .B2(n_261), .C1(n_395), .C2(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_62), .A2(n_162), .B1(n_348), .B2(n_362), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_63), .A2(n_118), .B1(n_419), .B2(n_420), .Y(n_418) );
INVx3_ASAP7_75t_L g248 ( .A(n_64), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_65), .B(n_335), .Y(n_334) );
XNOR2x2_ASAP7_75t_L g322 ( .A(n_67), .B(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_68), .A2(n_208), .B1(n_296), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_69), .A2(n_193), .B1(n_332), .B2(n_333), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_70), .A2(n_127), .B1(n_338), .B2(n_339), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_71), .A2(n_88), .B1(n_303), .B2(n_314), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_73), .A2(n_105), .B1(n_307), .B2(n_310), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_74), .B(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_75), .A2(n_126), .B1(n_303), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_97), .B1(n_310), .B2(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_78), .A2(n_102), .B1(n_419), .B2(n_543), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_79), .A2(n_87), .B1(n_315), .B2(n_339), .Y(n_616) );
INVx1_ASAP7_75t_SL g256 ( .A(n_80), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_80), .B(n_104), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_81), .A2(n_98), .B1(n_329), .B2(n_330), .Y(n_621) );
INVx2_ASAP7_75t_L g229 ( .A(n_83), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_86), .A2(n_138), .B1(n_339), .B2(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_89), .B(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_90), .A2(n_121), .B1(n_276), .B2(n_399), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_91), .A2(n_202), .B1(n_261), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_92), .A2(n_135), .B1(n_529), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_93), .A2(n_194), .B1(n_296), .B2(n_314), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_94), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_100), .A2(n_171), .B1(n_326), .B2(n_327), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_101), .A2(n_192), .B1(n_315), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_103), .A2(n_140), .B1(n_308), .B2(n_378), .Y(n_549) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_104), .A2(n_176), .B1(n_248), .B2(n_260), .Y(n_259) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_106), .A2(n_211), .B1(n_261), .B2(n_422), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_107), .A2(n_161), .B1(n_261), .B2(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_108), .A2(n_166), .B1(n_338), .B2(n_339), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_109), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_110), .A2(n_152), .B1(n_292), .B2(n_405), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_113), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_114), .A2(n_150), .B1(n_386), .B2(n_531), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_115), .A2(n_191), .B1(n_276), .B2(n_280), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_116), .A2(n_213), .B1(n_307), .B2(n_310), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_119), .A2(n_159), .B1(n_300), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_120), .A2(n_215), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g257 ( .A(n_122), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_123), .A2(n_153), .B1(n_266), .B2(n_270), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_124), .B(n_456), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_130), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_131), .A2(n_144), .B1(n_347), .B2(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_132), .B(n_367), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_133), .A2(n_204), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_134), .A2(n_141), .B1(n_344), .B2(n_345), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_139), .A2(n_158), .B1(n_438), .B2(n_439), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_143), .B(n_335), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_145), .A2(n_218), .B1(n_338), .B2(n_339), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_146), .A2(n_206), .B1(n_344), .B2(n_345), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g312 ( .A1(n_147), .A2(n_178), .B1(n_313), .B2(n_315), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_149), .A2(n_180), .B1(n_307), .B2(n_310), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_154), .A2(n_585), .B1(n_606), .B2(n_607), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_154), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_157), .A2(n_163), .B1(n_266), .B2(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_160), .A2(n_217), .B1(n_441), .B2(n_442), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_165), .B(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_167), .A2(n_210), .B1(n_307), .B2(n_310), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_168), .A2(n_177), .B1(n_378), .B2(n_380), .Y(n_377) );
XNOR2x1_ASAP7_75t_L g434 ( .A(n_172), .B(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_173), .A2(n_184), .B1(n_314), .B2(n_382), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_174), .A2(n_221), .B1(n_415), .B2(n_417), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_183), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_185), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g577 ( .A(n_185), .Y(n_577) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
AND2x2_ASAP7_75t_R g609 ( .A(n_188), .B(n_577), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_195), .A2(n_205), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_199), .A2(n_209), .B1(n_395), .B2(n_493), .Y(n_492) );
INVxp67_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_201), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_207), .B(n_261), .Y(n_602) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_212), .A2(n_240), .B1(n_318), .B2(n_319), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_212), .Y(n_318) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2x1_ASAP7_75t_R g224 ( .A(n_225), .B(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g626 ( .A(n_225), .B(n_228), .Y(n_626) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_226), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_500), .B1(n_572), .B2(n_573), .C(n_574), .Y(n_232) );
INVx1_ASAP7_75t_L g572 ( .A(n_233), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_430), .B2(n_432), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_352), .B2(n_429), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_320), .B1(n_349), .B2(n_350), .Y(n_237) );
INVx1_ASAP7_75t_L g349 ( .A(n_238), .Y(n_349) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_SL g319 ( .A(n_240), .Y(n_319) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_241), .B(n_290), .Y(n_240) );
NAND4xp25_ASAP7_75t_L g241 ( .A(n_242), .B(n_265), .C(n_275), .D(n_284), .Y(n_241) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g601 ( .A(n_244), .Y(n_601) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g395 ( .A(n_245), .Y(n_395) );
BUFx5_ASAP7_75t_L g422 ( .A(n_245), .Y(n_422) );
BUFx3_ASAP7_75t_L g623 ( .A(n_245), .Y(n_623) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
AND2x4_ASAP7_75t_L g267 ( .A(n_246), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g314 ( .A(n_246), .B(n_295), .Y(n_314) );
AND2x2_ASAP7_75t_L g329 ( .A(n_246), .B(n_268), .Y(n_329) );
AND2x4_ASAP7_75t_L g332 ( .A(n_246), .B(n_253), .Y(n_332) );
AND2x2_ASAP7_75t_L g348 ( .A(n_246), .B(n_295), .Y(n_348) );
AND2x2_ASAP7_75t_L g366 ( .A(n_246), .B(n_268), .Y(n_366) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g263 ( .A(n_247), .B(n_251), .Y(n_263) );
INVx1_ASAP7_75t_L g279 ( .A(n_247), .Y(n_279) );
INVx1_ASAP7_75t_L g289 ( .A(n_247), .Y(n_289) );
INVx2_ASAP7_75t_L g249 ( .A(n_248), .Y(n_249) );
INVx1_ASAP7_75t_L g252 ( .A(n_248), .Y(n_252) );
OAI22x1_ASAP7_75t_L g254 ( .A1(n_248), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_248), .Y(n_255) );
INVx1_ASAP7_75t_L g260 ( .A(n_248), .Y(n_260) );
INVxp67_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
AND2x4_ASAP7_75t_L g288 ( .A(n_250), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g277 ( .A(n_253), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g305 ( .A(n_253), .B(n_288), .Y(n_305) );
AND2x4_ASAP7_75t_L g326 ( .A(n_253), .B(n_278), .Y(n_326) );
AND2x2_ASAP7_75t_L g341 ( .A(n_253), .B(n_288), .Y(n_341) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_258), .Y(n_253) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_254), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_254), .Y(n_269) );
AND2x2_ASAP7_75t_L g274 ( .A(n_254), .B(n_259), .Y(n_274) );
AND2x4_ASAP7_75t_L g295 ( .A(n_258), .B(n_269), .Y(n_295) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g268 ( .A(n_259), .B(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g309 ( .A(n_259), .Y(n_309) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g494 ( .A(n_262), .Y(n_494) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x4_ASAP7_75t_L g302 ( .A(n_263), .B(n_295), .Y(n_302) );
AND2x4_ASAP7_75t_L g308 ( .A(n_263), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_263), .B(n_264), .Y(n_333) );
AND2x4_ASAP7_75t_L g342 ( .A(n_263), .B(n_295), .Y(n_342) );
AND2x4_ASAP7_75t_L g345 ( .A(n_263), .B(n_309), .Y(n_345) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g419 ( .A(n_267), .Y(n_419) );
AND2x2_ASAP7_75t_L g298 ( .A(n_268), .B(n_288), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_268), .B(n_278), .Y(n_311) );
AND2x6_ASAP7_75t_L g338 ( .A(n_268), .B(n_288), .Y(n_338) );
AND2x2_ASAP7_75t_L g344 ( .A(n_268), .B(n_278), .Y(n_344) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_268), .B(n_278), .Y(n_360) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g420 ( .A(n_271), .Y(n_420) );
INVx2_ASAP7_75t_SL g452 ( .A(n_271), .Y(n_452) );
INVx2_ASAP7_75t_L g512 ( .A(n_271), .Y(n_512) );
INVx2_ASAP7_75t_L g543 ( .A(n_271), .Y(n_543) );
INVx6_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g330 ( .A(n_273), .B(n_274), .Y(n_330) );
AND2x2_ASAP7_75t_L g365 ( .A(n_273), .B(n_274), .Y(n_365) );
AND2x4_ASAP7_75t_L g281 ( .A(n_274), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g287 ( .A(n_274), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g327 ( .A(n_274), .B(n_282), .Y(n_327) );
AND2x4_ASAP7_75t_L g367 ( .A(n_274), .B(n_288), .Y(n_367) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_277), .Y(n_398) );
INVx3_ASAP7_75t_L g416 ( .A(n_277), .Y(n_416) );
AND2x4_ASAP7_75t_L g294 ( .A(n_278), .B(n_295), .Y(n_294) );
AND2x6_ASAP7_75t_L g339 ( .A(n_278), .B(n_295), .Y(n_339) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
BUFx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_SL g399 ( .A(n_281), .Y(n_399) );
BUFx4f_ASAP7_75t_L g417 ( .A(n_281), .Y(n_417) );
INVx1_ASAP7_75t_L g497 ( .A(n_281), .Y(n_497) );
INVx2_ASAP7_75t_L g520 ( .A(n_281), .Y(n_520) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx4_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx4_ASAP7_75t_SL g335 ( .A(n_286), .Y(n_335) );
INVx3_ASAP7_75t_L g424 ( .A(n_286), .Y(n_424) );
INVx3_ASAP7_75t_SL g456 ( .A(n_286), .Y(n_456) );
INVx6_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g317 ( .A(n_288), .B(n_295), .Y(n_317) );
AND2x2_ASAP7_75t_L g362 ( .A(n_288), .B(n_295), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g290 ( .A(n_291), .B(n_299), .C(n_306), .D(n_312), .Y(n_290) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g442 ( .A(n_293), .Y(n_442) );
INVx2_ASAP7_75t_L g486 ( .A(n_293), .Y(n_486) );
INVx2_ASAP7_75t_L g551 ( .A(n_293), .Y(n_551) );
INVx2_ASAP7_75t_SL g596 ( .A(n_293), .Y(n_596) );
INVx8_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_SL g441 ( .A(n_297), .Y(n_441) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g405 ( .A(n_298), .Y(n_405) );
BUFx2_ASAP7_75t_L g524 ( .A(n_298), .Y(n_524) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_SL g408 ( .A(n_301), .Y(n_408) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g488 ( .A(n_302), .Y(n_488) );
BUFx3_ASAP7_75t_L g531 ( .A(n_302), .Y(n_531) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g407 ( .A(n_304), .Y(n_407) );
INVx2_ASAP7_75t_L g438 ( .A(n_304), .Y(n_438) );
INVx6_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g386 ( .A(n_305), .Y(n_386) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g380 ( .A(n_308), .Y(n_380) );
BUFx2_ASAP7_75t_L g446 ( .A(n_308), .Y(n_446) );
INVx5_ASAP7_75t_SL g482 ( .A(n_308), .Y(n_482) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g379 ( .A(n_311), .Y(n_379) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g389 ( .A(n_314), .Y(n_389) );
BUFx3_ASAP7_75t_L g439 ( .A(n_314), .Y(n_439) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_314), .Y(n_484) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_314), .Y(n_548) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx4_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
INVx2_ASAP7_75t_SL g411 ( .A(n_316), .Y(n_411) );
INVx2_ASAP7_75t_SL g448 ( .A(n_316), .Y(n_448) );
INVx2_ASAP7_75t_L g529 ( .A(n_316), .Y(n_529) );
INVx3_ASAP7_75t_SL g560 ( .A(n_316), .Y(n_560) );
INVx8_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g351 ( .A(n_322), .Y(n_351) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_336), .Y(n_323) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .C(n_331), .D(n_334), .Y(n_324) );
BUFx2_ASAP7_75t_L g508 ( .A(n_335), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .C(n_343), .D(n_346), .Y(n_336) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g429 ( .A(n_352), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_371), .B1(n_427), .B2(n_428), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
XNOR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_370), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_363), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .C(n_359), .D(n_361), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_368), .C(n_369), .Y(n_363) );
INVx2_ASAP7_75t_SL g392 ( .A(n_367), .Y(n_392) );
BUFx2_ASAP7_75t_L g568 ( .A(n_367), .Y(n_568) );
INVx2_ASAP7_75t_L g428 ( .A(n_371), .Y(n_428) );
OA22x2_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_401), .B1(n_425), .B2(n_426), .Y(n_371) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_372), .Y(n_426) );
XNOR2x1_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_375), .B(n_390), .Y(n_374) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_378), .Y(n_526) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
INVx1_ASAP7_75t_L g591 ( .A(n_379), .Y(n_591) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_396), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B(n_394), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_392), .A2(n_599), .B(n_600), .C(n_602), .Y(n_598) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_395), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
BUFx6f_ASAP7_75t_SL g518 ( .A(n_398), .Y(n_518) );
INVx1_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_403), .B(n_413), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .C(n_409), .D(n_410), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .C(n_421), .D(n_423), .Y(n_413) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g511 ( .A(n_419), .Y(n_511) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_457), .B2(n_458), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_449), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .C(n_443), .D(n_447), .Y(n_436) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .C(n_453), .D(n_454), .Y(n_449) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_477), .B2(n_499), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_476), .Y(n_460) );
NAND2x1_ASAP7_75t_SL g461 ( .A(n_462), .B(n_469), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_SL g499 ( .A(n_477), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_498), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .C(n_485), .D(n_487), .Y(n_479) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g527 ( .A(n_482), .Y(n_527) );
INVx2_ASAP7_75t_L g592 ( .A(n_482), .Y(n_592) );
NAND4xp25_ASAP7_75t_SL g489 ( .A(n_490), .B(n_491), .C(n_492), .D(n_495), .Y(n_489) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g516 ( .A(n_494), .Y(n_516) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_535), .B2(n_536), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g534 ( .A(n_505), .Y(n_534) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_521), .Y(n_505) );
NAND4xp25_ASAP7_75t_SL g506 ( .A(n_507), .B(n_509), .C(n_513), .D(n_517), .Y(n_506) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .C(n_528), .D(n_532), .Y(n_521) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AO22x1_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_555), .B1(n_570), .B2(n_571), .Y(n_537) );
INVx1_ASAP7_75t_L g570 ( .A(n_538), .Y(n_570) );
INVx1_ASAP7_75t_L g554 ( .A(n_539), .Y(n_554) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .C(n_544), .D(n_545), .Y(n_540) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .C(n_550), .D(n_552), .Y(n_546) );
INVx1_ASAP7_75t_SL g571 ( .A(n_555), .Y(n_571) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_564), .D(n_567), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_576), .B(n_579), .Y(n_625) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_608), .B1(n_610), .B2(n_612), .C1(n_625), .C2(n_626), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_585), .Y(n_607) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_597), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_619), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .C(n_617), .D(n_618), .Y(n_614) );
NAND4xp25_ASAP7_75t_SL g619 ( .A(n_620), .B(n_621), .C(n_622), .D(n_624), .Y(n_619) );
endmodule