module fake_jpeg_15124_n_354 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_70),
.B1(n_32),
.B2(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_1),
.B(n_37),
.Y(n_99)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_71),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_38),
.B1(n_30),
.B2(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_77),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_12),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_25),
.B1(n_20),
.B2(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_111),
.B1(n_18),
.B2(n_38),
.Y(n_116)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_25),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_95),
.Y(n_125)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_94),
.Y(n_132)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_19),
.B1(n_34),
.B2(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_112),
.B1(n_114),
.B2(n_29),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_102),
.Y(n_137)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_1),
.B(n_2),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_104),
.Y(n_144)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_20),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_18),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_26),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_52),
.B1(n_42),
.B2(n_49),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_115),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_126),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_89),
.B1(n_93),
.B2(n_4),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_29),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_47),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_29),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_128),
.B(n_46),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_29),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_50),
.B1(n_52),
.B2(n_49),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_84),
.B1(n_92),
.B2(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_142),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_111),
.B(n_87),
.C(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_21),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_26),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_112),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_153),
.B(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_137),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_47),
.A3(n_46),
.B1(n_43),
.B2(n_27),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_163),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_128),
.B1(n_127),
.B2(n_138),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_103),
.B1(n_115),
.B2(n_40),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_160),
.B1(n_174),
.B2(n_118),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_129),
.Y(n_184)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_87),
.C(n_108),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_120),
.C(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_146),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

BUFx24_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_43),
.B1(n_27),
.B2(n_40),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_170),
.B1(n_138),
.B2(n_133),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_119),
.A2(n_36),
.B1(n_79),
.B2(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_26),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_184),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_119),
.B(n_126),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_190),
.B(n_192),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_153),
.B1(n_143),
.B2(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_198),
.B1(n_134),
.B2(n_26),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_188),
.A2(n_36),
.B1(n_21),
.B2(n_48),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_119),
.B(n_128),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_149),
.B(n_162),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_170),
.C(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_200),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_125),
.B1(n_127),
.B2(n_131),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_154),
.A2(n_140),
.B1(n_134),
.B2(n_122),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_163),
.B1(n_153),
.B2(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_118),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_204),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_202),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_216),
.C(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_204),
.B1(n_192),
.B2(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_230),
.B1(n_235),
.B2(n_176),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_153),
.B(n_137),
.C(n_165),
.D(n_141),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_219),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_224),
.B1(n_226),
.B2(n_234),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_124),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_145),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_26),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_22),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_22),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_36),
.B1(n_22),
.B2(n_21),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_233),
.Y(n_240)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_204),
.B1(n_189),
.B2(n_180),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_248),
.B1(n_261),
.B2(n_241),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_247),
.C(n_222),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_175),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_214),
.B(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_188),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_210),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_180),
.B1(n_197),
.B2(n_191),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_191),
.B1(n_199),
.B2(n_7),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_216),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_211),
.B1(n_230),
.B2(n_235),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_283),
.B1(n_245),
.B2(n_247),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_281),
.C(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_199),
.C(n_48),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_240),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_2),
.B1(n_5),
.B2(n_10),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_300),
.C(n_301),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_294),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_303),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_248),
.B1(n_256),
.B2(n_238),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_302),
.B1(n_271),
.B2(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_260),
.C(n_261),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_257),
.C(n_250),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_242),
.B1(n_248),
.B2(n_12),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_271),
.A2(n_268),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_278),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_306),
.B(n_315),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_316),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_281),
.B1(n_284),
.B2(n_12),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_300),
.B1(n_291),
.B2(n_14),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_10),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_11),
.C(n_13),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_296),
.C(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_287),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_322),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_287),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_289),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_305),
.C(n_304),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_303),
.B(n_293),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_308),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_329),
.B1(n_312),
.B2(n_314),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_317),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_334),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_323),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_336),
.Y(n_340)
);

NOR2x1_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_337),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_15),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_15),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_326),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_343),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_331),
.A2(n_319),
.B1(n_324),
.B2(n_15),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_17),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_345),
.B(n_346),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_334),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_347),
.B(n_339),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_350),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_341),
.Y(n_352)
);

O2A1O1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_342),
.B(n_348),
.C(n_340),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_333),
.Y(n_354)
);


endmodule