module fake_jpeg_10811_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_42),
.B(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_18),
.B(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_0),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_22),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_32),
.B1(n_38),
.B2(n_35),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_29),
.B1(n_20),
.B2(n_45),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_28),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_87),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_16),
.B1(n_38),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_87),
.B1(n_41),
.B2(n_52),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_25),
.CON(n_87),
.SN(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_25),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_107),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_100),
.B1(n_105),
.B2(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_33),
.B1(n_39),
.B2(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_57),
.B1(n_55),
.B2(n_53),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_115),
.B1(n_121),
.B2(n_81),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_24),
.B1(n_39),
.B2(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_34),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_113),
.C(n_119),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_46),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_29),
.B1(n_24),
.B2(n_20),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_34),
.B(n_2),
.C(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_34),
.C(n_2),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_1),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_4),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_1),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_92),
.B1(n_94),
.B2(n_81),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_122),
.B1(n_120),
.B2(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_121),
.B1(n_106),
.B2(n_111),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_67),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_143),
.B(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_73),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_86),
.B(n_70),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_4),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_120),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_71),
.Y(n_146)
);

XNOR2x2_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_71),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_135),
.B1(n_149),
.B2(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_113),
.C(n_117),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.C(n_165),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_113),
.C(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_163),
.Y(n_171)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_118),
.B(n_121),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_121),
.C(n_86),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_9),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_138),
.A3(n_146),
.B1(n_127),
.B2(n_142),
.C1(n_148),
.C2(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_156),
.B1(n_168),
.B2(n_155),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_126),
.CI(n_130),
.CON(n_180),
.SN(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_130),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_147),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_169),
.A2(n_147),
.B1(n_133),
.B2(n_128),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_165),
.B1(n_169),
.B2(n_152),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_193),
.B1(n_180),
.B2(n_174),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_160),
.B1(n_158),
.B2(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_185),
.B(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_157),
.B(n_153),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_181),
.C(n_176),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_179),
.B1(n_170),
.B2(n_176),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_199),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_180),
.C(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_190),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_175),
.B1(n_183),
.B2(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_206),
.B1(n_187),
.B2(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_214),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_174),
.B1(n_197),
.B2(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_201),
.C(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_173),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_207),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_220),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_218),
.C(n_204),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_209),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_227),
.A2(n_175),
.B(n_225),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_224),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_206),
.Y(n_232)
);


endmodule