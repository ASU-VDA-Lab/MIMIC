module fake_netlist_1_6162_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
AND2x6_ASAP7_75t_L g5 ( .A(n_0), .B(n_1), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
NAND2x1p5_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_6), .B(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
AO22x1_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_5), .B1(n_9), .B2(n_2), .Y(n_12) );
OAI211xp5_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_0), .B(n_2), .C(n_6), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_2), .B(n_12), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
endmodule