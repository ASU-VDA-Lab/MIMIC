module fake_jpeg_8538_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_10),
.B(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_23),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_23),
.B1(n_22),
.B2(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_30),
.B1(n_16),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_64),
.B1(n_65),
.B2(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_30),
.B1(n_25),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_62),
.B1(n_27),
.B2(n_19),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_18),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_35),
.B(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_30),
.B1(n_20),
.B2(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_36),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_35),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_62),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_75),
.B1(n_59),
.B2(n_22),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_33),
.B(n_60),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_33),
.B1(n_32),
.B2(n_42),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_63),
.B1(n_58),
.B2(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_15),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_36),
.B1(n_22),
.B2(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_50),
.B1(n_60),
.B2(n_43),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_11),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_94),
.B1(n_109),
.B2(n_78),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_103),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_60),
.B1(n_43),
.B2(n_56),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_35),
.B(n_32),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_75),
.B(n_87),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_32),
.C(n_33),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_75),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_111),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_75),
.B(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_33),
.Y(n_149)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_114),
.B(n_120),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_122),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_133),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_107),
.B1(n_104),
.B2(n_77),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_75),
.B1(n_71),
.B2(n_77),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_92),
.B1(n_133),
.B2(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_78),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_18),
.B(n_17),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_132),
.B(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_105),
.B(n_97),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_139),
.B(n_142),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_102),
.B(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_156),
.B1(n_126),
.B2(n_129),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_95),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_88),
.B1(n_94),
.B2(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_153),
.C(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_33),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_127),
.B1(n_93),
.B2(n_25),
.Y(n_189)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_171),
.C(n_170),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_124),
.A3(n_118),
.B1(n_116),
.B2(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_128),
.B1(n_123),
.B2(n_121),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_170),
.A2(n_172),
.B1(n_146),
.B2(n_144),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_125),
.B1(n_120),
.B2(n_115),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_107),
.B1(n_93),
.B2(n_47),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_174),
.B1(n_141),
.B2(n_140),
.Y(n_178)
);

NOR2x1p5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_17),
.Y(n_174)
);

BUFx4f_ASAP7_75t_SL g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_182),
.B(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_68),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_191),
.C(n_192),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_144),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_146),
.B(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_189),
.B1(n_161),
.B2(n_174),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_48),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_127),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_48),
.C(n_47),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_173),
.B1(n_160),
.B2(n_177),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_205),
.B(n_206),
.Y(n_219)
);

AO221x1_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_179),
.B1(n_176),
.B2(n_167),
.C(n_185),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_9),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_166),
.B(n_15),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_207),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_205)
);

INVxp33_ASAP7_75t_SL g206 ( 
.A(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_26),
.B1(n_25),
.B2(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_192),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_191),
.C(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_18),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_8),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_26),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_197),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_8),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_195),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_202),
.B1(n_205),
.B2(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_228),
.B1(n_220),
.B2(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_100),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_208),
.B1(n_209),
.B2(n_207),
.Y(n_228)
);

AOI221xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_12),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_10),
.B(n_4),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_4),
.B(n_5),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_230),
.B(n_210),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_235),
.B(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_211),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_226),
.B1(n_5),
.B2(n_6),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_4),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_226),
.B(n_5),
.C(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_246),
.A3(n_0),
.B1(n_13),
.B2(n_14),
.C1(n_242),
.C2(n_230),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_225),
.B(n_9),
.C(n_13),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_243),
.C(n_14),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_249),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_247),
.Y(n_251)
);


endmodule