module fake_netlist_5_2394_n_452 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_452);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_452;

wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_444;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_397;
wire n_155;
wire n_423;
wire n_284;
wire n_245;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_314;
wire n_368;
wire n_247;
wire n_433;
wire n_321;
wire n_292;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_355;
wire n_336;
wire n_430;
wire n_337;
wire n_313;
wire n_216;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_213;
wire n_342;
wire n_361;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_239;
wire n_420;
wire n_310;
wire n_358;
wire n_362;
wire n_332;
wire n_170;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_441;
wire n_450;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_25),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_47),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_31),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_18),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_10),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_30),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

INVxp33_ASAP7_75t_SL g167 ( 
.A(n_54),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_36),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_37),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_32),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_86),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_33),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_55),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_92),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_9),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_44),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_43),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_130),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_15),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_79),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_72),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_57),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_91),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_41),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_76),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_104),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_120),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_140),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_66),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_56),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_45),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_20),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_98),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_97),
.Y(n_231)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_53),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_49),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_117),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_121),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_71),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_105),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_39),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_42),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_17),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_61),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_115),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_110),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_84),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_65),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_19),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_63),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_138),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_67),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_75),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_23),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_14),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_116),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_101),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_88),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_127),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_119),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_136),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_196),
.B(n_1),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_153),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_159),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_212),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_224),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_R g280 ( 
.A(n_237),
.B(n_2),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_201),
.B(n_5),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_210),
.B(n_8),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_154),
.B(n_177),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_151),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_228),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_152),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_240),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_245),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_216),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_156),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_R g297 ( 
.A(n_243),
.B(n_12),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_162),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_267),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_268),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_233),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_167),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_157),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_163),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_169),
.B(n_16),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_R g311 ( 
.A(n_186),
.B(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_161),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_180),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_164),
.B(n_168),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_255),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_190),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_165),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_R g318 ( 
.A(n_171),
.B(n_21),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

AND3x2_ASAP7_75t_L g320 ( 
.A(n_150),
.B(n_22),
.C(n_27),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_251),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_172),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_175),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_176),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_187),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_188),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_195),
.Y(n_330)
);

NAND2x1p5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_178),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_257),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

AO22x2_ASAP7_75t_L g337 ( 
.A1(n_272),
.A2(n_199),
.B1(n_265),
.B2(n_264),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

OAI221xp5_ASAP7_75t_L g339 ( 
.A1(n_271),
.A2(n_277),
.B1(n_304),
.B2(n_308),
.C(n_317),
.Y(n_339)
);

AND2x6_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_179),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_191),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

OR2x2_ASAP7_75t_SL g343 ( 
.A(n_300),
.B(n_181),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_200),
.B1(n_262),
.B2(n_261),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_197),
.B1(n_260),
.B2(n_258),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_276),
.B(n_158),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_194),
.B1(n_256),
.B2(n_253),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_182),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_274),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_160),
.Y(n_355)
);

NAND2x1p5_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_183),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_248),
.B1(n_221),
.B2(n_219),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_289),
.B(n_193),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_322),
.B(n_220),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_355),
.A2(n_283),
.B(n_302),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_SL g365 ( 
.A(n_327),
.B(n_313),
.C(n_309),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_336),
.A2(n_323),
.B(n_269),
.C(n_254),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_359),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_343),
.B1(n_345),
.B2(n_348),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_360),
.A2(n_326),
.B1(n_330),
.B2(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_342),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_292),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_351),
.A2(n_202),
.B(n_185),
.C(n_174),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_294),
.B(n_298),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_301),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_362),
.B(n_333),
.Y(n_376)
);

NOR3xp33_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_305),
.C(n_230),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_295),
.B1(n_299),
.B2(n_203),
.Y(n_379)
);

NAND2x1p5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_184),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_280),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g382 ( 
.A1(n_357),
.A2(n_198),
.B1(n_204),
.B2(n_189),
.Y(n_382)
);

CKINVDCx8_ASAP7_75t_R g383 ( 
.A(n_352),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_170),
.B(n_226),
.C(n_225),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

AOI21x1_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_208),
.B(n_205),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_334),
.B(n_231),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_376),
.A2(n_207),
.B(n_206),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_209),
.B1(n_211),
.B2(n_213),
.Y(n_389)
);

O2A1O1Ixp33_ASAP7_75t_SL g390 ( 
.A1(n_372),
.A2(n_244),
.B(n_215),
.C(n_217),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_252),
.B(n_218),
.Y(n_391)
);

AOI221x1_ASAP7_75t_L g392 ( 
.A1(n_368),
.A2(n_347),
.B1(n_344),
.B2(n_247),
.C(n_242),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_364),
.A2(n_250),
.B(n_222),
.C(n_223),
.Y(n_393)
);

AO21x2_ASAP7_75t_L g394 ( 
.A1(n_371),
.A2(n_375),
.B(n_373),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_SL g395 ( 
.A(n_383),
.B(n_270),
.Y(n_395)
);

CKINVDCx9p33_ASAP7_75t_R g396 ( 
.A(n_381),
.Y(n_396)
);

OR2x6_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_354),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_246),
.B(n_236),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_370),
.A2(n_214),
.B(n_238),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_378),
.A2(n_284),
.B1(n_297),
.B2(n_239),
.Y(n_400)
);

NAND2x1p5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_352),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_241),
.B(n_335),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_377),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_379),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_402),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_389),
.A2(n_366),
.B(n_365),
.C(n_384),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_391),
.A2(n_382),
.B1(n_318),
.B2(n_320),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_393),
.A2(n_328),
.B1(n_356),
.B2(n_38),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_29),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_396),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_35),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_40),
.C(n_46),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_418),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_415),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_408),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_414),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_407),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_416),
.A2(n_398),
.B(n_405),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_409),
.A2(n_399),
.B(n_390),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_421),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_428),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_432),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_392),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_430),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_429),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_433),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_425),
.Y(n_441)
);

AND4x1_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_395),
.C(n_410),
.D(n_437),
.Y(n_442)
);

NAND4xp25_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_438),
.C(n_417),
.D(n_426),
.Y(n_443)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_411),
.Y(n_444)
);

AOI221x1_ASAP7_75t_L g445 ( 
.A1(n_442),
.A2(n_431),
.B1(n_50),
.B2(n_52),
.C(n_58),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_445),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_444),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_424),
.B(n_64),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_448),
.Y(n_449)
);

NAND5xp2_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_447),
.C(n_69),
.D(n_78),
.E(n_80),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_48),
.B1(n_81),
.B2(n_82),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.Y(n_452)
);


endmodule