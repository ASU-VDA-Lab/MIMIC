module fake_jpeg_26082_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_21),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_8),
.CI(n_12),
.CON(n_27),
.SN(n_27)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_15),
.B1(n_9),
.B2(n_16),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_25),
.B1(n_17),
.B2(n_18),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.C(n_31),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_16),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR3xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_11),
.C(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_39),
.C(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_13),
.B1(n_16),
.B2(n_10),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_29),
.C(n_25),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR3xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_44),
.C(n_27),
.Y(n_46)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_36),
.A3(n_27),
.B1(n_26),
.B2(n_34),
.C(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_37),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_42),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.A3(n_10),
.B1(n_8),
.B2(n_6),
.C1(n_5),
.C2(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_43),
.B1(n_38),
.B2(n_28),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_50),
.C(n_51),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_8),
.B(n_50),
.Y(n_54)
);


endmodule