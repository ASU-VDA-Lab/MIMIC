module fake_ariane_1280_n_1731 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1731);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1731;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_2),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_15),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_43),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_43),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_23),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_51),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_20),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_48),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_45),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_81),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_108),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_85),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_36),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_48),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_36),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_60),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_39),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_83),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_128),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_59),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_62),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

BUFx8_ASAP7_75t_SL g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_10),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_117),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_35),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_74),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_63),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_69),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_44),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_27),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_101),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_16),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_4),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_70),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_7),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_75),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_114),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_87),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_1),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_40),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_103),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_13),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_29),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_38),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_91),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_96),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_99),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_134),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_50),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_32),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_40),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_38),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_139),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_46),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_97),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_37),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_52),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_122),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_79),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_125),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_89),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_132),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_119),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_16),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_66),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_12),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_80),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_22),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_19),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_126),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_52),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_129),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_73),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_130),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_42),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_37),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_0),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_49),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_19),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_247),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_191),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_230),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_155),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_157),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_170),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_170),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_157),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_153),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_161),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_161),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_186),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_149),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_186),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_150),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_173),
.B(n_2),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_173),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_156),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_174),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_174),
.B(n_3),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_203),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_179),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_187),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_207),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_196),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_187),
.B(n_3),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_188),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_160),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_180),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_190),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_188),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_162),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_196),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_180),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_199),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_190),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_180),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_199),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_202),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_202),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_208),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_190),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_208),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_180),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_213),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_203),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_213),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_167),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_159),
.B(n_5),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_167),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_205),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_167),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_159),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_205),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_217),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_167),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_217),
.B(n_6),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_228),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_169),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_228),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_240),
.B(n_7),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_190),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_240),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_215),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_252),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_171),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_374),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_276),
.Y(n_378)
);

BUFx8_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_252),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_276),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_210),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_336),
.B(n_344),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_260),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

CKINVDCx11_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_336),
.B(n_249),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_249),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_330),
.A2(n_266),
.B1(n_256),
.B2(n_258),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_304),
.A2(n_296),
.B1(n_269),
.B2(n_300),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_306),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_340),
.B(n_249),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_309),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_312),
.B(n_313),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_312),
.B(n_260),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_319),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_321),
.B(n_264),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_340),
.B(n_241),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_195),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_264),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_269),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_342),
.B(n_284),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_305),
.B(n_249),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_346),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_347),
.B(n_284),
.Y(n_434)
);

CKINVDCx11_ASAP7_75t_R g435 ( 
.A(n_332),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_303),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_348),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_317),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_305),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_377),
.B(n_344),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_381),
.B(n_310),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_415),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_314),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_364),
.C(n_318),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_377),
.B(n_310),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_L g467 ( 
.A1(n_399),
.A2(n_328),
.B1(n_356),
.B2(n_333),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_322),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_377),
.B(n_328),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_286),
.Y(n_479)
);

BUFx6f_ASAP7_75t_SL g480 ( 
.A(n_384),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_425),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_322),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_398),
.B(n_311),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g485 ( 
.A1(n_399),
.A2(n_356),
.B1(n_333),
.B2(n_360),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_366),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_427),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_437),
.B(n_320),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_429),
.B(n_326),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_386),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_385),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_427),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_391),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_435),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_436),
.B(n_339),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_431),
.B(n_314),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_426),
.B(n_316),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_426),
.B(n_316),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

BUFx4f_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_411),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_395),
.B(n_405),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_382),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_437),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_406),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_437),
.B(n_354),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_395),
.B(n_286),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_426),
.A2(n_369),
.B1(n_365),
.B2(n_372),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_362),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_385),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_416),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_426),
.B(n_378),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_413),
.B(n_362),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_392),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_392),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_382),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_397),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_397),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_413),
.B(n_418),
.C(n_417),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_378),
.B(n_324),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_384),
.B(n_296),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_397),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_400),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_408),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_400),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_413),
.B(n_375),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_400),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_413),
.B(n_341),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_405),
.B(n_302),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_438),
.B(n_351),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_L g551 ( 
.A(n_387),
.B(n_282),
.C(n_324),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_378),
.A2(n_372),
.B1(n_368),
.B2(n_365),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_420),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_420),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_408),
.B(n_190),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_421),
.B(n_368),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_389),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_378),
.B(n_353),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_419),
.B(n_353),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_390),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_422),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_390),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_430),
.B(n_360),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_393),
.B(n_371),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_432),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_389),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_433),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_379),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_390),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_419),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_390),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_409),
.Y(n_582)
);

AND3x1_ASAP7_75t_L g583 ( 
.A(n_409),
.B(n_256),
.C(n_241),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_390),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_439),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_396),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_441),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_441),
.B(n_288),
.C(n_212),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_479),
.A2(n_515),
.B1(n_523),
.B2(n_454),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_562),
.B(n_443),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_569),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_577),
.B(n_443),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_569),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_444),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_582),
.B(n_444),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_572),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_448),
.B(n_507),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_473),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_572),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_448),
.B(n_303),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_494),
.B(n_414),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_515),
.B(n_422),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_544),
.B(n_414),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_577),
.B(n_424),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_479),
.B(n_424),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_451),
.B(n_428),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_580),
.B(n_355),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_473),
.B(n_434),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_479),
.B(n_428),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_479),
.A2(n_434),
.B1(n_422),
.B2(n_299),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_479),
.B(n_422),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_479),
.B(n_422),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_448),
.A2(n_285),
.B(n_295),
.C(n_272),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_479),
.B(n_422),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_584),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_473),
.B(n_178),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_533),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

BUFx6f_ASAP7_75t_SL g627 ( 
.A(n_564),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_577),
.B(n_299),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_533),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_379),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_577),
.B(n_402),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_484),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_578),
.B(n_379),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_523),
.B(n_460),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_578),
.B(n_541),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_534),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_357),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_512),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_507),
.A2(n_396),
.B1(n_367),
.B2(n_373),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_523),
.B(n_379),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_473),
.B(n_183),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_500),
.B(n_301),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_465),
.B(n_184),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_212),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_477),
.B(n_516),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_534),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_518),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_515),
.B(n_212),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_523),
.B(n_194),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_516),
.B(n_192),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_515),
.A2(n_181),
.B1(n_222),
.B2(n_204),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_484),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_517),
.B(n_402),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_536),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_517),
.B(n_510),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_486),
.B(n_371),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_541),
.B(n_507),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_518),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_536),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_517),
.B(n_402),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_519),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_523),
.B(n_307),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_541),
.B(n_307),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_490),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_523),
.B(n_358),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_502),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_507),
.A2(n_358),
.B1(n_373),
.B2(n_367),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_460),
.B(n_361),
.Y(n_672)
);

AOI22x1_ASAP7_75t_L g673 ( 
.A1(n_445),
.A2(n_258),
.B1(n_285),
.B2(n_272),
.Y(n_673)
);

BUFx5_ASAP7_75t_L g674 ( 
.A(n_446),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_504),
.B(n_361),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_510),
.B(n_402),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_519),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_548),
.B(n_211),
.C(n_193),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_504),
.B(n_359),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_540),
.B(n_363),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_535),
.B(n_221),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_522),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_540),
.B(n_546),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_541),
.A2(n_164),
.B1(n_273),
.B2(n_218),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_540),
.B(n_164),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_540),
.B(n_218),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_L g688 ( 
.A(n_573),
.B(n_402),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_535),
.B(n_223),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_510),
.B(n_529),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_510),
.B(n_224),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_526),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_509),
.B(n_273),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_542),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_528),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_509),
.B(n_279),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_529),
.B(n_226),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_525),
.A2(n_295),
.B(n_294),
.C(n_279),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_509),
.B(n_563),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_515),
.B(n_212),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_564),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_509),
.B(n_280),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_515),
.B(n_212),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_528),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_563),
.B(n_280),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_231),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_564),
.B(n_292),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_564),
.B(n_292),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_521),
.B(n_288),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_542),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_530),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_529),
.B(n_531),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_587),
.A2(n_294),
.B1(n_283),
.B2(n_181),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_531),
.B(n_232),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_531),
.B(n_233),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_549),
.B(n_244),
.C(n_262),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_480),
.A2(n_468),
.B1(n_482),
.B2(n_467),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_531),
.B(n_234),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_456),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_530),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_538),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_543),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_524),
.B(n_237),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_553),
.B(n_238),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_538),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_468),
.A2(n_245),
.B1(n_268),
.B2(n_293),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_554),
.B(n_242),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_554),
.B(n_246),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_555),
.B(n_250),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_513),
.B(n_402),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_480),
.B(n_251),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_493),
.B(n_551),
.C(n_464),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_555),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_456),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_545),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_513),
.B(n_195),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_SL g740 ( 
.A(n_480),
.B(n_253),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_556),
.B(n_254),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_556),
.B(n_259),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_557),
.B(n_277),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_557),
.A2(n_151),
.B(n_291),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_468),
.B(n_281),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_559),
.B(n_290),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_468),
.B(n_283),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_456),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_513),
.B(n_567),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_490),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_485),
.A2(n_283),
.B1(n_288),
.B2(n_219),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_547),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_559),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_464),
.B(n_288),
.C(n_289),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_468),
.A2(n_298),
.B1(n_152),
.B2(n_287),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_567),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_565),
.B(n_154),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_565),
.B(n_163),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_571),
.B(n_165),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_547),
.Y(n_761)
);

BUFx4f_ASAP7_75t_L g762 ( 
.A(n_666),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_683),
.A2(n_539),
.B(n_532),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_603),
.A2(n_482),
.B1(n_541),
.B2(n_550),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_613),
.B(n_482),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_670),
.B(n_570),
.Y(n_767)
);

BUFx4f_ASAP7_75t_L g768 ( 
.A(n_666),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_610),
.A2(n_539),
.B(n_482),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_610),
.A2(n_482),
.B(n_571),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_595),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_606),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_609),
.A2(n_576),
.B(n_574),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_660),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_647),
.A2(n_576),
.B(n_574),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_615),
.A2(n_475),
.B(n_472),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_701),
.B(n_586),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_613),
.B(n_701),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_648),
.B(n_561),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_645),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_634),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_612),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_680),
.B(n_501),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_651),
.A2(n_588),
.B(n_586),
.Y(n_784)
);

CKINVDCx6p67_ASAP7_75t_R g785 ( 
.A(n_627),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_648),
.B(n_588),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_679),
.B(n_461),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_607),
.B(n_590),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_615),
.A2(n_475),
.B(n_472),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_604),
.B(n_590),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_606),
.B(n_583),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_604),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_702),
.A2(n_705),
.B(n_598),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_598),
.A2(n_591),
.B(n_449),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_645),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_628),
.A2(n_591),
.B(n_449),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_703),
.A2(n_660),
.B1(n_594),
.B2(n_646),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_628),
.A2(n_450),
.B(n_446),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_640),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_692),
.A2(n_453),
.B(n_450),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_660),
.A2(n_583),
.B1(n_461),
.B2(n_459),
.Y(n_801)
);

AO21x1_ASAP7_75t_L g802 ( 
.A1(n_739),
.A2(n_481),
.B(n_478),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_646),
.B(n_481),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_611),
.A2(n_616),
.B(n_735),
.C(n_748),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_692),
.A2(n_455),
.B(n_453),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_650),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_658),
.A2(n_462),
.B(n_455),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_665),
.B(n_461),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_659),
.B(n_487),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_614),
.B(n_639),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_666),
.B(n_461),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_693),
.B(n_487),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_630),
.B(n_456),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_637),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_669),
.B(n_567),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_720),
.B(n_458),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_714),
.B(n_459),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_672),
.B(n_469),
.C(n_459),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_693),
.B(n_488),
.C(n_491),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_748),
.A2(n_452),
.B(n_457),
.C(n_447),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_699),
.A2(n_469),
.B1(n_459),
.B2(n_508),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_739),
.A2(n_658),
.B(n_656),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_699),
.B(n_488),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_637),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_636),
.A2(n_447),
.B1(n_452),
.B2(n_457),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_637),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_645),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_755),
.A2(n_491),
.B(n_498),
.Y(n_828)
);

AOI21xp33_ASAP7_75t_L g829 ( 
.A1(n_745),
.A2(n_498),
.B(n_508),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_708),
.B(n_698),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_596),
.A2(n_470),
.B(n_445),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_752),
.A2(n_499),
.B(n_476),
.C(n_492),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_661),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_600),
.A2(n_469),
.B(n_503),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_663),
.A2(n_568),
.B(n_589),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_708),
.B(n_463),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_664),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_698),
.B(n_463),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_752),
.A2(n_499),
.B(n_476),
.C(n_492),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_601),
.A2(n_469),
.B(n_506),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_645),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_677),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_682),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_635),
.B(n_283),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_624),
.B(n_458),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_757),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_671),
.B(n_466),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_633),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_663),
.A2(n_608),
.B(n_690),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_675),
.B(n_466),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_671),
.B(n_471),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_685),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_593),
.A2(n_511),
.B(n_495),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_642),
.B(n_471),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_624),
.B(n_458),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_714),
.B(n_496),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_729),
.A2(n_496),
.B(n_503),
.C(n_505),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_717),
.A2(n_505),
.B(n_511),
.C(n_552),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_641),
.B(n_552),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_643),
.B(n_560),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_694),
.A2(n_474),
.B(n_483),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_697),
.A2(n_474),
.B1(n_483),
.B2(n_585),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_706),
.A2(n_474),
.B(n_483),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_676),
.A2(n_474),
.B(n_483),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_643),
.B(n_560),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_655),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_676),
.A2(n_489),
.B(n_585),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_678),
.B(n_489),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_713),
.A2(n_489),
.B(n_585),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_625),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_625),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_629),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_695),
.B(n_687),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_734),
.B(n_489),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_723),
.A2(n_585),
.B(n_581),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_704),
.B(n_581),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_709),
.B(n_710),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_629),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_707),
.B(n_581),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_632),
.A2(n_589),
.B(n_579),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_653),
.B(n_568),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_745),
.A2(n_558),
.B1(n_579),
.B2(n_566),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_724),
.A2(n_458),
.B(n_566),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_718),
.A2(n_592),
.B(n_10),
.C(n_14),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_654),
.B(n_458),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_728),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_641),
.B(n_288),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_736),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_757),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_652),
.A2(n_458),
.B(n_566),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_644),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_734),
.B(n_490),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_754),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_653),
.A2(n_592),
.B(n_566),
.C(n_527),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_667),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_599),
.A2(n_566),
.B1(n_527),
.B2(n_497),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_681),
.A2(n_527),
.B(n_497),
.C(n_490),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_632),
.A2(n_527),
.B(n_497),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_668),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_597),
.A2(n_527),
.B(n_497),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_668),
.Y(n_903)
);

OAI321xp33_ASAP7_75t_L g904 ( 
.A1(n_684),
.A2(n_219),
.A3(n_497),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_904)
);

BUFx12f_ASAP7_75t_L g905 ( 
.A(n_667),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_623),
.A2(n_278),
.B1(n_275),
.B2(n_274),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_618),
.A2(n_219),
.B(n_270),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_681),
.B(n_166),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_689),
.B(n_168),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_689),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_715),
.B(n_9),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_730),
.B(n_172),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_740),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_620),
.B(n_176),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_731),
.A2(n_17),
.B(n_21),
.C(n_23),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_619),
.A2(n_219),
.B(n_267),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_667),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_617),
.A2(n_271),
.B(n_265),
.C(n_263),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_712),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_602),
.A2(n_261),
.B(n_257),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_626),
.A2(n_255),
.B(n_248),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_756),
.A2(n_243),
.B1(n_239),
.B2(n_236),
.Y(n_922)
);

NOR2x2_ASAP7_75t_L g923 ( 
.A(n_605),
.B(n_26),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_622),
.A2(n_229),
.B(n_227),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_631),
.A2(n_225),
.B1(n_220),
.B2(n_182),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_732),
.B(n_185),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_721),
.B(n_189),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_758),
.A2(n_206),
.B(n_216),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_621),
.A2(n_219),
.B(n_93),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_214),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_759),
.A2(n_209),
.B(n_201),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_722),
.A2(n_200),
.B(n_198),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_712),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_742),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_743),
.B(n_197),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_688),
.A2(n_86),
.B(n_143),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_722),
.A2(n_76),
.B(n_142),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_747),
.A2(n_29),
.B(n_30),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_760),
.A2(n_30),
.B(n_31),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_716),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_715),
.B(n_33),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_726),
.B(n_94),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_744),
.A2(n_727),
.B(n_719),
.Y(n_943)
);

INVx11_ASAP7_75t_L g944 ( 
.A(n_673),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_767),
.B(n_778),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_771),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_772),
.B(n_700),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_910),
.B(n_737),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_783),
.A2(n_750),
.B1(n_749),
.B2(n_737),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_766),
.A2(n_749),
.B1(n_751),
.B2(n_750),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_788),
.A2(n_751),
.B(n_733),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_782),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_848),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_791),
.A2(n_674),
.B1(n_733),
.B2(n_711),
.Y(n_954)
);

OAI22x1_ASAP7_75t_L g955 ( 
.A1(n_764),
.A2(n_761),
.B1(n_753),
.B2(n_746),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_812),
.A2(n_751),
.B(n_753),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_868),
.A2(n_751),
.B1(n_761),
.B2(n_746),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_830),
.B(n_638),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_893),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_781),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_823),
.A2(n_738),
.B(n_716),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_810),
.Y(n_962)
);

CKINVDCx11_ASAP7_75t_R g963 ( 
.A(n_785),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_889),
.A2(n_738),
.B1(n_725),
.B2(n_696),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_804),
.A2(n_686),
.B(n_662),
.C(n_657),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_779),
.B(n_649),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_836),
.A2(n_674),
.B(n_100),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_775),
.A2(n_674),
.B(n_88),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_SL g969 ( 
.A(n_792),
.B(n_674),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_799),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_911),
.A2(n_674),
.B1(n_39),
.B2(n_41),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_775),
.A2(n_674),
.B(n_109),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_784),
.A2(n_867),
.B(n_862),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_770),
.A2(n_34),
.B(n_45),
.C(n_46),
.Y(n_974)
);

INVx8_ASAP7_75t_L g975 ( 
.A(n_905),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_786),
.A2(n_34),
.B1(n_50),
.B2(n_54),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_765),
.B(n_54),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_845),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_777),
.B(n_55),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_827),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_762),
.B(n_57),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_806),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_833),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_908),
.A2(n_58),
.B(n_59),
.C(n_72),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_943),
.B(n_58),
.C(n_104),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_SL g986 ( 
.A1(n_944),
.A2(n_116),
.B(n_118),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_762),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_850),
.B(n_847),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_851),
.B(n_138),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_909),
.A2(n_146),
.B(n_938),
.C(n_803),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_827),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_837),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_939),
.B(n_931),
.C(n_928),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_842),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_773),
.A2(n_793),
.B(n_856),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_768),
.B(n_797),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_838),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_770),
.A2(n_787),
.B(n_793),
.C(n_769),
.Y(n_998)
);

BUFx4f_ASAP7_75t_L g999 ( 
.A(n_913),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_769),
.B(n_876),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_768),
.B(n_811),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_914),
.A2(n_927),
.B1(n_857),
.B2(n_844),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_912),
.A2(n_930),
.B(n_926),
.C(n_935),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_852),
.B(n_809),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_827),
.B(n_857),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_792),
.A2(n_888),
.B1(n_843),
.B2(n_895),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_861),
.B(n_879),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_858),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_890),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_846),
.B(n_774),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_SL g1011 ( 
.A(n_922),
.B(n_941),
.C(n_939),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_819),
.A2(n_776),
.B1(n_789),
.B2(n_817),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_820),
.A2(n_904),
.B(n_818),
.C(n_883),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_800),
.A2(n_805),
.B(n_877),
.Y(n_1014)
);

BUFx4f_ASAP7_75t_L g1015 ( 
.A(n_780),
.Y(n_1015)
);

INVx6_ASAP7_75t_L g1016 ( 
.A(n_774),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_915),
.A2(n_934),
.B(n_860),
.C(n_918),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_903),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_817),
.A2(n_801),
.B1(n_821),
.B2(n_894),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_872),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_849),
.A2(n_763),
.B1(n_774),
.B2(n_827),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_800),
.A2(n_805),
.B(n_877),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_875),
.B(n_774),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_814),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_873),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_863),
.A2(n_865),
.B(n_871),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_919),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_849),
.A2(n_763),
.B1(n_932),
.B2(n_824),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_SL g1029 ( 
.A(n_846),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_824),
.Y(n_1030)
);

INVx3_ASAP7_75t_SL g1031 ( 
.A(n_923),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_829),
.A2(n_870),
.B(n_859),
.C(n_796),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_SL g1033 ( 
.A(n_780),
.B(n_795),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_826),
.B(n_881),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_940),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_863),
.A2(n_871),
.B(n_865),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_874),
.B(n_901),
.Y(n_1037)
);

AND3x1_ASAP7_75t_SL g1038 ( 
.A(n_921),
.B(n_931),
.C(n_928),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_880),
.A2(n_933),
.B1(n_878),
.B2(n_816),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_907),
.A2(n_916),
.B(n_882),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_891),
.B(n_839),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_790),
.A2(n_825),
.B(n_886),
.C(n_906),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_835),
.A2(n_902),
.B(n_900),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_891),
.B(n_780),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_795),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_854),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_900),
.A2(n_834),
.B(n_840),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_832),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_925),
.A2(n_899),
.B(n_864),
.C(n_828),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_815),
.B(n_808),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_902),
.A2(n_822),
.B(n_885),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_917),
.B(n_855),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_795),
.B(n_897),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_917),
.B(n_841),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_841),
.B(n_897),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_855),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_920),
.A2(n_924),
.B(n_796),
.C(n_794),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_884),
.A2(n_887),
.B1(n_813),
.B2(n_936),
.Y(n_1058)
);

INVxp33_ASAP7_75t_SL g1059 ( 
.A(n_920),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_841),
.B(n_853),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_794),
.Y(n_1061)
);

AND2x6_ASAP7_75t_SL g1062 ( 
.A(n_855),
.B(n_924),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_942),
.A2(n_802),
.B1(n_937),
.B2(n_929),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_853),
.B(n_897),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_834),
.A2(n_840),
.B(n_831),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_798),
.A2(n_885),
.B(n_896),
.C(n_831),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_853),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_898),
.B(n_798),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_807),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_866),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_807),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_869),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_892),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_781),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_910),
.A2(n_766),
.B(n_613),
.C(n_454),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_910),
.A2(n_766),
.B(n_613),
.C(n_454),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_781),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_910),
.A2(n_766),
.B(n_613),
.C(n_454),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_810),
.A2(n_454),
.B1(n_485),
.B2(n_671),
.C(n_641),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_782),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_781),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1007),
.B(n_988),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_971),
.A2(n_1075),
.B1(n_1076),
.B2(n_1078),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1000),
.A2(n_969),
.B(n_1003),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1040),
.A2(n_1068),
.B(n_995),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_971),
.A2(n_945),
.B(n_974),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1014),
.A2(n_1022),
.B(n_1065),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_960),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_1012),
.A2(n_1011),
.B(n_1059),
.C(n_1006),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_980),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_946),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_958),
.B(n_966),
.Y(n_1093)
);

AO21x2_ASAP7_75t_L g1094 ( 
.A1(n_1047),
.A2(n_1066),
.B(n_1073),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_976),
.A2(n_1028),
.B(n_981),
.C(n_990),
.Y(n_1095)
);

OAI22x1_ASAP7_75t_L g1096 ( 
.A1(n_1031),
.A2(n_1002),
.B1(n_996),
.B2(n_1001),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1068),
.A2(n_967),
.B(n_968),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_958),
.B(n_1023),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_962),
.B(n_1031),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1023),
.B(n_997),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_972),
.A2(n_1036),
.B(n_1026),
.Y(n_1101)
);

AO32x2_ASAP7_75t_L g1102 ( 
.A1(n_957),
.A2(n_1019),
.A3(n_1021),
.B1(n_950),
.B2(n_985),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1013),
.A2(n_1032),
.B(n_1049),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_951),
.A2(n_956),
.B(n_961),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1079),
.A2(n_979),
.B1(n_977),
.B2(n_947),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1017),
.A2(n_1057),
.B(n_1042),
.Y(n_1107)
);

CKINVDCx11_ASAP7_75t_R g1108 ( 
.A(n_975),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_965),
.A2(n_1061),
.B(n_1069),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_975),
.B(n_1030),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1063),
.A2(n_1041),
.B(n_1070),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1070),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_949),
.A2(n_984),
.B(n_1060),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1048),
.A2(n_1046),
.B(n_1071),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1020),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1058),
.A2(n_955),
.B(n_989),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1039),
.A2(n_1005),
.B(n_1050),
.Y(n_1117)
);

AOI221x1_ASAP7_75t_L g1118 ( 
.A1(n_1050),
.A2(n_979),
.B1(n_977),
.B2(n_948),
.C(n_1004),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_997),
.B(n_1004),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1025),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_985),
.A2(n_993),
.B(n_948),
.C(n_986),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_970),
.Y(n_1122)
);

AO21x1_ASAP7_75t_L g1123 ( 
.A1(n_1034),
.A2(n_1052),
.B(n_1005),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1072),
.A2(n_1053),
.B(n_1044),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_987),
.B(n_959),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1080),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_982),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1039),
.A2(n_1064),
.B(n_1056),
.Y(n_1128)
);

AOI221x1_ASAP7_75t_L g1129 ( 
.A1(n_1052),
.A2(n_1018),
.B1(n_1035),
.B2(n_1027),
.C(n_1081),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_993),
.B(n_978),
.C(n_954),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1037),
.A2(n_964),
.B(n_1010),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_999),
.A2(n_953),
.B1(n_1029),
.B2(n_1024),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_983),
.A2(n_992),
.B(n_1074),
.C(n_1009),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1015),
.A2(n_1054),
.B(n_1077),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_975),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_994),
.Y(n_1136)
);

AND2x2_ASAP7_75t_SL g1137 ( 
.A(n_980),
.B(n_991),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1008),
.B(n_964),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1045),
.A2(n_1067),
.B(n_1038),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1055),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_1038),
.A2(n_1045),
.B(n_1067),
.Y(n_1141)
);

INVx2_ASAP7_75t_R g1142 ( 
.A(n_1062),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1033),
.A2(n_1055),
.B(n_991),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_1016),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_980),
.A2(n_991),
.B(n_1016),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_980),
.A2(n_991),
.B(n_1016),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_963),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_980),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_997),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1007),
.B(n_988),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_946),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1031),
.A2(n_1002),
.B1(n_399),
.B2(n_484),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1030),
.B(n_774),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_960),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_1078),
.C(n_1003),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1157)
);

AO32x2_ASAP7_75t_L g1158 ( 
.A1(n_1028),
.A2(n_957),
.A3(n_1012),
.B1(n_1019),
.B2(n_1021),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_980),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_946),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_1078),
.C(n_766),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1030),
.B(n_774),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_960),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_952),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_946),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1007),
.B(n_988),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1007),
.B(n_988),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_971),
.A2(n_1076),
.B1(n_1078),
.B2(n_1075),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_960),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_980),
.B(n_991),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1007),
.B(n_988),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1066),
.A2(n_998),
.A3(n_1058),
.B(n_955),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_945),
.B(n_670),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_960),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1002),
.B(n_945),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_960),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1079),
.A2(n_454),
.B1(n_485),
.B2(n_381),
.C(n_467),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1190)
);

AOI31xp67_ASAP7_75t_L g1191 ( 
.A1(n_1000),
.A2(n_1068),
.A3(n_1071),
.B(n_1073),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1007),
.B(n_988),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_975),
.B(n_603),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_960),
.Y(n_1194)
);

INVx8_ASAP7_75t_L g1195 ( 
.A(n_975),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1066),
.A2(n_998),
.A3(n_1058),
.B(n_955),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_SL g1198 ( 
.A(n_987),
.B(n_762),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1007),
.B(n_988),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_1078),
.C(n_1003),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_960),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_960),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_1078),
.C(n_1003),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_980),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_973),
.A2(n_1000),
.B(n_998),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_971),
.A2(n_1076),
.B1(n_1078),
.B2(n_1075),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1036),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_1000),
.A2(n_1068),
.B(n_998),
.C(n_995),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1007),
.B(n_988),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1007),
.B(n_988),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_998),
.A3(n_1058),
.B(n_955),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_960),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_971),
.A2(n_1076),
.B1(n_1078),
.B2(n_1075),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1075),
.A2(n_804),
.B(n_1076),
.Y(n_1215)
);

O2A1O1Ixp5_ASAP7_75t_SL g1216 ( 
.A1(n_1070),
.A2(n_1068),
.B(n_1000),
.C(n_1061),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1075),
.A2(n_454),
.B(n_670),
.C(n_1076),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_960),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_997),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_960),
.Y(n_1220)
);

AOI221x1_ASAP7_75t_L g1221 ( 
.A1(n_974),
.A2(n_1028),
.B1(n_1011),
.B2(n_938),
.C(n_976),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1108),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1181),
.B(n_1099),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_1156),
.B2(n_1200),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1195),
.Y(n_1225)
);

INVx8_ASAP7_75t_L g1226 ( 
.A(n_1195),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1084),
.A2(n_1174),
.B1(n_1207),
.B2(n_1214),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1089),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1153),
.A2(n_1087),
.B1(n_1184),
.B2(n_1142),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1096),
.A2(n_1214),
.B1(n_1084),
.B2(n_1174),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1207),
.A2(n_1103),
.B1(n_1215),
.B2(n_1098),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1195),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1122),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1118),
.A2(n_1103),
.B1(n_1221),
.B2(n_1215),
.Y(n_1234)
);

BUFx4f_ASAP7_75t_L g1235 ( 
.A(n_1105),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1119),
.B(n_1083),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1083),
.A2(n_1199),
.B1(n_1177),
.B2(n_1150),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1151),
.Y(n_1238)
);

BUFx8_ASAP7_75t_L g1239 ( 
.A(n_1147),
.Y(n_1239)
);

INVx11_ASAP7_75t_L g1240 ( 
.A(n_1176),
.Y(n_1240)
);

INVx2_ASAP7_75t_R g1241 ( 
.A(n_1216),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1150),
.A2(n_1192),
.B1(n_1172),
.B2(n_1173),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1172),
.A2(n_1211),
.B1(n_1173),
.B2(n_1177),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1135),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1192),
.A2(n_1199),
.B1(n_1210),
.B2(n_1211),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1176),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1217),
.A2(n_1204),
.B(n_1121),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1098),
.A2(n_1119),
.B1(n_1093),
.B2(n_1210),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1127),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1115),
.A2(n_1126),
.B1(n_1120),
.B2(n_1169),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1093),
.A2(n_1138),
.B1(n_1149),
.B2(n_1219),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1130),
.A2(n_1095),
.B1(n_1107),
.B2(n_1092),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1136),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_1125),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1111),
.A2(n_1107),
.B1(n_1130),
.B2(n_1198),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1162),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1155),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1138),
.A2(n_1100),
.B1(n_1123),
.B2(n_1213),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1171),
.A2(n_1193),
.B1(n_1132),
.B2(n_1085),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1193),
.A2(n_1110),
.B1(n_1100),
.B2(n_1140),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1094),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1110),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1140),
.A2(n_1082),
.B1(n_1206),
.B2(n_1197),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1175),
.A2(n_1220),
.B1(n_1218),
.B2(n_1203),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1176),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1152),
.A2(n_1165),
.B1(n_1168),
.B2(n_1183),
.Y(n_1267)
);

BUFx2_ASAP7_75t_SL g1268 ( 
.A(n_1144),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1178),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1182),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1187),
.B(n_1201),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1143),
.B(n_1091),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1148),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_1148),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1194),
.A2(n_1113),
.B1(n_1198),
.B2(n_1154),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1109),
.A2(n_1114),
.B1(n_1164),
.B2(n_1154),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1133),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1134),
.A2(n_1090),
.B1(n_1164),
.B2(n_1163),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1157),
.A2(n_1190),
.B1(n_1186),
.B2(n_1097),
.Y(n_1279)
);

OAI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1088),
.A2(n_1109),
.B(n_1101),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1114),
.A2(n_1117),
.B1(n_1131),
.B2(n_1128),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1129),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1124),
.A2(n_1141),
.B1(n_1091),
.B2(n_1158),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1141),
.A2(n_1159),
.B1(n_1205),
.B2(n_1145),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1191),
.Y(n_1285)
);

CKINVDCx16_ASAP7_75t_R g1286 ( 
.A(n_1159),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1158),
.A2(n_1205),
.B1(n_1159),
.B2(n_1102),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1102),
.A2(n_1158),
.B1(n_1139),
.B2(n_1205),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1146),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1104),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1209),
.Y(n_1291)
);

CKINVDCx6p67_ASAP7_75t_R g1292 ( 
.A(n_1102),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1178),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1196),
.A2(n_1212),
.B1(n_1116),
.B2(n_1112),
.Y(n_1294)
);

CKINVDCx6p67_ASAP7_75t_R g1295 ( 
.A(n_1086),
.Y(n_1295)
);

CKINVDCx14_ASAP7_75t_R g1296 ( 
.A(n_1196),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1160),
.A2(n_1161),
.B1(n_1166),
.B2(n_1170),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1179),
.A2(n_1180),
.B1(n_1185),
.B2(n_1189),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1202),
.A2(n_1188),
.B(n_1106),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1208),
.A2(n_1106),
.B1(n_1188),
.B2(n_454),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1195),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1153),
.A2(n_1188),
.B1(n_1079),
.B2(n_587),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1089),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1105),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1106),
.A2(n_910),
.B1(n_1076),
.B2(n_1075),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1108),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_454),
.B2(n_1079),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1137),
.B(n_774),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_1118),
.B2(n_1174),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1106),
.A2(n_910),
.B1(n_1076),
.B2(n_1075),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1195),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1108),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1110),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_1118),
.B2(n_1174),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1195),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1153),
.A2(n_1188),
.B1(n_1079),
.B2(n_587),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1153),
.A2(n_1188),
.B1(n_1079),
.B2(n_587),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1089),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_1110),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1108),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1188),
.A2(n_1079),
.B1(n_1106),
.B2(n_1087),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1151),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1106),
.A2(n_1184),
.B1(n_844),
.B2(n_587),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_454),
.B2(n_1079),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1089),
.Y(n_1330)
);

BUFx2_ASAP7_75t_SL g1331 ( 
.A(n_1144),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1144),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1176),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1089),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1089),
.Y(n_1335)
);

BUFx10_ASAP7_75t_L g1336 ( 
.A(n_1110),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1188),
.A2(n_1079),
.B1(n_1106),
.B2(n_1087),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1188),
.A2(n_1079),
.B1(n_1106),
.B2(n_1087),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1089),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1084),
.A2(n_396),
.B1(n_311),
.B2(n_587),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1285),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1269),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1292),
.B(n_1296),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1227),
.B(n_1271),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1228),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1303),
.A2(n_1342),
.B1(n_1304),
.B2(n_1324),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1234),
.A2(n_1282),
.B(n_1262),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1246),
.B(n_1293),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1290),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1279),
.A2(n_1267),
.B(n_1297),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1227),
.B(n_1231),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1298),
.A2(n_1264),
.B(n_1281),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1233),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1249),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1253),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1291),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1309),
.A2(n_1329),
.B(n_1224),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1231),
.B(n_1257),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1270),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1295),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1305),
.B(n_1322),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1262),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1330),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1334),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1335),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1326),
.A2(n_1337),
.B(n_1338),
.C(n_1230),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1339),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1261),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1277),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1287),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1294),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1294),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1288),
.A2(n_1272),
.B(n_1258),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1284),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1311),
.A2(n_1317),
.B(n_1300),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1265),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1289),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1316),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1248),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1223),
.B(n_1255),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1289),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1234),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1311),
.A2(n_1312),
.B1(n_1307),
.B2(n_1340),
.C(n_1341),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1266),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1256),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1240),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1252),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1236),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1276),
.A2(n_1299),
.B(n_1247),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1255),
.A2(n_1342),
.B(n_1341),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1251),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1278),
.A2(n_1260),
.B(n_1241),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1313),
.B(n_1243),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1276),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1259),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1333),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1241),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1316),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1275),
.A2(n_1229),
.B(n_1243),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1263),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1303),
.A2(n_1340),
.B1(n_1304),
.B2(n_1324),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1273),
.Y(n_1405)
);

CKINVDCx6p67_ASAP7_75t_R g1406 ( 
.A(n_1222),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1242),
.B(n_1245),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1321),
.A2(n_1302),
.B1(n_1320),
.B2(n_1319),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1323),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1336),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1242),
.A2(n_1245),
.B(n_1310),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1250),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1237),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1238),
.B(n_1327),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1274),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1274),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1286),
.B(n_1268),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1328),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1225),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1331),
.B(n_1332),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1232),
.B(n_1301),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1386),
.A2(n_1321),
.B(n_1235),
.C(n_1226),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1363),
.B(n_1254),
.Y(n_1423)
);

NOR2x1_ASAP7_75t_L g1424 ( 
.A(n_1417),
.B(n_1362),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1386),
.A2(n_1235),
.B1(n_1308),
.B2(n_1325),
.C(n_1315),
.Y(n_1425)
);

AOI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1393),
.A2(n_1226),
.B1(n_1306),
.B2(n_1239),
.C(n_1244),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1388),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1393),
.A2(n_1226),
.B(n_1314),
.C(n_1318),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1347),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1406),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1378),
.A2(n_1239),
.B(n_1359),
.C(n_1369),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1359),
.A2(n_1378),
.B(n_1353),
.C(n_1390),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1396),
.B(n_1391),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1409),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1404),
.A2(n_1348),
.B1(n_1353),
.B2(n_1408),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1383),
.B(n_1346),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1360),
.B(n_1390),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1345),
.B(n_1420),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1358),
.B(n_1373),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1373),
.B(n_1407),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1392),
.A2(n_1385),
.B(n_1382),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1392),
.A2(n_1404),
.B(n_1408),
.C(n_1385),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1350),
.B(n_1364),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1357),
.B(n_1361),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1349),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1398),
.A2(n_1414),
.B1(n_1413),
.B2(n_1389),
.Y(n_1448)
);

AO32x2_ASAP7_75t_L g1449 ( 
.A1(n_1381),
.A2(n_1410),
.A3(n_1401),
.B1(n_1349),
.B2(n_1394),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1413),
.A2(n_1375),
.B1(n_1374),
.B2(n_1394),
.C(n_1418),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1414),
.B(n_1357),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1365),
.A2(n_1352),
.B(n_1354),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1402),
.A2(n_1374),
.B1(n_1375),
.B2(n_1418),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1389),
.A2(n_1387),
.B1(n_1397),
.B2(n_1362),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1361),
.B(n_1366),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1365),
.A2(n_1354),
.B(n_1376),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1402),
.A2(n_1411),
.B(n_1400),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1402),
.A2(n_1411),
.B(n_1400),
.Y(n_1458)
);

AO32x2_ASAP7_75t_L g1459 ( 
.A1(n_1381),
.A2(n_1401),
.A3(n_1410),
.B1(n_1349),
.B2(n_1379),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1379),
.A2(n_1349),
.B1(n_1397),
.B2(n_1372),
.C(n_1367),
.Y(n_1460)
);

INVx5_ASAP7_75t_SL g1461 ( 
.A(n_1406),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1411),
.A2(n_1351),
.B(n_1365),
.Y(n_1462)
);

AO32x2_ASAP7_75t_L g1463 ( 
.A1(n_1371),
.A2(n_1351),
.A3(n_1370),
.B1(n_1368),
.B2(n_1395),
.Y(n_1463)
);

NOR3xp33_ASAP7_75t_SL g1464 ( 
.A(n_1405),
.B(n_1399),
.C(n_1421),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1354),
.A2(n_1376),
.B(n_1377),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1403),
.B(n_1405),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1463),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1395),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1429),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1435),
.A2(n_1395),
.B1(n_1412),
.B2(n_1376),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1463),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1427),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1463),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1446),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1424),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1444),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1452),
.B(n_1343),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1447),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1452),
.B(n_1384),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1344),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1455),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1466),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1440),
.B(n_1436),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1454),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1451),
.Y(n_1487)
);

OAI211xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1422),
.A2(n_1415),
.B(n_1416),
.C(n_1419),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1456),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1439),
.B(n_1380),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1434),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1476),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1485),
.B(n_1438),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1476),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1477),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1468),
.B(n_1442),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1469),
.Y(n_1499)
);

AOI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1488),
.A2(n_1422),
.B(n_1432),
.C(n_1431),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1457),
.Y(n_1501)
);

NAND4xp25_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1425),
.C(n_1435),
.D(n_1431),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1480),
.B(n_1464),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1443),
.C(n_1426),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1476),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1469),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1478),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1472),
.B(n_1449),
.Y(n_1509)
);

BUFx2_ASAP7_75t_SL g1510 ( 
.A(n_1486),
.Y(n_1510)
);

NAND2x1_ASAP7_75t_L g1511 ( 
.A(n_1491),
.B(n_1464),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1469),
.Y(n_1512)
);

OAI31xp33_ASAP7_75t_L g1513 ( 
.A1(n_1488),
.A2(n_1443),
.A3(n_1428),
.B(n_1448),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1486),
.B(n_1434),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1488),
.A2(n_1450),
.B1(n_1428),
.B2(n_1453),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1445),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1467),
.A2(n_1447),
.B(n_1462),
.Y(n_1517)
);

INVxp67_ASAP7_75t_SL g1518 ( 
.A(n_1479),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1470),
.A2(n_1460),
.B1(n_1471),
.B2(n_1467),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.B(n_1458),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1490),
.B(n_1459),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1459),
.Y(n_1522)
);

INVxp67_ASAP7_75t_SL g1523 ( 
.A(n_1479),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1495),
.B(n_1498),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1495),
.B(n_1484),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1496),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1495),
.B(n_1484),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.B(n_1484),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1506),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1520),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1506),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1498),
.B(n_1487),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1520),
.B(n_1475),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1520),
.B(n_1475),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1499),
.Y(n_1536)
);

AND2x2_ASAP7_75t_SL g1537 ( 
.A(n_1503),
.B(n_1465),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1487),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1430),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1486),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1497),
.B(n_1482),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1499),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1481),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1506),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1482),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1497),
.B(n_1482),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1507),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1507),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1477),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1504),
.A2(n_1473),
.B1(n_1423),
.B2(n_1481),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1503),
.B(n_1489),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1512),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1481),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1552),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1552),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1536),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1551),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1554),
.B(n_1504),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1554),
.A2(n_1500),
.B1(n_1515),
.B2(n_1502),
.Y(n_1565)
);

NAND2x1_ASAP7_75t_SL g1566 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1551),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1430),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1545),
.B(n_1510),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1510),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1556),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1556),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1544),
.Y(n_1574)
);

NAND2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1493),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1544),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1529),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1543),
.B(n_1494),
.Y(n_1582)
);

CKINVDCx16_ASAP7_75t_R g1583 ( 
.A(n_1541),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1545),
.B(n_1501),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1545),
.A2(n_1505),
.B(n_1514),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1526),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1526),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1549),
.B(n_1494),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1529),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1553),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1539),
.B(n_1516),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1550),
.B(n_1505),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1509),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1539),
.B(n_1516),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1541),
.Y(n_1598)
);

OR2x6_ASAP7_75t_L g1599 ( 
.A(n_1555),
.B(n_1514),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1570),
.B(n_1541),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1583),
.B(n_1539),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1602)
);

INVxp33_ASAP7_75t_L g1603 ( 
.A(n_1568),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1574),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1581),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1564),
.B(n_1557),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1577),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1578),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

NAND4xp25_ASAP7_75t_L g1611 ( 
.A(n_1564),
.B(n_1500),
.C(n_1542),
.D(n_1513),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1534),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1575),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1560),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1578),
.B(n_1533),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1598),
.B(n_1533),
.Y(n_1618)
);

AO21x1_ASAP7_75t_L g1619 ( 
.A1(n_1598),
.A2(n_1555),
.B(n_1523),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1561),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1562),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1542),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1567),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1571),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1570),
.A2(n_1513),
.B(n_1537),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1572),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1534),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1558),
.Y(n_1631)
);

NAND2x1_ASAP7_75t_L g1632 ( 
.A(n_1570),
.B(n_1525),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1559),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1584),
.B(n_1535),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1611),
.A2(n_1515),
.B1(n_1599),
.B2(n_1575),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1593),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1626),
.A2(n_1585),
.B(n_1595),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.B(n_1606),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1603),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1612),
.B(n_1586),
.Y(n_1642)
);

OAI332xp33_ASAP7_75t_L g1643 ( 
.A1(n_1631),
.A2(n_1569),
.A3(n_1594),
.B1(n_1596),
.B2(n_1590),
.B3(n_1582),
.C1(n_1588),
.C2(n_1518),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1631),
.Y(n_1644)
);

AOI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1519),
.B1(n_1537),
.B2(n_1467),
.C1(n_1483),
.C2(n_1471),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1604),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1619),
.A2(n_1595),
.B(n_1599),
.C(n_1523),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1608),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1609),
.B(n_1597),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1619),
.A2(n_1519),
.B1(n_1474),
.B2(n_1471),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1618),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1461),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1615),
.A2(n_1563),
.B(n_1597),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1608),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1614),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1630),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1615),
.A2(n_1563),
.B(n_1502),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1641),
.B(n_1634),
.Y(n_1660)
);

AOI321xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1643),
.A2(n_1632),
.A3(n_1600),
.B1(n_1617),
.B2(n_1613),
.C(n_1634),
.Y(n_1661)
);

AOI22x1_ASAP7_75t_SL g1662 ( 
.A1(n_1635),
.A2(n_1615),
.B1(n_1633),
.B2(n_1461),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1651),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1651),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1639),
.B(n_1623),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1652),
.A2(n_1632),
.B1(n_1600),
.B2(n_1566),
.C(n_1599),
.Y(n_1666)
);

INVxp33_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1653),
.B(n_1613),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1653),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1654),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

AOI31xp33_ASAP7_75t_L g1672 ( 
.A1(n_1639),
.A2(n_1563),
.A3(n_1624),
.B(n_1627),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1637),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1637),
.B(n_1600),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1659),
.A2(n_1600),
.B1(n_1628),
.B2(n_1492),
.Y(n_1675)
);

NAND2x1_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1622),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1642),
.B(n_1576),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1645),
.A2(n_1607),
.B1(n_1605),
.B2(n_1503),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1659),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1672),
.A2(n_1636),
.B1(n_1655),
.B2(n_1648),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1660),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1674),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1672),
.B(n_1658),
.Y(n_1684)
);

XOR2x2_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1642),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1662),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1675),
.A2(n_1644),
.B(n_1656),
.C(n_1657),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1668),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1678),
.A2(n_1607),
.B1(n_1605),
.B2(n_1517),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1683),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1688),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1680),
.B(n_1675),
.C(n_1666),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1663),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1679),
.A2(n_1661),
.B(n_1670),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1682),
.B(n_1664),
.Y(n_1696)
);

NOR3x1_ASAP7_75t_L g1697 ( 
.A(n_1685),
.B(n_1669),
.C(n_1671),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1686),
.B(n_1640),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1687),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1689),
.B(n_1686),
.C(n_1646),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1694),
.A2(n_1649),
.B1(n_1657),
.B2(n_1656),
.C(n_1647),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1694),
.A2(n_1649),
.B1(n_1647),
.B2(n_1627),
.C(n_1624),
.Y(n_1702)
);

AOI221x1_ASAP7_75t_L g1703 ( 
.A1(n_1695),
.A2(n_1616),
.B1(n_1621),
.B2(n_1620),
.C(n_1625),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1693),
.A2(n_1616),
.B1(n_1677),
.B2(n_1614),
.C(n_1591),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1703),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1692),
.C(n_1690),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1704),
.A2(n_1698),
.B1(n_1691),
.B2(n_1697),
.C(n_1696),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1701),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1702),
.A2(n_1650),
.B(n_1617),
.C(n_1622),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1703),
.Y(n_1710)
);

INVxp33_ASAP7_75t_L g1711 ( 
.A(n_1706),
.Y(n_1711)
);

XOR2xp5_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_1461),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1710),
.B(n_1650),
.Y(n_1713)
);

NAND4xp75_ASAP7_75t_L g1714 ( 
.A(n_1707),
.B(n_1629),
.C(n_1591),
.D(n_1525),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1629),
.Y(n_1715)
);

OAI211xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1713),
.A2(n_1709),
.B(n_1518),
.C(n_1530),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1711),
.B(n_1492),
.C(n_1555),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1715),
.B(n_1492),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1718),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1719),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1720),
.B(n_1714),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1712),
.B1(n_1717),
.B2(n_1716),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1721),
.A2(n_1722),
.B1(n_1389),
.B2(n_1492),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1721),
.A2(n_1530),
.B1(n_1548),
.B2(n_1547),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1723),
.A2(n_1555),
.B1(n_1517),
.B2(n_1547),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1538),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1532),
.B(n_1548),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1726),
.B(n_1525),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1728),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_R g1730 ( 
.A1(n_1729),
.A2(n_1527),
.B1(n_1528),
.B2(n_1555),
.C(n_1546),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1423),
.B(n_1555),
.C(n_1535),
.Y(n_1731)
);


endmodule