module fake_ariane_1975_n_1705 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1705);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1705;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_46),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_57),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_50),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_35),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_26),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_95),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_10),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_134),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_45),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

BUFx8_ASAP7_75t_SL g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_35),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_12),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_52),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_29),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_14),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_90),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_29),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_100),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_64),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_4),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_113),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_59),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_55),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_38),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_16),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_14),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_69),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_153),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_48),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_118),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_102),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_97),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_20),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_18),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_34),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_144),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_65),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_78),
.Y(n_239)
);

INVxp33_ASAP7_75t_R g240 ( 
.A(n_48),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_16),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_117),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_141),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_89),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_54),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_23),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_80),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_88),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_32),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_60),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_66),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_42),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_4),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_3),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_33),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_96),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_15),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_140),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_59),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_128),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_19),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_73),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_47),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_103),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_31),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_83),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_98),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_81),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_21),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_9),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_39),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_130),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_27),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_61),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_104),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_137),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_23),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_5),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_31),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_18),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_79),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_156),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_93),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_8),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_63),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_91),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_149),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_24),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_146),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_37),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_87),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_116),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_20),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_49),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_24),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_21),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_216),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_171),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_185),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_175),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_182),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_278),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_216),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_186),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_220),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_250),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_216),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_216),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_216),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_261),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_269),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_216),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_194),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_216),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_276),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_175),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_162),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_231),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_275),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_197),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_275),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_275),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_263),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_224),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_224),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_224),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_281),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_321),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_224),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_224),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_246),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_246),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_246),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_204),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_221),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_208),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_246),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_246),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_249),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_211),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_265),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_265),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_160),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_249),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_265),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_265),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_265),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_193),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_195),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_193),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_168),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_217),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_212),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_256),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_256),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_260),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_260),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_295),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_215),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_196),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_177),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_353),
.A2(n_240),
.B1(n_160),
.B2(n_187),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_380),
.B(n_196),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_164),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_295),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_334),
.A2(n_210),
.B1(n_242),
.B2(n_191),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_369),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_325),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_332),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_343),
.A2(n_187),
.B1(n_184),
.B2(n_180),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_356),
.B(n_190),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_163),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_218),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_333),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_342),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_385),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_200),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_335),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_337),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_372),
.B(n_379),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_337),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_338),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_213),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_328),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_339),
.Y(n_451)
);

CKINVDCx8_ASAP7_75t_R g452 ( 
.A(n_327),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_344),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_327),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_344),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_346),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_345),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_348),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_388),
.B(n_200),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_389),
.B(n_227),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_350),
.B(n_167),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_350),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_354),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_389),
.B(n_258),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_355),
.B(n_181),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_301),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_340),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_371),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_411),
.B(n_349),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_460),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_347),
.B1(n_352),
.B2(n_376),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_455),
.B(n_363),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

NOR2x1p5_ASAP7_75t_L g496 ( 
.A(n_450),
.B(n_375),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_351),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_423),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_467),
.B(n_377),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_455),
.B(n_381),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_395),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_425),
.A2(n_403),
.B1(n_285),
.B2(n_316),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_427),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_432),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_408),
.B(n_402),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_453),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_371),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_411),
.B(n_391),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_202),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_444),
.B(n_373),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_391),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_475),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_477),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

BUFx6f_ASAP7_75t_SL g536 ( 
.A(n_432),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_444),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_441),
.B(n_373),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_432),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_421),
.B(n_364),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_440),
.B(n_393),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_440),
.B(n_393),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_473),
.A2(n_294),
.B1(n_322),
.B2(n_270),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_429),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_436),
.B(n_394),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_408),
.B(n_341),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_473),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_394),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_165),
.C(n_164),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_434),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_473),
.A2(n_293),
.B1(n_262),
.B2(n_268),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_471),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_452),
.B(n_161),
.Y(n_562)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_471),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_452),
.B(n_161),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g570 ( 
.A(n_467),
.B(n_165),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_441),
.A2(n_299),
.B1(n_305),
.B2(n_280),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_433),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_459),
.B(n_170),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_418),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_170),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_435),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_441),
.B(n_374),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_446),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_435),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_198),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_434),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_451),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_451),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_425),
.B(n_173),
.C(n_169),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_457),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_426),
.B(n_172),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_461),
.B(n_374),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_433),
.Y(n_594)
);

AND3x2_ASAP7_75t_L g595 ( 
.A(n_426),
.B(n_317),
.C(n_287),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_433),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_463),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_436),
.B(n_396),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_436),
.B(n_396),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_172),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_461),
.A2(n_282),
.B1(n_302),
.B2(n_309),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_461),
.B(n_378),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_466),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_437),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_416),
.A2(n_184),
.B1(n_180),
.B2(n_174),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_434),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_461),
.B(n_214),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_461),
.B(n_219),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_416),
.B(n_173),
.C(n_169),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_464),
.B(n_285),
.C(n_174),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_462),
.B(n_397),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_420),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_434),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_462),
.A2(n_314),
.B1(n_226),
.B2(n_166),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_439),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_462),
.A2(n_289),
.B1(n_297),
.B2(n_303),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_439),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_439),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_406),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_469),
.B(n_397),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_480),
.B(n_421),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_579),
.B(n_464),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_480),
.B(n_454),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_583),
.B(n_470),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_538),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_556),
.B(n_470),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_538),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_538),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_480),
.B(n_454),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_623),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_556),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_563),
.B(n_439),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_623),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_526),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_304),
.C(n_289),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_616),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_519),
.B(n_368),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_480),
.B(n_439),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_563),
.B(n_469),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_482),
.B(n_476),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_525),
.B(n_469),
.Y(n_650)
);

AO221x1_ASAP7_75t_L g651 ( 
.A1(n_608),
.A2(n_407),
.B1(n_308),
.B2(n_206),
.C(n_319),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_499),
.B(n_176),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_526),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_525),
.B(n_406),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_499),
.B(n_222),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_581),
.B(n_176),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_545),
.B(n_424),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_525),
.B(n_415),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_581),
.B(n_178),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_581),
.B(n_178),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_544),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_415),
.Y(n_664)
);

NAND2x1p5_ASAP7_75t_L g665 ( 
.A(n_567),
.B(n_244),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_398),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_534),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_499),
.B(n_223),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_499),
.B(n_230),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_500),
.B(n_232),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_179),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_512),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_545),
.A2(n_316),
.B1(n_313),
.B2(n_235),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_512),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_512),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_537),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_179),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_581),
.B(n_183),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_537),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_612),
.B(n_183),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_542),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_479),
.Y(n_683)
);

INVxp33_ASAP7_75t_L g684 ( 
.A(n_543),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_518),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_523),
.B(n_188),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_543),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_558),
.B(n_189),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_523),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_531),
.B(n_189),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_548),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_509),
.B(n_233),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_479),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_531),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_544),
.B(n_296),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_481),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_573),
.B(n_298),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_545),
.B(n_494),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_481),
.Y(n_700)
);

BUFx12f_ASAP7_75t_SL g701 ( 
.A(n_545),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_573),
.B(n_298),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_483),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_544),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_544),
.B(n_306),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_551),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_594),
.B(n_306),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_496),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_508),
.B(n_237),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_576),
.A2(n_301),
.B1(n_311),
.B2(n_315),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_507),
.B(n_307),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_596),
.B(n_311),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_551),
.A2(n_387),
.B(n_382),
.C(n_383),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_620),
.B(n_410),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_533),
.B(n_315),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_533),
.B(n_252),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_483),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_562),
.B(n_241),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_536),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_568),
.B(n_248),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_620),
.B(n_553),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_533),
.B(n_253),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_481),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_489),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_552),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_557),
.B(n_599),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_SL g727 ( 
.A1(n_521),
.A2(n_407),
.B1(n_410),
.B2(n_313),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_491),
.B(n_399),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_557),
.B(n_257),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_554),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_489),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_552),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_577),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_510),
.B(n_323),
.C(n_259),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_489),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_490),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_490),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_557),
.B(n_266),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_530),
.B(n_272),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_577),
.A2(n_387),
.B(n_383),
.C(n_382),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_599),
.B(n_274),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_496),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_599),
.B(n_283),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_601),
.A2(n_312),
.B1(n_267),
.B2(n_288),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_574),
.B(n_501),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_570),
.B(n_284),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_615),
.B(n_192),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_490),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_615),
.B(n_600),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_589),
.B(n_201),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_530),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_615),
.B(n_203),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_613),
.A2(n_401),
.B1(n_400),
.B2(n_399),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_571),
.A2(n_400),
.B1(n_401),
.B2(n_318),
.C(n_310),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_516),
.A2(n_300),
.B(n_290),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_578),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_492),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_600),
.B(n_205),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_624),
.B(n_592),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_492),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_567),
.A2(n_243),
.B1(n_202),
.B2(n_251),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_614),
.B(n_472),
.C(n_474),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_604),
.B(n_472),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_624),
.B(n_243),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_501),
.B(n_207),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_501),
.B(n_209),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_SL g767 ( 
.A(n_483),
.B(n_225),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_578),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_501),
.B(n_228),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_582),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_582),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_513),
.B(n_251),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_492),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_513),
.B(n_524),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_513),
.B(n_254),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_536),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_641),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_703),
.B(n_516),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_645),
.B(n_517),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_626),
.B(n_602),
.Y(n_780)
);

AOI21x1_ASAP7_75t_L g781 ( 
.A1(n_772),
.A2(n_588),
.B(n_587),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_643),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_703),
.B(n_516),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_648),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_R g785 ( 
.A(n_701),
.B(n_536),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_630),
.B(n_618),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_714),
.A2(n_560),
.B1(n_547),
.B2(n_605),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_658),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_749),
.B(n_604),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_645),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_742),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_653),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_719),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_686),
.B(n_604),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_SL g796 ( 
.A(n_629),
.B(n_588),
.C(n_587),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_629),
.B(n_524),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_663),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_667),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_688),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_656),
.B(n_541),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_656),
.B(n_524),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_649),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_704),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_R g805 ( 
.A(n_776),
.B(n_536),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_719),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_627),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_668),
.B(n_524),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_636),
.B(n_699),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_635),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_636),
.B(n_487),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_666),
.B(n_487),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_668),
.B(n_528),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_669),
.B(n_528),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_727),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_654),
.B(n_528),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_699),
.B(n_487),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_676),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_669),
.B(n_528),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_726),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_693),
.B(n_590),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_666),
.B(n_522),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_625),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_690),
.A2(n_527),
.B1(n_580),
.B2(n_593),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_682),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_625),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_717),
.B(n_631),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_644),
.B(n_595),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_683),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_715),
.A2(n_772),
.B(n_775),
.C(n_716),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_685),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_670),
.B(n_764),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_717),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_692),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_650),
.B(n_520),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_632),
.A2(n_569),
.B1(n_605),
.B2(n_546),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_670),
.B(n_569),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_L g841 ( 
.A1(n_715),
.A2(n_591),
.B(n_550),
.C(n_549),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_695),
.B(n_520),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_683),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_651),
.A2(n_535),
.B1(n_546),
.B2(n_549),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_694),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_662),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_706),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_759),
.B(n_529),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_730),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_725),
.B(n_540),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_764),
.B(n_535),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_733),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_734),
.A2(n_603),
.B1(n_535),
.B2(n_546),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_759),
.B(n_549),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_662),
.A2(n_555),
.B1(n_550),
.B2(n_572),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_732),
.B(n_550),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_673),
.B(n_564),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_687),
.B(n_555),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_691),
.B(n_572),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_759),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_751),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_694),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_756),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_633),
.B(n_529),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_722),
.B(n_572),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_768),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_634),
.B(n_586),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_751),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_728),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_722),
.B(n_586),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_718),
.A2(n_598),
.B1(n_586),
.B2(n_591),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_665),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_703),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_703),
.Y(n_876)
);

AO22x1_ASAP7_75t_L g877 ( 
.A1(n_684),
.A2(n_254),
.B1(n_264),
.B2(n_598),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_771),
.A2(n_597),
.B1(n_598),
.B2(n_511),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_597),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_637),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_640),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_741),
.B(n_478),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_652),
.B(n_539),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_697),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_697),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_R g886 ( 
.A(n_703),
.B(n_539),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_700),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_754),
.A2(n_511),
.B1(n_505),
.B2(n_484),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_758),
.B(n_478),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_700),
.Y(n_890)
);

AND3x2_ASAP7_75t_SL g891 ( 
.A(n_628),
.B(n_264),
.C(n_514),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_678),
.B(n_484),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_745),
.Y(n_893)
);

AND2x2_ASAP7_75t_SL g894 ( 
.A(n_646),
.B(n_505),
.Y(n_894)
);

AND3x1_ASAP7_75t_L g895 ( 
.A(n_709),
.B(n_488),
.C(n_503),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_723),
.Y(n_896)
);

NOR2x1p5_ASAP7_75t_L g897 ( 
.A(n_743),
.B(n_486),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_723),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_SL g899 ( 
.A1(n_709),
.A2(n_277),
.B1(n_229),
.B2(n_234),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_681),
.B(n_488),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_705),
.B(n_539),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_724),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_724),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_774),
.B(n_495),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_755),
.A2(n_720),
.B1(n_773),
.B2(n_736),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_763),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_763),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_731),
.Y(n_909)
);

NOR2x2_ASAP7_75t_L g910 ( 
.A(n_638),
.B(n_493),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_774),
.A2(n_504),
.B(n_495),
.C(n_497),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_729),
.B(n_497),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_720),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_913)
);

AND3x1_ASAP7_75t_L g914 ( 
.A(n_710),
.B(n_502),
.C(n_559),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_731),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_735),
.A2(n_514),
.B1(n_515),
.B2(n_565),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_642),
.B(n_236),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_735),
.A2(n_515),
.B1(n_566),
.B2(n_561),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_746),
.B(n_539),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_744),
.B(n_619),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_738),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_753),
.B(n_561),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_711),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_639),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_657),
.A2(n_559),
.B1(n_585),
.B2(n_621),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_736),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_737),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_689),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_698),
.B(n_565),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_702),
.B(n_566),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_748),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_707),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_748),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_657),
.A2(n_585),
.B1(n_621),
.B2(n_617),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_712),
.B(n_585),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_753),
.B(n_585),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_660),
.B(n_619),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_716),
.B(n_765),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_752),
.B(n_622),
.Y(n_939)
);

BUFx4f_ASAP7_75t_SL g940 ( 
.A(n_750),
.Y(n_940)
);

OAI22xp33_ASAP7_75t_L g941 ( 
.A1(n_786),
.A2(n_661),
.B1(n_671),
.B2(n_761),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_866),
.A2(n_661),
.B(n_679),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_823),
.A2(n_775),
.B(n_769),
.C(n_766),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_807),
.B(n_810),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_871),
.A2(n_659),
.B(n_664),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_800),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_782),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_822),
.A2(n_797),
.B1(n_894),
.B2(n_784),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_834),
.B(n_757),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_804),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_809),
.B(n_762),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_840),
.A2(n_713),
.B(n_740),
.C(n_739),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_787),
.B(n_760),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_812),
.B(n_655),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_893),
.A2(n_773),
.B(n_628),
.C(n_675),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_787),
.B(n_647),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_825),
.B(n_647),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_777),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_937),
.A2(n_674),
.B(n_672),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_893),
.A2(n_796),
.B(n_860),
.C(n_859),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_931),
.Y(n_961)
);

NOR2x1_ASAP7_75t_R g962 ( 
.A(n_791),
.B(n_238),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_778),
.A2(n_674),
.B(n_672),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_803),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_824),
.B(n_767),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_828),
.B(n_619),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_894),
.A2(n_622),
.B1(n_621),
.B2(n_617),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_841),
.A2(n_617),
.B(n_610),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_793),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_783),
.A2(n_610),
.B(n_619),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_801),
.A2(n_610),
.B(n_619),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_784),
.A2(n_609),
.B1(n_607),
.B2(n_247),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_782),
.B(n_607),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_812),
.B(n_609),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_824),
.B(n_0),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_889),
.A2(n_892),
.B(n_900),
.C(n_789),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_899),
.A2(n_245),
.B1(n_239),
.B2(n_271),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_804),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_780),
.B(n_2),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_905),
.A2(n_474),
.B(n_378),
.C(n_417),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_793),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_848),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_905),
.B(n_6),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_938),
.A2(n_498),
.B(n_412),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_792),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_858),
.A2(n_417),
.B(n_414),
.C(n_412),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_795),
.A2(n_414),
.B(n_417),
.C(n_10),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_851),
.B(n_7),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_911),
.A2(n_414),
.B(n_11),
.C(n_17),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_895),
.A2(n_474),
.B1(n_498),
.B2(n_319),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_931),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_781),
.A2(n_474),
.B(n_308),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_SL g993 ( 
.A1(n_802),
.A2(n_9),
.B(n_11),
.C(n_17),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_855),
.A2(n_474),
.B1(n_308),
.B2(n_319),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_846),
.B(n_793),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_L g996 ( 
.A(n_917),
.B(n_255),
.C(n_206),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_826),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_790),
.B(n_413),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_855),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_830),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_793),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_816),
.B(n_25),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_932),
.B(n_921),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_831),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_879),
.A2(n_255),
.B(n_206),
.C(n_195),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_826),
.A2(n_33),
.B(n_37),
.C(n_39),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_835),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_855),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_843),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_816),
.B(n_41),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_788),
.B(n_41),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_806),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_873),
.B(n_798),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_SL g1014 ( 
.A(n_870),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_808),
.B(n_44),
.C(n_46),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_815),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_845),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_794),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_806),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_873),
.B(n_44),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_861),
.B(n_47),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_904),
.A2(n_195),
.B(n_413),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_813),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_841),
.A2(n_53),
.B(n_56),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_814),
.A2(n_413),
.B(n_409),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_790),
.B(n_413),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_799),
.A2(n_58),
.B1(n_413),
.B2(n_409),
.C(n_77),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_819),
.A2(n_413),
.B(n_409),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_940),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_897),
.A2(n_409),
.B1(n_58),
.B2(n_74),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_L g1032 ( 
.A(n_811),
.B(n_409),
.C(n_84),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_928),
.B(n_72),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_839),
.A2(n_94),
.B(n_99),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_818),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_835),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_820),
.B(n_101),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_879),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_821),
.A2(n_106),
.B1(n_111),
.B2(n_120),
.C(n_121),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_940),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_827),
.B(n_122),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_833),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_123),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_857),
.A2(n_126),
.B(n_129),
.C(n_131),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_837),
.B(n_133),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_852),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_847),
.B(n_158),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_856),
.A2(n_138),
.B1(n_139),
.B2(n_147),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_922),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_832),
.A2(n_854),
.B(n_872),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_863),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_790),
.B(n_785),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_907),
.B(n_850),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_853),
.A2(n_880),
.B1(n_867),
.B2(n_864),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_874),
.B(n_881),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_849),
.B(n_862),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_882),
.B(n_842),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_785),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_878),
.A2(n_842),
.B1(n_913),
.B2(n_912),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_884),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_875),
.A2(n_876),
.B(n_930),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_886),
.B(n_805),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_817),
.A2(n_929),
.B(n_901),
.C(n_865),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_887),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_862),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_805),
.B(n_914),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_924),
.B(n_877),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_906),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_878),
.A2(n_913),
.B1(n_906),
.B2(n_865),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_885),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_919),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_936),
.B(n_868),
.Y(n_1072)
);

AOI221x1_ASAP7_75t_L g1073 ( 
.A1(n_1015),
.A2(n_901),
.B1(n_939),
.B2(n_927),
.C(n_896),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1038),
.B(n_1057),
.Y(n_1074)
);

AO22x2_ASAP7_75t_L g1075 ( 
.A1(n_948),
.A2(n_891),
.B1(n_939),
.B2(n_910),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_946),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1050),
.A2(n_934),
.B(n_925),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_957),
.B(n_836),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_944),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1038),
.B(n_898),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_947),
.B(n_919),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1003),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_868),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_945),
.A2(n_903),
.A3(n_890),
.B(n_926),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_960),
.A2(n_935),
.B(n_844),
.C(n_883),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_982),
.B(n_1072),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_941),
.A2(n_844),
.B(n_920),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1055),
.Y(n_1088)
);

INVx3_ASAP7_75t_SL g1089 ( 
.A(n_1014),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_958),
.Y(n_1090)
);

NAND3x1_ASAP7_75t_L g1091 ( 
.A(n_1022),
.B(n_908),
.C(n_891),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_950),
.B(n_836),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_951),
.A2(n_888),
.B(n_838),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_1062),
.B(n_829),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_982),
.B(n_915),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_978),
.B(n_1013),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_985),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_964),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1061),
.A2(n_779),
.B(n_869),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1069),
.A2(n_888),
.B(n_838),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_968),
.A2(n_916),
.B(n_918),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_SL g1102 ( 
.A1(n_1030),
.A2(n_829),
.B1(n_869),
.B2(n_908),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1035),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_978),
.B(n_909),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1046),
.B(n_902),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1040),
.B(n_933),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1059),
.B(n_933),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_966),
.B(n_933),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_973),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_941),
.A2(n_838),
.B(n_1025),
.C(n_1034),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_960),
.A2(n_838),
.B(n_942),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1042),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_943),
.A2(n_970),
.B(n_963),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1005),
.A2(n_955),
.A3(n_956),
.B(n_953),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_986),
.A2(n_971),
.B(n_984),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1002),
.A2(n_1010),
.B1(n_983),
.B2(n_979),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_974),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1008),
.B(n_974),
.Y(n_1118)
);

BUFx10_ASAP7_75t_L g1119 ( 
.A(n_991),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1053),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_1056),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1016),
.B(n_1021),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1054),
.B(n_988),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_1071),
.A2(n_1066),
.B1(n_1048),
.B2(n_977),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_997),
.A2(n_1006),
.B(n_989),
.Y(n_1125)
);

CKINVDCx11_ASAP7_75t_R g1126 ( 
.A(n_961),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1011),
.B(n_975),
.Y(n_1127)
);

OR2x6_ASAP7_75t_L g1128 ( 
.A(n_1058),
.B(n_1052),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_962),
.B(n_1000),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1019),
.B(n_999),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_999),
.B(n_949),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1004),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_995),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1018),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_954),
.B(n_1068),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_954),
.B(n_1064),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_967),
.A2(n_1063),
.B(n_1041),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_997),
.A2(n_1006),
.B(n_989),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1018),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1033),
.A2(n_1043),
.B1(n_1015),
.B2(n_1047),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_990),
.A2(n_952),
.B(n_980),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_952),
.A2(n_1032),
.B(n_1045),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1009),
.B(n_1060),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_987),
.A2(n_1028),
.B(n_1031),
.C(n_1037),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_1018),
.B(n_1036),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1067),
.A2(n_1070),
.A3(n_1017),
.B(n_1051),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1020),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1024),
.A2(n_965),
.B1(n_993),
.B2(n_1032),
.C(n_1049),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1039),
.B(n_1044),
.C(n_972),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_959),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1065),
.B(n_981),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_998),
.A2(n_1027),
.B(n_994),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1018),
.B(n_1036),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_959),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1012),
.B(n_981),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1012),
.B(n_969),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1014),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_996),
.A2(n_969),
.B1(n_1001),
.B2(n_1007),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_976),
.A2(n_871),
.B(n_866),
.Y(n_1159)
);

NAND2x1_ASAP7_75t_L g1160 ( 
.A(n_1065),
.B(n_1007),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_946),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_976),
.A2(n_871),
.B(n_866),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_976),
.A2(n_948),
.B(n_1059),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1055),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1055),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_948),
.A2(n_1069),
.B1(n_1059),
.B2(n_823),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1055),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_812),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1018),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_957),
.B(n_606),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1050),
.A2(n_832),
.B(n_893),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1008),
.B(n_812),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_997),
.B(n_1006),
.C(n_668),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_945),
.A2(n_1005),
.A3(n_1069),
.B(n_1023),
.Y(n_1179)
);

AOI221x1_ASAP7_75t_L g1180 ( 
.A1(n_1015),
.A2(n_1025),
.B1(n_1024),
.B2(n_1048),
.C(n_942),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1015),
.B(n_606),
.C(n_708),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_945),
.A2(n_1005),
.A3(n_1069),
.B(n_1023),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_944),
.B(n_721),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1055),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1015),
.A2(n_449),
.B(n_656),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_992),
.A2(n_1029),
.B(n_1026),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_957),
.B(n_721),
.Y(n_1189)
);

NAND2x1_ASAP7_75t_L g1190 ( 
.A(n_1065),
.B(n_1007),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_957),
.A2(n_721),
.B1(n_714),
.B2(n_438),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1008),
.B(n_812),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_948),
.B(n_825),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_945),
.A2(n_1005),
.A3(n_1069),
.B(n_1023),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1055),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_946),
.Y(n_1196)
);

NOR2x1_ASAP7_75t_R g1197 ( 
.A(n_1040),
.B(n_606),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_950),
.B(n_947),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_946),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1062),
.B(n_835),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_957),
.B(n_721),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_944),
.B(n_721),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_948),
.B(n_825),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_957),
.B(n_606),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1139),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1140),
.B(n_1168),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1169),
.A2(n_1172),
.B(n_1171),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1187),
.A2(n_1116),
.B(n_1168),
.C(n_1144),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1074),
.B(n_1189),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1116),
.A2(n_1138),
.B(n_1142),
.C(n_1178),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1142),
.A2(n_1165),
.B(n_1110),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1184),
.A2(n_1188),
.B(n_1186),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1100),
.A2(n_1093),
.B(n_1178),
.C(n_1138),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1090),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1193),
.A2(n_1203),
.B(n_1123),
.C(n_1148),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1125),
.A2(n_1201),
.B1(n_1087),
.B2(n_1100),
.C(n_1191),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1157),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1139),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1124),
.A2(n_1075),
.B1(n_1087),
.B2(n_1093),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1175),
.A2(n_1204),
.B1(n_1124),
.B2(n_1075),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1118),
.B(n_1094),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1183),
.A2(n_1202),
.B1(n_1149),
.B2(n_1086),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1161),
.Y(n_1224)
);

CKINVDCx6p67_ASAP7_75t_R g1225 ( 
.A(n_1089),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1074),
.B(n_1109),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1079),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1149),
.A2(n_1181),
.B1(n_1198),
.B2(n_1141),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1137),
.A2(n_1141),
.B(n_1180),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1150),
.A2(n_1154),
.A3(n_1073),
.B(n_1085),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1076),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1196),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1122),
.B(n_1088),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1097),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1176),
.A2(n_1077),
.B(n_1111),
.C(n_1107),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1082),
.A2(n_1081),
.B1(n_1176),
.B2(n_1078),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_1147),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1107),
.A2(n_1135),
.A3(n_1158),
.B(n_1131),
.Y(n_1238)
);

BUFx8_ASAP7_75t_L g1239 ( 
.A(n_1199),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1135),
.A2(n_1158),
.A3(n_1080),
.B(n_1143),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1133),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_SL g1242 ( 
.A1(n_1151),
.A2(n_1099),
.B(n_1155),
.Y(n_1242)
);

AO32x2_ASAP7_75t_L g1243 ( 
.A1(n_1102),
.A2(n_1084),
.A3(n_1146),
.B1(n_1114),
.B2(n_1194),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1077),
.A2(n_1152),
.B(n_1101),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1094),
.B(n_1128),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1086),
.A2(n_1096),
.B1(n_1195),
.B2(n_1185),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1092),
.A2(n_1106),
.B(n_1174),
.C(n_1134),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_SL g1248 ( 
.A1(n_1160),
.A2(n_1190),
.B(n_1108),
.C(n_1156),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1117),
.B(n_1173),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1083),
.B(n_1098),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1095),
.A2(n_1136),
.B(n_1143),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1166),
.A2(n_1167),
.B1(n_1170),
.B2(n_1127),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1095),
.A2(n_1136),
.B(n_1112),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1120),
.B(n_1173),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1103),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_1128),
.B1(n_1091),
.B2(n_1104),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1126),
.Y(n_1257)
);

AOI222xp33_ASAP7_75t_L g1258 ( 
.A1(n_1105),
.A2(n_1197),
.B1(n_1177),
.B2(n_1192),
.C1(n_1130),
.C2(n_1117),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1145),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1132),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1177),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1179),
.A2(n_1194),
.B(n_1182),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1153),
.A2(n_1179),
.B(n_1182),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1200),
.A2(n_1179),
.B(n_1182),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1194),
.A2(n_1114),
.B(n_1129),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1119),
.B(n_1114),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1119),
.A2(n_721),
.B1(n_1191),
.B2(n_714),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1090),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1142),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1113),
.A2(n_1164),
.B(n_1162),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1165),
.B(n_1100),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1187),
.A2(n_1116),
.B(n_1168),
.C(n_1144),
.Y(n_1273)
);

AOI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1116),
.A2(n_1140),
.B(n_1178),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1079),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1087),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1090),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_1164),
.B(n_1162),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1140),
.A2(n_1178),
.B1(n_1187),
.B2(n_825),
.Y(n_1280)
);

BUFx8_ASAP7_75t_L g1281 ( 
.A(n_1161),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1168),
.A2(n_1189),
.B1(n_1201),
.B2(n_1100),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1197),
.B(n_575),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1187),
.B(n_1116),
.C(n_1140),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1140),
.A2(n_1178),
.B1(n_1187),
.B2(n_825),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1090),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1076),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1124),
.A2(n_714),
.B1(n_721),
.B2(n_1168),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1140),
.A2(n_1178),
.B1(n_1187),
.B2(n_825),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1116),
.A2(n_1163),
.B(n_1159),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1157),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1189),
.B(n_1201),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1189),
.B(n_1201),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1191),
.A2(n_721),
.B1(n_714),
.B2(n_1175),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1118),
.B(n_1094),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1113),
.A2(n_1164),
.B(n_1162),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1118),
.B(n_1094),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1146),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1124),
.A2(n_714),
.B1(n_721),
.B2(n_1075),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1142),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1124),
.A2(n_714),
.B1(n_721),
.B2(n_1168),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1183),
.B(n_1202),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1079),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1074),
.B(n_1189),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1115),
.A2(n_1164),
.B(n_1162),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1124),
.A2(n_714),
.B1(n_721),
.B2(n_1168),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1128),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1146),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1142),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1121),
.B(n_835),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1087),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1142),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1272),
.B(n_1276),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1226),
.B(n_1227),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1215),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1207),
.A2(n_1274),
.B(n_1273),
.C(n_1209),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1233),
.B(n_1290),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1294),
.B(n_1297),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1221),
.B(n_1288),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1275),
.B(n_1310),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1306),
.A2(n_1289),
.B1(n_1308),
.B2(n_1313),
.Y(n_1329)
);

O2A1O1Ixp5_ASAP7_75t_L g1330 ( 
.A1(n_1207),
.A2(n_1229),
.B(n_1214),
.C(n_1291),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1280),
.A2(n_1286),
.B(n_1211),
.C(n_1284),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1272),
.B(n_1314),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1276),
.B(n_1318),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1311),
.B(n_1295),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1289),
.A2(n_1313),
.B(n_1308),
.C(n_1217),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1234),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1318),
.B(n_1255),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1263),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1295),
.B(n_1299),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1319),
.A2(n_1212),
.B(n_1213),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1300),
.A2(n_1214),
.B1(n_1306),
.B2(n_1267),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1220),
.A2(n_1282),
.B1(n_1228),
.B2(n_1216),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1268),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1277),
.B(n_1287),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1282),
.A2(n_1235),
.B(n_1245),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1254),
.B(n_1232),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1250),
.B(n_1223),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1220),
.A2(n_1223),
.B1(n_1235),
.B2(n_1236),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1299),
.B(n_1246),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1250),
.B(n_1224),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1253),
.B(n_1251),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1246),
.B(n_1252),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1241),
.A2(n_1292),
.B1(n_1256),
.B2(n_1237),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1231),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1252),
.B(n_1253),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1218),
.A2(n_1293),
.B(n_1225),
.Y(n_1356)
);

INVx3_ASAP7_75t_SL g1357 ( 
.A(n_1218),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1249),
.B(n_1301),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1251),
.B(n_1258),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1222),
.B(n_1303),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1241),
.A2(n_1293),
.B1(n_1303),
.B2(n_1301),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1238),
.B(n_1240),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1247),
.A2(n_1283),
.B(n_1242),
.C(n_1248),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1265),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1222),
.A2(n_1303),
.B1(n_1301),
.B2(n_1257),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1281),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1257),
.A2(n_1317),
.B1(n_1261),
.B2(n_1206),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1238),
.B(n_1240),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1262),
.B(n_1238),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1208),
.A2(n_1205),
.B(n_1279),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1271),
.A2(n_1285),
.B(n_1296),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1239),
.A2(n_1281),
.B1(n_1317),
.B2(n_1262),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_1219),
.A2(n_1315),
.B(n_1304),
.C(n_1298),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1239),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1281),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1259),
.A2(n_1244),
.B1(n_1260),
.B2(n_1278),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1259),
.A2(n_1244),
.B1(n_1270),
.B2(n_1278),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1243),
.B(n_1264),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1243),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1230),
.B(n_1302),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1312),
.B(n_1230),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1230),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1269),
.A2(n_1316),
.B(n_1307),
.Y(n_1385)
);

OAI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1289),
.A2(n_1308),
.B1(n_1313),
.B2(n_1300),
.C(n_1221),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1284),
.A2(n_1308),
.B1(n_1313),
.B2(n_1289),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1250),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1266),
.B(n_1272),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1209),
.A2(n_1273),
.B(n_1187),
.C(n_1289),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1225),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1226),
.B(n_1210),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1226),
.B(n_1210),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1233),
.B(n_1290),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1215),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1226),
.B(n_1210),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1209),
.A2(n_1168),
.B(n_1273),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1233),
.B(n_1290),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1269),
.A2(n_1316),
.B(n_1307),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1225),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1226),
.B(n_1210),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1330),
.A2(n_1397),
.B(n_1323),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1329),
.A2(n_1341),
.B1(n_1386),
.B2(n_1387),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1351),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1392),
.B(n_1393),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1369),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1369),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1385),
.B(n_1399),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1364),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1385),
.B(n_1399),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1399),
.B(n_1376),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1337),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1391),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1396),
.B(n_1401),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1376),
.B(n_1380),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1380),
.B(n_1382),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1322),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1383),
.B(n_1340),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1383),
.B(n_1340),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1336),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1343),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1364),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1362),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1377),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1338),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1349),
.B(n_1355),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1364),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1395),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1333),
.A2(n_1384),
.B(n_1378),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1348),
.A2(n_1342),
.B1(n_1347),
.B2(n_1352),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1344),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1381),
.B(n_1368),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1379),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1320),
.B(n_1333),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1370),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1373),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1321),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1370),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1345),
.B(n_1332),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1359),
.A2(n_1335),
.B(n_1390),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1328),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1389),
.B(n_1324),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.B(n_1345),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1370),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1426),
.B(n_1339),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1426),
.B(n_1346),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1325),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1425),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1445),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_L g1453 ( 
.A(n_1427),
.B(n_1353),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1403),
.A2(n_1441),
.B1(n_1431),
.B2(n_1402),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1411),
.B(n_1326),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1411),
.B(n_1350),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1434),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1436),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1434),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1436),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1403),
.A2(n_1327),
.B1(n_1334),
.B2(n_1335),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1441),
.A2(n_1397),
.B1(n_1390),
.B2(n_1365),
.Y(n_1463)
);

AND2x2_ASAP7_75t_SL g1464 ( 
.A(n_1445),
.B(n_1360),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1440),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1413),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1404),
.B(n_1331),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1439),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1446),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1412),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1415),
.B(n_1416),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1441),
.A2(n_1372),
.B1(n_1367),
.B2(n_1358),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1413),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1445),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1454),
.A2(n_1441),
.B1(n_1402),
.B2(n_1431),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1454),
.B(n_1424),
.C(n_1418),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1463),
.A2(n_1418),
.B1(n_1419),
.B2(n_1424),
.C(n_1410),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1463),
.A2(n_1441),
.B1(n_1435),
.B2(n_1416),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1462),
.A2(n_1424),
.B1(n_1437),
.B2(n_1433),
.C(n_1405),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1467),
.B(n_1363),
.C(n_1354),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1462),
.A2(n_1414),
.B1(n_1405),
.B2(n_1440),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1457),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1466),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1448),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1472),
.A2(n_1440),
.B1(n_1438),
.B2(n_1361),
.Y(n_1485)
);

AOI222xp33_ASAP7_75t_L g1486 ( 
.A1(n_1467),
.A2(n_1416),
.B1(n_1415),
.B2(n_1406),
.C1(n_1407),
.C2(n_1423),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1487)
);

AND4x1_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1418),
.C(n_1419),
.D(n_1375),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1457),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1460),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1438),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1458),
.A2(n_1446),
.B(n_1430),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1448),
.B(n_1430),
.C(n_1410),
.D(n_1408),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1440),
.Y(n_1495)
);

NOR4xp25_ASAP7_75t_SL g1496 ( 
.A(n_1473),
.B(n_1375),
.C(n_1374),
.D(n_1422),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1460),
.Y(n_1497)
);

NAND2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1466),
.B(n_1357),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1473),
.B(n_1374),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1450),
.B(n_1443),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1450),
.B(n_1443),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

AOI31xp33_ASAP7_75t_L g1503 ( 
.A1(n_1452),
.A2(n_1366),
.A3(n_1443),
.B(n_1444),
.Y(n_1503)
);

OAI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1474),
.A2(n_1419),
.B(n_1408),
.C(n_1410),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_SL g1505 ( 
.A(n_1450),
.B(n_1357),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1464),
.A2(n_1449),
.B1(n_1453),
.B2(n_1447),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1507)
);

AOI33xp33_ASAP7_75t_L g1508 ( 
.A1(n_1456),
.A2(n_1444),
.A3(n_1417),
.B1(n_1428),
.B2(n_1420),
.B3(n_1421),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_R g1509 ( 
.A(n_1448),
.B(n_1391),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1505),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1482),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1492),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1482),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1476),
.A2(n_1461),
.B(n_1468),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1500),
.B(n_1455),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1509),
.B(n_1400),
.C(n_1451),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1502),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1508),
.B(n_1456),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1491),
.B(n_1449),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1476),
.A2(n_1459),
.B(n_1469),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1480),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1499),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1484),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1494),
.A2(n_1459),
.B(n_1469),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1497),
.B(n_1456),
.Y(n_1528)
);

INVx3_ASAP7_75t_SL g1529 ( 
.A(n_1483),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1484),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1488),
.B(n_1464),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1507),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1492),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1455),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1514),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1514),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1523),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1527),
.B(n_1500),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1518),
.B(n_1477),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1527),
.B(n_1501),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1527),
.B(n_1515),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1529),
.B(n_1488),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1531),
.A2(n_1475),
.B1(n_1481),
.B2(n_1478),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1527),
.B(n_1487),
.Y(n_1546)
);

NAND2x1_ASAP7_75t_SL g1547 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1514),
.B(n_1504),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1493),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1510),
.B(n_1493),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1455),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1506),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1525),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1479),
.C(n_1486),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

AND2x4_ASAP7_75t_SL g1561 ( 
.A(n_1516),
.B(n_1495),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1513),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1517),
.Y(n_1563)
);

CKINVDCx16_ASAP7_75t_R g1564 ( 
.A(n_1524),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1522),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1522),
.A2(n_1485),
.B1(n_1429),
.B2(n_1437),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1530),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1513),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1538),
.B(n_1532),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1532),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1565),
.B(n_1529),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1569),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1569),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1554),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1556),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1554),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1554),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1558),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1526),
.C(n_1498),
.D(n_1528),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1534),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1554),
.B(n_1464),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1465),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1561),
.B(n_1512),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1550),
.B(n_1496),
.Y(n_1589)
);

OAI322xp33_ASAP7_75t_L g1590 ( 
.A1(n_1540),
.A2(n_1536),
.A3(n_1548),
.B1(n_1545),
.B2(n_1563),
.C1(n_1566),
.C2(n_1559),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1540),
.B(n_1528),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1568),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1568),
.Y(n_1596)
);

OAI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1540),
.A2(n_1533),
.B(n_1519),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1549),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1556),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1560),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1561),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1583),
.A2(n_1547),
.B1(n_1567),
.B2(n_1548),
.C(n_1536),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1598),
.B(n_1536),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1595),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1604),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1580),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1580),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1577),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1599),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1590),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1597),
.B(n_1550),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1574),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1574),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1599),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1593),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1589),
.B(n_1551),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1400),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1600),
.Y(n_1621)
);

AO21x2_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1559),
.B(n_1535),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1596),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1579),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1601),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1593),
.A2(n_1545),
.B1(n_1567),
.B2(n_1548),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1586),
.A2(n_1553),
.B1(n_1561),
.B2(n_1551),
.Y(n_1630)
);

OAI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1613),
.A2(n_1592),
.B(n_1553),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1612),
.Y(n_1632)
);

OAI32xp33_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1586),
.A3(n_1592),
.B1(n_1587),
.B2(n_1553),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1629),
.A2(n_1547),
.B(n_1571),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1616),
.B(n_1625),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1614),
.A2(n_1589),
.B(n_1586),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1611),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1575),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1573),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1622),
.A2(n_1533),
.B1(n_1559),
.B2(n_1566),
.C(n_1535),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1622),
.A2(n_1559),
.B1(n_1566),
.B2(n_1535),
.C(n_1537),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1611),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1606),
.A2(n_1566),
.B1(n_1587),
.B2(n_1537),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1626),
.A2(n_1573),
.B(n_1537),
.C(n_1581),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1625),
.B(n_1551),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1549),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1628),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1651),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1631),
.A2(n_1630),
.B1(n_1606),
.B2(n_1561),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1651),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1636),
.B(n_1608),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1647),
.B(n_1607),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1648),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1641),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1644),
.B(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1632),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1656),
.B(n_1644),
.C(n_1635),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1659),
.A2(n_1633),
.B(n_1646),
.Y(n_1664)
);

NOR4xp25_ASAP7_75t_L g1665 ( 
.A(n_1660),
.B(n_1640),
.C(n_1639),
.D(n_1634),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1654),
.A2(n_1645),
.B1(n_1642),
.B2(n_1643),
.C(n_1637),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1655),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1654),
.A2(n_1645),
.B1(n_1618),
.B2(n_1649),
.C(n_1628),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1661),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1658),
.A2(n_1623),
.B(n_1650),
.C(n_1617),
.Y(n_1670)
);

O2A1O1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1653),
.A2(n_1618),
.B(n_1621),
.C(n_1609),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1620),
.Y(n_1672)
);

XNOR2xp5_ASAP7_75t_L g1673 ( 
.A(n_1667),
.B(n_1657),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1664),
.A2(n_1652),
.B(n_1662),
.C(n_1610),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1666),
.A2(n_1619),
.B1(n_1588),
.B2(n_1587),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1676)
);

AOI32xp33_ASAP7_75t_L g1677 ( 
.A1(n_1663),
.A2(n_1542),
.A3(n_1546),
.B1(n_1539),
.B2(n_1541),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1673),
.B(n_1672),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1675),
.B(n_1665),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1674),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1676),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1677),
.B(n_1668),
.Y(n_1682)
);

XNOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1552),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1678),
.B(n_1670),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1683),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1681),
.Y(n_1686)
);

XOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1680),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_SL g1689 ( 
.A(n_1686),
.B(n_1682),
.C(n_1680),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1686),
.B(n_1578),
.C(n_1576),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1688),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1685),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1692),
.B(n_1689),
.C(n_1690),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1693),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1693),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1694),
.B(n_1684),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1687),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1697),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1696),
.A2(n_1578),
.B(n_1576),
.C(n_1581),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1698),
.Y(n_1700)
);

XNOR2xp5_ASAP7_75t_L g1701 ( 
.A(n_1700),
.B(n_1699),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1701),
.A2(n_1582),
.B1(n_1601),
.B2(n_1603),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1582),
.B(n_1602),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1542),
.B1(n_1552),
.B2(n_1546),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1555),
.B(n_1544),
.C(n_1356),
.Y(n_1705)
);


endmodule