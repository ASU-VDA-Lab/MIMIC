module real_jpeg_32050_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_0),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_1),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_1),
.A2(n_175),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_1),
.A2(n_175),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_1),
.A2(n_175),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_100),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_2),
.A2(n_100),
.B1(n_319),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_2),
.A2(n_47),
.B1(n_100),
.B2(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_33),
.B1(n_64),
.B2(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_4),
.A2(n_199),
.B(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_4),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g381 ( 
.A1(n_4),
.A2(n_165),
.A3(n_382),
.B1(n_386),
.B2(n_389),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_4),
.A2(n_347),
.B1(n_423),
.B2(n_428),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_4),
.B(n_138),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_4),
.A2(n_26),
.B1(n_506),
.B2(n_520),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_6),
.A2(n_86),
.B1(n_89),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_6),
.A2(n_93),
.B1(n_150),
.B2(n_154),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_6),
.A2(n_93),
.B1(n_336),
.B2(n_340),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_7),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_117),
.B1(n_120),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_9),
.A2(n_124),
.B1(n_301),
.B2(n_305),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_9),
.A2(n_67),
.B1(n_124),
.B2(n_433),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_9),
.A2(n_124),
.B1(n_494),
.B2(n_497),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_12),
.A2(n_117),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_12),
.A2(n_217),
.B1(n_326),
.B2(n_329),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_12),
.A2(n_217),
.B1(n_460),
.B2(n_465),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_12),
.A2(n_217),
.B1(n_507),
.B2(n_509),
.Y(n_506)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_14),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_14),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_14),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_15),
.A2(n_64),
.B1(n_67),
.B2(n_71),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_48),
.B1(n_71),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_15),
.A2(n_71),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_16),
.A2(n_34),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_16),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_17),
.A2(n_46),
.B1(n_67),
.B2(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_292),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_R g19 ( 
.A(n_20),
.B(n_288),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_246),
.Y(n_20)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_21),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_179),
.C(n_234),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_22),
.B(n_235),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_94),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_24),
.B(n_249),
.C(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_25),
.B(n_53),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_41),
.B2(n_45),
.Y(n_25)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_26),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_26),
.A2(n_45),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_26),
.A2(n_474),
.B1(n_480),
.B2(n_483),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_26),
.A2(n_493),
.B1(n_506),
.B2(n_513),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_29),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_31),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_31),
.Y(n_339)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_32),
.Y(n_210)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_37),
.Y(n_400)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_37),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_37),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_38),
.Y(n_497)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_39),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_40),
.Y(n_449)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_40),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_204),
.B1(n_205),
.B2(n_210),
.Y(n_203)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_44),
.Y(n_242)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_49),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_50),
.Y(n_508)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_63),
.B1(n_72),
.B2(n_85),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_54),
.A2(n_63),
.B1(n_72),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_54),
.A2(n_72),
.B1(n_237),
.B2(n_255),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_54),
.A2(n_72),
.B1(n_85),
.B2(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_54),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_54),
.A2(n_72),
.B1(n_432),
.B2(n_458),
.Y(n_486)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AO21x2_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_73),
.B(n_79),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_58),
.Y(n_451)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_66),
.Y(n_464)
);

BUFx6f_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_69),
.Y(n_257)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_72),
.A2(n_315),
.B1(n_375),
.B2(n_377),
.Y(n_374)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_72),
.Y(n_437)
);

NAND2xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_78),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_79),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_88),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_92),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_137),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_95),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_105),
.B1(n_116),
.B2(n_125),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_96),
.A2(n_105),
.B1(n_125),
.B2(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_98),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_105),
.A2(n_125),
.B1(n_216),
.B2(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_105),
.B(n_347),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_108),
.Y(n_427)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_126),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_135),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_133),
.Y(n_313)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_149),
.B1(n_157),
.B2(n_172),
.Y(n_137)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_138),
.A2(n_149),
.B1(n_157),
.B2(n_172),
.Y(n_250)
);

AOI22x1_ASAP7_75t_L g268 ( 
.A1(n_138),
.A2(n_149),
.B1(n_157),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_138),
.A2(n_157),
.B1(n_299),
.B2(n_307),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_159),
.B(n_165),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_139)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_145),
.Y(n_388)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_173),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g324 ( 
.A1(n_158),
.A2(n_224),
.B1(n_300),
.B2(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_158),
.A2(n_224),
.B1(n_325),
.B2(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_178),
.Y(n_274)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_179),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_211),
.C(n_222),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_202),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_181),
.B(n_202),
.Y(n_358)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.A3(n_187),
.B1(n_192),
.B2(n_198),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g349 ( 
.A1(n_182),
.A2(n_184),
.A3(n_187),
.B1(n_192),
.B2(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_202),
.A2(n_203),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_204),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_204),
.A2(n_205),
.B1(n_335),
.B2(n_342),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_204),
.A2(n_335),
.B1(n_397),
.B2(n_405),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_204),
.A2(n_492),
.B1(n_498),
.B2(n_499),
.Y(n_491)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_212),
.A2(n_222),
.B1(n_223),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_229),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_230),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_241),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_263),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_258),
.B(n_262),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_259),
.Y(n_262)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_286),
.B2(n_287),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_275),
.B2(n_276),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_368),
.B(n_541),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_359),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_351),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_296),
.B(n_351),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_322),
.C(n_348),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_297),
.B(n_538),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_308),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_320),
.C(n_321),
.Y(n_354)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_320),
.B2(n_321),
.Y(n_308)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_323),
.B(n_348),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_333),
.C(n_346),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_333),
.A2(n_334),
.B1(n_346),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_344),
.Y(n_524)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_345),
.Y(n_516)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_347),
.B(n_453),
.Y(n_452)
);

OA21x2_ASAP7_75t_SL g467 ( 
.A1(n_347),
.A2(n_452),
.B(n_468),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_347),
.B(n_375),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_347),
.B(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_353),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_361),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.C(n_364),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_365),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AOI21x1_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_536),
.B(n_540),
.Y(n_369)
);

OAI21x1_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_438),
.B(n_535),
.Y(n_370)
);

AOI211xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_411),
.B(n_416),
.C(n_417),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_372),
.A2(n_411),
.B(n_416),
.C(n_417),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_413),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_380),
.B1(n_409),
.B2(n_410),
.Y(n_373)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_374),
.B(n_409),
.C(n_412),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_375),
.A2(n_458),
.B1(n_466),
.B2(n_467),
.Y(n_457)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_378),
.B1(n_431),
.B2(n_437),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_395),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_381),
.A2(n_395),
.B1(n_396),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_403),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.C(n_430),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_418),
.B(n_532),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_420),
.A2(n_421),
.B1(n_430),
.B2(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_437),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_529),
.B(n_534),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_489),
.B(n_528),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_472),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_441),
.B(n_472),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_457),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_442),
.B(n_457),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_445),
.B(n_446),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_450),
.B(n_452),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx4f_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_464),
.Y(n_471)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_484),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_473),
.B(n_486),
.C(n_487),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_485),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_486),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_503),
.B(n_527),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_502),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_491),
.B(n_502),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_SL g499 ( 
.A(n_500),
.Y(n_499)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_504),
.A2(n_518),
.B(n_526),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_517),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_505),
.B(n_517),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_530),
.B(n_531),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_537),
.B(n_539),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_537),
.B(n_539),
.Y(n_540)
);

OAI21xp33_ASAP7_75t_L g541 ( 
.A1(n_542),
.A2(n_543),
.B(n_548),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_544),
.B(n_546),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_544),
.B(n_546),
.Y(n_548)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);


endmodule