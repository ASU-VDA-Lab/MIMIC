module fake_jpeg_13710_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_44),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_6),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_11),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_30),
.B1(n_45),
.B2(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_50),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_60),
.B1(n_53),
.B2(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_22),
.B1(n_35),
.B2(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_59),
.B1(n_64),
.B2(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.C(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_51),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_83),
.C(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_75),
.B1(n_79),
.B2(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_59),
.B1(n_64),
.B2(n_57),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_74),
.B1(n_81),
.B2(n_57),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_96),
.B1(n_87),
.B2(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_98),
.C(n_86),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_102),
.B(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_108),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_91),
.Y(n_111)
);


endmodule