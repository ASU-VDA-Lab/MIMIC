module fake_jpeg_24446_n_323 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_0),
.Y(n_71)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_70),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_10),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_59),
.B(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_30),
.B1(n_37),
.B2(n_22),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_69),
.B1(n_73),
.B2(n_40),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_27),
.B1(n_36),
.B2(n_24),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_27),
.B1(n_36),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_27),
.B1(n_24),
.B2(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_19),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_32),
.B1(n_37),
.B2(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_38),
.B1(n_28),
.B2(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_81),
.Y(n_102)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_21),
.B1(n_34),
.B2(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_0),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_40),
.B1(n_26),
.B2(n_35),
.Y(n_86)
);

CKINVDCx9p33_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_12),
.C(n_17),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_100),
.C(n_12),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_47),
.B1(n_40),
.B2(n_35),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_49),
.B1(n_62),
.B2(n_52),
.Y(n_155)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_11),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_43),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_43),
.A3(n_48),
.B1(n_49),
.B2(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_116),
.Y(n_136)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_122),
.B(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_31),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_119),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_10),
.B1(n_12),
.B2(n_17),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_63),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_83),
.C(n_43),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_48),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_55),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_143),
.B1(n_123),
.B2(n_144),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_79),
.B1(n_51),
.B2(n_74),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_129),
.B1(n_141),
.B2(n_155),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_137),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_128),
.B(n_110),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_66),
.B1(n_51),
.B2(n_61),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_48),
.B1(n_49),
.B2(n_61),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_52),
.B(n_62),
.C(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_43),
.Y(n_180)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_153),
.B1(n_117),
.B2(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_92),
.B1(n_104),
.B2(n_113),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_121),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_118),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_87),
.Y(n_166)
);

CKINVDCx12_ASAP7_75t_R g151 ( 
.A(n_88),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_0),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_116),
.C(n_102),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_93),
.A2(n_53),
.B1(n_13),
.B2(n_16),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_93),
.B1(n_120),
.B2(n_95),
.Y(n_178)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_162),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_159),
.B(n_8),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_8),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_102),
.CI(n_101),
.CON(n_163),
.SN(n_163)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_173),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_168),
.B(n_175),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_172),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_107),
.B(n_87),
.C(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_179),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_182),
.B1(n_186),
.B2(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_142),
.C(n_134),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_141),
.A2(n_132),
.B1(n_123),
.B2(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_144),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_188),
.B1(n_179),
.B2(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_96),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_125),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_218),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_133),
.B1(n_132),
.B2(n_139),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_196),
.B1(n_187),
.B2(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_143),
.B1(n_129),
.B2(n_124),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_212),
.B1(n_215),
.B2(n_173),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_144),
.B(n_110),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_219),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_152),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_152),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_146),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_140),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_62),
.B1(n_135),
.B2(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_171),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_231),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_186),
.B(n_160),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_163),
.C(n_175),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_241),
.C(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_163),
.B1(n_174),
.B2(n_166),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_174),
.B1(n_187),
.B2(n_176),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_235),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_176),
.A3(n_4),
.B1(n_5),
.B2(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_9),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_209),
.B(n_11),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_157),
.B1(n_5),
.B2(n_4),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_238)
);

NAND2x1p5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_6),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_193),
.Y(n_240)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_15),
.C(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_201),
.C(n_207),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_200),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_254),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_205),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_204),
.B1(n_212),
.B2(n_208),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_253),
.B1(n_258),
.B2(n_232),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_237),
.B(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_192),
.C(n_206),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_256),
.C(n_241),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_215),
.B1(n_195),
.B2(n_217),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_219),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_209),
.C(n_210),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_195),
.B1(n_203),
.B2(n_213),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_200),
.Y(n_261)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_268),
.C(n_273),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_276),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_257),
.B1(n_262),
.B2(n_231),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_275),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_236),
.C(n_230),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_224),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_274),
.B(n_252),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_224),
.C(n_221),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_235),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_239),
.A3(n_231),
.B1(n_225),
.B2(n_221),
.C1(n_190),
.C2(n_234),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_190),
.C(n_231),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_240),
.B1(n_191),
.B2(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_249),
.B1(n_253),
.B2(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_248),
.C(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.C(n_291),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_262),
.B1(n_245),
.B2(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_276),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_274),
.B(n_275),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_191),
.C(n_13),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_13),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_263),
.C(n_270),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_299),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_271),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_291),
.B1(n_271),
.B2(n_280),
.Y(n_309)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_301),
.A2(n_264),
.B1(n_288),
.B2(n_267),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_264),
.C(n_270),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_267),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_310),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_306),
.C(n_302),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_309),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_297),
.B(n_265),
.C(n_293),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_285),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_301),
.B(n_264),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_315),
.A3(n_303),
.B1(n_307),
.B2(n_298),
.C1(n_292),
.C2(n_284),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_318),
.B(n_315),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_312),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_14),
.Y(n_323)
);


endmodule