module fake_jpeg_6320_n_276 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_276);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_15),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_17),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_25),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_33),
.B1(n_26),
.B2(n_17),
.Y(n_47)
);

OAI22x1_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_48),
.B1(n_37),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_17),
.B1(n_13),
.B2(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_17),
.B1(n_32),
.B2(n_14),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_13),
.B1(n_14),
.B2(n_25),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_46),
.B1(n_56),
.B2(n_54),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_40),
.C(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_44),
.B1(n_40),
.B2(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_48),
.B1(n_55),
.B2(n_58),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_40),
.C(n_43),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_49),
.Y(n_87)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_44),
.B1(n_51),
.B2(n_14),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_49),
.B1(n_14),
.B2(n_41),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_62),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_58),
.B1(n_28),
.B2(n_29),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_71),
.B(n_72),
.C(n_75),
.Y(n_97)
);

AOI22x1_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_63),
.B1(n_72),
.B2(n_66),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_69),
.B(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_103),
.B1(n_107),
.B2(n_114),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_93),
.B(n_91),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_63),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_108),
.C(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_71),
.B1(n_69),
.B2(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_60),
.B1(n_51),
.B2(n_57),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_60),
.C(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_89),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_44),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_92),
.A3(n_97),
.B1(n_112),
.B2(n_88),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_92),
.B(n_79),
.C(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_80),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_96),
.B(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_79),
.B1(n_92),
.B2(n_90),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_92),
.B1(n_80),
.B2(n_81),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_92),
.B1(n_94),
.B2(n_42),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_136),
.Y(n_152)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_100),
.C(n_102),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_140),
.C(n_147),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_104),
.C(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_143),
.Y(n_176)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_117),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_101),
.B1(n_113),
.B2(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_121),
.B1(n_158),
.B2(n_115),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_101),
.C(n_78),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_41),
.B1(n_19),
.B2(n_35),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_117),
.B(n_116),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_86),
.C(n_43),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_155),
.C(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_86),
.C(n_94),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_42),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_16),
.B1(n_23),
.B2(n_15),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_121),
.B1(n_129),
.B2(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_166),
.B1(n_177),
.B2(n_18),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_169),
.B(n_149),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_129),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_171),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_121),
.B(n_122),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_99),
.C(n_42),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_178),
.C(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_22),
.B(n_18),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_42),
.C(n_41),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_18),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_199),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_138),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_184),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_19),
.B(n_23),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_156),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_150),
.C(n_139),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_148),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_42),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_24),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_24),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_163),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_41),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_16),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_176),
.B(n_173),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_162),
.B1(n_177),
.B2(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_35),
.C(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_23),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_197),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_35),
.C(n_16),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_35),
.C(n_29),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_190),
.A2(n_11),
.B(n_10),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_228),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_182),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_222),
.B(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_232),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_24),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_202),
.B(n_35),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_208),
.A3(n_216),
.B1(n_205),
.B2(n_209),
.C1(n_215),
.C2(n_214),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_238),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_224),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_239),
.B(n_241),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_218),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_204),
.A3(n_20),
.B1(n_34),
.B2(n_24),
.C1(n_21),
.C2(n_5),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_204),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_244),
.C(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_0),
.C(n_1),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_241),
.C(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_244),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_250),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_1),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_2),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_2),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_3),
.B(n_4),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_3),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_259),
.B(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_261),
.C(n_6),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_4),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_9),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_4),
.C(n_6),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_269),
.B(n_7),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_270),
.B1(n_9),
.B2(n_7),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_6),
.C(n_7),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_6),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_268),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_239),
.C(n_259),
.Y(n_275)
);


endmodule