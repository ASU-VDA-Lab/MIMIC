module fake_jpeg_28253_n_58 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_14),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_10),
.B(n_20),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_8),
.B1(n_19),
.B2(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_22),
.B1(n_23),
.B2(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_32),
.B1(n_7),
.B2(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_5),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_38),
.C(n_41),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_44),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_48),
.B1(n_45),
.B2(n_49),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_55),
.B(n_51),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_53),
.Y(n_58)
);


endmodule