module real_jpeg_22047_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_0),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_84),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_84),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_72),
.B1(n_77),
.B2(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_72),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_74),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_82),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_14),
.B(n_29),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_4),
.A2(n_26),
.B1(n_31),
.B2(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_66),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_66),
.B(n_175),
.Y(n_179)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_8),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_91)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_80),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_40),
.B(n_43),
.C(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_43),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_105),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_52),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_26),
.A2(n_36),
.B1(n_133),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_26),
.A2(n_135),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_27),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_27),
.A2(n_30),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_27),
.A2(n_35),
.B(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_28),
.B(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_91),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_31),
.B(n_78),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_36),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_40),
.A2(n_50),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_40),
.B(n_78),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_40),
.A2(n_50),
.B1(n_143),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_40),
.A2(n_50),
.B1(n_163),
.B2(n_182),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_41),
.A2(n_44),
.B(n_78),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_44),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_43),
.A2(n_67),
.A3(n_70),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_44),
.B(n_64),
.Y(n_176)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_50),
.A2(n_182),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.C(n_75),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_57),
.B(n_60),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_63),
.A2(n_69),
.B1(n_120),
.B2(n_179),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_66),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_80),
.Y(n_89)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_76),
.B1(n_81),
.B2(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_71),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.CON(n_76),
.SN(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_80),
.Y(n_81)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.C(n_111),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_107),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_118),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_200),
.B(n_204),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_187),
.B(n_199),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_169),
.B(n_186),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_155),
.B(n_168),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_144),
.B(n_154),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_136),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_153),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_177),
.B1(n_184),
.B2(n_185),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_183),
.C(n_184),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_189),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_196),
.C(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);


endmodule