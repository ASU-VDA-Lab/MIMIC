module fake_netlist_6_614_n_15 (n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_15);

input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_15;

wire n_7;
wire n_14;
wire n_10;
wire n_13;
wire n_9;
wire n_11;
wire n_8;
wire n_12;

INVx8_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVxp67_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_7),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_10),
.B(n_9),
.Y(n_13)
);

O2A1O1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_7),
.B(n_0),
.C(n_2),
.Y(n_14)
);

BUFx2_ASAP7_75t_SL g15 ( 
.A(n_14),
.Y(n_15)
);


endmodule