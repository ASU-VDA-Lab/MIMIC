module fake_jpeg_28279_n_100 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_53),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_30),
.B(n_24),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_54),
.B(n_55),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_28),
.B1(n_18),
.B2(n_22),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_24),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_14),
.CON(n_56),
.SN(n_56)
);

XOR2x1_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_47),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_33),
.B(n_36),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_58),
.B(n_57),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_62),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_45),
.C(n_46),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_76),
.C(n_39),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_64),
.B(n_63),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_64),
.B1(n_65),
.B2(n_53),
.C(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_45),
.C(n_34),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_77),
.B(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_44),
.C(n_30),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_70),
.B(n_77),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_78),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_42),
.B(n_12),
.C(n_17),
.D(n_75),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_93),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_9),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.C(n_94),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_12),
.B(n_17),
.C(n_4),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_2),
.C(n_4),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_5),
.Y(n_100)
);


endmodule