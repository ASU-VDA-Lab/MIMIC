module fake_jpeg_586_n_502 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_56),
.Y(n_127)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_93),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_26),
.B(n_0),
.CON(n_85),
.SN(n_85)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_85),
.B(n_91),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_88),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

AND2x4_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_98),
.Y(n_164)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_7),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_99),
.B(n_22),
.Y(n_144)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_105),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_43),
.B1(n_37),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_107),
.A2(n_112),
.B1(n_120),
.B2(n_40),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_54),
.A2(n_43),
.B1(n_50),
.B2(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_53),
.A2(n_60),
.B1(n_49),
.B2(n_37),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_49),
.C(n_34),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_20),
.C(n_25),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_22),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_20),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_144),
.B(n_162),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_61),
.A2(n_51),
.B1(n_52),
.B2(n_50),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_148),
.B1(n_167),
.B2(n_16),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_65),
.A2(n_105),
.B1(n_102),
.B2(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_17),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_75),
.B(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_64),
.B(n_45),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_66),
.B(n_25),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_41),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_69),
.A2(n_51),
.B1(n_52),
.B2(n_50),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_71),
.B(n_41),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_70),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_183),
.Y(n_219)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_149),
.B1(n_113),
.B2(n_156),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_74),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_177),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_40),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_39),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_188),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_107),
.A2(n_97),
.B1(n_89),
.B2(n_83),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_184),
.A2(n_201),
.B1(n_206),
.B2(n_164),
.Y(n_238)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_29),
.B1(n_48),
.B2(n_46),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_187),
.A2(n_195),
.B1(n_213),
.B2(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_117),
.B(n_131),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_39),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_194),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_119),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_112),
.A2(n_79),
.B1(n_78),
.B2(n_51),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_207),
.C(n_208),
.Y(n_220)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_127),
.Y(n_200)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_110),
.A2(n_120),
.B1(n_133),
.B2(n_164),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_209),
.B1(n_214),
.B2(n_149),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_132),
.B(n_40),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_116),
.B(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_127),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_209),
.B1(n_200),
.B2(n_172),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_139),
.B(n_42),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_218),
.B1(n_44),
.B2(n_113),
.Y(n_229)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_141),
.C(n_123),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_118),
.A2(n_44),
.B1(n_38),
.B2(n_50),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_16),
.B1(n_34),
.B2(n_36),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_42),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_177),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_226),
.A2(n_243),
.B1(n_252),
.B2(n_208),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_154),
.C(n_158),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_248),
.C(n_208),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_241),
.B1(n_254),
.B2(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_118),
.B1(n_156),
.B2(n_138),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_166),
.B1(n_159),
.B2(n_138),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_177),
.C(n_198),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_180),
.A2(n_29),
.B1(n_48),
.B2(n_46),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_268),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_239),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_238),
.A2(n_184),
.B1(n_190),
.B2(n_211),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_262),
.A2(n_266),
.B1(n_283),
.B2(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_188),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_265),
.Y(n_301)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_185),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_194),
.B1(n_159),
.B2(n_128),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_179),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_274),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_286),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_241),
.A2(n_207),
.B1(n_178),
.B2(n_196),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_278),
.A2(n_202),
.B1(n_199),
.B2(n_150),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_207),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_280),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_232),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_220),
.B(n_231),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_166),
.B1(n_128),
.B2(n_178),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_192),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_287),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_245),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_273),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_253),
.B1(n_226),
.B2(n_236),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_297),
.A2(n_283),
.B1(n_266),
.B2(n_262),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_231),
.B(n_220),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_299),
.A2(n_302),
.B(n_304),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_236),
.B(n_240),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_240),
.B(n_226),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_260),
.A2(n_226),
.A3(n_186),
.B1(n_169),
.B2(n_244),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_266),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_258),
.A2(n_226),
.B(n_214),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_278),
.B(n_277),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_311),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_267),
.B1(n_283),
.B2(n_269),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_224),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.C(n_279),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_230),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_343),
.C(n_315),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_325),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_265),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_327),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_346),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_331),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_291),
.A2(n_277),
.B1(n_278),
.B2(n_261),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_337),
.B1(n_344),
.B2(n_345),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_257),
.B1(n_280),
.B2(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_303),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_339),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_303),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_340),
.A2(n_306),
.B1(n_299),
.B2(n_310),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_275),
.B(n_284),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_230),
.C(n_174),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_227),
.B(n_249),
.C(n_246),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_264),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_360),
.C(n_367),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_292),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_370),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_295),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_365),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_374),
.B1(n_345),
.B2(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_292),
.C(n_306),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_310),
.B1(n_313),
.B2(n_307),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_362),
.A2(n_364),
.B1(n_318),
.B2(n_335),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_337),
.A2(n_298),
.B1(n_290),
.B2(n_311),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_333),
.B(n_294),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_298),
.C(n_203),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_205),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_332),
.C(n_346),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_375),
.C(n_340),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_323),
.A2(n_290),
.B1(n_312),
.B2(n_256),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_204),
.C(n_227),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_348),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_383),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_378),
.A2(n_394),
.B1(n_334),
.B2(n_173),
.Y(n_422)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_369),
.Y(n_383)
);

FAx1_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_339),
.CI(n_345),
.CON(n_384),
.SN(n_384)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_150),
.B(n_191),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_326),
.Y(n_385)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_395),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_342),
.C(n_338),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_387),
.B(n_392),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_393),
.B1(n_397),
.B2(n_399),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_SL g389 ( 
.A(n_359),
.B(n_350),
.C(n_355),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_391),
.Y(n_417)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_331),
.B1(n_320),
.B2(n_319),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_344),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_210),
.C(n_228),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_401),
.Y(n_421)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_228),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_367),
.Y(n_404)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_356),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_357),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_351),
.B(n_249),
.C(n_246),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_334),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_334),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_410),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_347),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_409),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_362),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_356),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_400),
.B(n_356),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_378),
.A2(n_357),
.B1(n_368),
.B2(n_363),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_422),
.B1(n_382),
.B2(n_213),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_389),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_419),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_382),
.B(n_147),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_423),
.A2(n_398),
.B(n_402),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_396),
.C(n_387),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_377),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_434),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_408),
.B(n_384),
.CI(n_386),
.CON(n_427),
.SN(n_427)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_428),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g428 ( 
.A(n_410),
.B(n_423),
.CI(n_409),
.CON(n_428),
.SN(n_428)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_416),
.A2(n_394),
.B1(n_401),
.B2(n_381),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_435),
.A2(n_407),
.B1(n_86),
.B2(n_163),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_411),
.A2(n_175),
.B(n_36),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_437),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_158),
.C(n_237),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_417),
.B(n_415),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_421),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_215),
.B1(n_88),
.B2(n_86),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_439),
.B(n_442),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_424),
.A2(n_237),
.B(n_163),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_406),
.B(n_9),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_420),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_449),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_426),
.A2(n_419),
.B1(n_404),
.B2(n_412),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_446),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_426),
.A2(n_431),
.B1(n_429),
.B2(n_428),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_421),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_450),
.B(n_427),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_451),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_438),
.A2(n_163),
.B(n_1),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_452),
.A2(n_433),
.B(n_440),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_7),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_456),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_436),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_0),
.C(n_3),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_458),
.B(n_0),
.Y(n_464)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_441),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_463),
.Y(n_478)
);

NAND2xp67_ASAP7_75t_SL g463 ( 
.A(n_457),
.B(n_427),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_458),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_466),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_428),
.C(n_5),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_470),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_469),
.A2(n_472),
.B1(n_454),
.B2(n_447),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_445),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_4),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_471),
.B(n_6),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

OAI211xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_483),
.B(n_467),
.C(n_463),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_474),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_462),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_476),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_468),
.A2(n_444),
.B(n_450),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_481),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_484),
.A2(n_486),
.B(n_489),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_473),
.A2(n_466),
.B(n_10),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_6),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_11),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_10),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_493),
.C(n_487),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_485),
.B(n_476),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_494),
.B(n_478),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_496),
.C(n_497),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_478),
.C(n_482),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_11),
.C(n_13),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_11),
.C(n_14),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_14),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_498),
.Y(n_502)
);


endmodule