module fake_netlist_5_655_n_2129 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2129);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2129;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_2031;
wire n_556;
wire n_1728;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_2111;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_2102;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

INVxp33_ASAP7_75t_SL g219 ( 
.A(n_38),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_19),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_148),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_120),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_119),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_113),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_155),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_160),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_21),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_77),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_102),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_60),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_75),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_54),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_159),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_165),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_27),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_136),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_141),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_135),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_81),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_33),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_179),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_66),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_92),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_7),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_65),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_68),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_45),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_156),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_197),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_193),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_86),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_94),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_122),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_111),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_61),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_8),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_147),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_126),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_110),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_138),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_143),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_77),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_161),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_62),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_173),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_163),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_185),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_11),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_44),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_123),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_150),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_169),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_206),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_166),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_153),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_17),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_187),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_58),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_64),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_59),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_82),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_37),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_112),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_149),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_68),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_37),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_158),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_75),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_22),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_101),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_190),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_0),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_188),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_16),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_133),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_130),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_207),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_36),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_90),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_69),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_108),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_54),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_8),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_14),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_43),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_18),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_24),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_3),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_21),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_174),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_208),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_48),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_170),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_74),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_1),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_29),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_4),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_117),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_62),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_131),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_104),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_31),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_66),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_25),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_212),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_105),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_24),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_26),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_42),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_34),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_5),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_64),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_29),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_76),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_184),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_211),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_85),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_96),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_34),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_10),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_56),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_50),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_168),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_132),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_125),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_87),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_1),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_139),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_76),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_3),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_202),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_178),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_5),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_28),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_6),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_13),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_196),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_78),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_36),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_201),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_114),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_6),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_142),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_89),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_55),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_46),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_204),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_38),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_20),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_60),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_199),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_182),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_198),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_115),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_91),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_14),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_47),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_67),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_233),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_0),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_217),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_229),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_229),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_266),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_239),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_239),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_252),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_350),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_288),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_251),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_220),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_252),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_230),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_422),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_2),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_246),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_7),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_254),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_254),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_255),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_271),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_256),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_270),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_265),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_258),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_271),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_272),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_310),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_233),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_288),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_273),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_362),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_288),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_382),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_388),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_286),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_218),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_284),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_288),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_221),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_284),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_R g467 ( 
.A(n_224),
.B(n_84),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_310),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_292),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_293),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_293),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_295),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_297),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_295),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_296),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_296),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_215),
.B(n_12),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_301),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_225),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_270),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_222),
.B(n_13),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_303),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_308),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_309),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_316),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_270),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_227),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_318),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_215),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_301),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_319),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_288),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_304),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_304),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_310),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_306),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_320),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_326),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_306),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_232),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_312),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_312),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_222),
.B(n_15),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_329),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_336),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_313),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_347),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_348),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_313),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_234),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_324),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_236),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_324),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_237),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_335),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_323),
.B(n_15),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_335),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_238),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_338),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_349),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_338),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_351),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_356),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_341),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_243),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_345),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_245),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_248),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_280),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_433),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_370),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_425),
.A2(n_242),
.B1(n_247),
.B2(n_244),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_533),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_433),
.A2(n_458),
.B(n_455),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_458),
.A2(n_372),
.B(n_345),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_464),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_493),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_518),
.B(n_267),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_487),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_487),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_503),
.B(n_323),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_528),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_323),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_280),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_529),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_530),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_505),
.A2(n_328),
.B(n_214),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_R g561 ( 
.A(n_435),
.B(n_219),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_430),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_424),
.B(n_441),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_466),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_472),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_475),
.A2(n_410),
.B(n_372),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_476),
.B(n_399),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_478),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_491),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_481),
.B(n_370),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_497),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_434),
.B(n_278),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_439),
.B(n_450),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_508),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_511),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_513),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_515),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_519),
.A2(n_328),
.B(n_214),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_521),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_523),
.B(n_399),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

AND2x2_ASAP7_75t_SL g602 ( 
.A(n_477),
.B(n_352),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_477),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_447),
.B(n_270),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_461),
.B(n_404),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_423),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_423),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_352),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_435),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_437),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_437),
.B(n_341),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_440),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_440),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_444),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_444),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_446),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g619 ( 
.A(n_428),
.B(n_269),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_446),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_448),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_586),
.B(n_499),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_553),
.B(n_343),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_589),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_538),
.B(n_480),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_589),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_602),
.A2(n_363),
.B1(n_420),
.B2(n_269),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_582),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_557),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_557),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_603),
.B(n_448),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_452),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_542),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_607),
.B(n_486),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_542),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_R g640 ( 
.A(n_620),
.B(n_428),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_603),
.B(n_452),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_612),
.B(n_614),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_553),
.B(n_602),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_607),
.B(n_456),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_539),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_568),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_582),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_542),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_553),
.B(n_602),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_456),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_535),
.B(n_469),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_607),
.B(n_469),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_539),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_604),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_539),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_580),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_582),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_612),
.B(n_462),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_580),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_607),
.B(n_473),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_603),
.B(n_473),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_538),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_603),
.B(n_482),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_580),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_580),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_482),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_552),
.Y(n_669)
);

OR2x2_ASAP7_75t_SL g670 ( 
.A(n_607),
.B(n_410),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_614),
.B(n_615),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_552),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_615),
.B(n_465),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_556),
.B(n_483),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_618),
.B(n_479),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_580),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_543),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_574),
.A2(n_420),
.B1(n_363),
.B2(n_223),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_541),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_541),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_541),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_541),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_611),
.B(n_216),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_543),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_611),
.B(n_357),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_607),
.B(n_483),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_609),
.B(n_276),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_556),
.B(n_484),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_591),
.B(n_485),
.C(n_484),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_591),
.B(n_489),
.C(n_485),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_567),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_607),
.B(n_489),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_543),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_618),
.B(n_488),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_611),
.B(n_357),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_567),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_545),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_607),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_567),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_608),
.B(n_492),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_608),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_545),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_570),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_620),
.B(n_611),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_556),
.B(n_606),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_552),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_608),
.B(n_621),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_581),
.B(n_492),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_606),
.B(n_498),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_620),
.B(n_616),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_582),
.B(n_498),
.Y(n_718)
);

INVx6_ASAP7_75t_L g719 ( 
.A(n_550),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_568),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_609),
.B(n_506),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_621),
.B(n_343),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_562),
.B(n_432),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_570),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_507),
.C(n_506),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_545),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_608),
.B(n_507),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_571),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_571),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_571),
.Y(n_730)
);

BUFx4f_ASAP7_75t_L g731 ( 
.A(n_621),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_616),
.B(n_501),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_572),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_550),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_548),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_548),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_548),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_581),
.B(n_355),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_572),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_608),
.B(n_509),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_552),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_548),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_549),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_572),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_616),
.B(n_512),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_604),
.A2(n_299),
.B1(n_360),
.B2(n_358),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_608),
.B(n_509),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_608),
.B(n_510),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_573),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_608),
.B(n_621),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_550),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_552),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_613),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_574),
.B(n_522),
.C(n_510),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_552),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_581),
.B(n_522),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_621),
.B(n_524),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_609),
.B(n_524),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_613),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_573),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_609),
.B(n_525),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_616),
.B(n_276),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_537),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_605),
.C(n_613),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_609),
.B(n_525),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_549),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_575),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_621),
.B(n_432),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_575),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_537),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_575),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_549),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_609),
.B(n_276),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_640),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_696),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_710),
.B(n_617),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_SL g779 ( 
.A(n_656),
.B(n_449),
.Y(n_779)
);

BUFx4f_ASAP7_75t_L g780 ( 
.A(n_723),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_734),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_624),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_693),
.B(n_617),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_624),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_625),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_633),
.B(n_617),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_722),
.A2(n_609),
.B1(n_223),
.B2(n_226),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_633),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_622),
.B(n_617),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_696),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_717),
.B(n_621),
.Y(n_791)
);

NOR2xp67_ASAP7_75t_L g792 ( 
.A(n_694),
.B(n_605),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_637),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_644),
.B(n_621),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_734),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_641),
.B(n_610),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_753),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_650),
.B(n_609),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_753),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_651),
.B(n_619),
.C(n_561),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_722),
.B(n_711),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_719),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_702),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_731),
.A2(n_547),
.B(n_559),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_634),
.B(n_609),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_755),
.A2(n_561),
.B1(n_516),
.B2(n_520),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_664),
.B(n_589),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_702),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_725),
.B(n_536),
.C(n_619),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_755),
.A2(n_527),
.B1(n_531),
.B2(n_514),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_641),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_652),
.B(n_609),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_658),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_668),
.B(n_609),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_623),
.B(n_547),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_719),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_658),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_705),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_719),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_732),
.B(n_457),
.Y(n_820)
);

AO22x2_ASAP7_75t_L g821 ( 
.A1(n_761),
.A2(n_364),
.B1(n_379),
.B2(n_355),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_731),
.B(n_276),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_663),
.B(n_600),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_663),
.Y(n_824)
);

BUFx6f_ASAP7_75t_SL g825 ( 
.A(n_739),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_623),
.B(n_568),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_642),
.B(n_532),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_623),
.B(n_568),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_671),
.B(n_563),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_761),
.A2(n_460),
.B1(n_459),
.B2(n_302),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_705),
.B(n_568),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_731),
.B(n_276),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_600),
.C(n_590),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_709),
.B(n_568),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_625),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_637),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_721),
.B(n_568),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_709),
.B(n_568),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_716),
.B(n_577),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_716),
.B(n_577),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_665),
.B(n_600),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_724),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_629),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_760),
.B(n_577),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_724),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_714),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_728),
.B(n_577),
.Y(n_848)
);

NAND2x1_ASAP7_75t_L g849 ( 
.A(n_661),
.B(n_550),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_756),
.B(n_536),
.C(n_563),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_629),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_661),
.B(n_550),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_763),
.B(n_577),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_648),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_648),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_728),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_730),
.Y(n_857)
);

INVx8_ASAP7_75t_L g858 ( 
.A(n_685),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_729),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_730),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_659),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_733),
.B(n_577),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_628),
.A2(n_592),
.B(n_595),
.C(n_590),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_733),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_740),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_767),
.B(n_577),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_592),
.Y(n_867)
);

BUFx4f_ASAP7_75t_L g868 ( 
.A(n_723),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_674),
.A2(n_379),
.B1(n_380),
.B2(n_364),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_746),
.B(n_596),
.C(n_595),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_664),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_659),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_740),
.B(n_577),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_692),
.B(n_596),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_688),
.B(n_249),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_660),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_745),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_745),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_718),
.B(n_599),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_747),
.B(n_579),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_627),
.B(n_599),
.C(n_578),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_747),
.B(n_579),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_751),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_751),
.B(n_579),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_762),
.B(n_769),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_762),
.B(n_769),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_771),
.B(n_579),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_771),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_773),
.B(n_579),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_673),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_704),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_714),
.B(n_576),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_773),
.B(n_579),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_713),
.A2(n_559),
.B(n_550),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_628),
.Y(n_895)
);

INVx8_ASAP7_75t_L g896 ( 
.A(n_685),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_635),
.Y(n_897)
);

BUFx5_ASAP7_75t_L g898 ( 
.A(n_666),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_654),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_L g900 ( 
.A(n_688),
.B(n_250),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_635),
.B(n_646),
.Y(n_901)
);

INVxp33_ASAP7_75t_L g902 ( 
.A(n_758),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_704),
.Y(n_903)
);

INVx8_ASAP7_75t_L g904 ( 
.A(n_685),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_707),
.B(n_579),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_758),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_707),
.B(n_579),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_752),
.B(n_585),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_646),
.B(n_585),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_654),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_765),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_765),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_759),
.B(n_231),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_670),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_654),
.B(n_585),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_655),
.B(n_585),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_666),
.B(n_585),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_645),
.B(n_337),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_655),
.B(n_585),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_655),
.B(n_657),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_657),
.B(n_585),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_657),
.B(n_667),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_653),
.B(n_339),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_662),
.B(n_576),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_667),
.B(n_585),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_676),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_L g927 ( 
.A1(n_676),
.A2(n_226),
.B1(n_228),
.B2(n_216),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_690),
.B(n_576),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_765),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_772),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_739),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_739),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_697),
.B(n_578),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_678),
.B(n_594),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_678),
.B(n_594),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_772),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_706),
.A2(n_305),
.B1(n_257),
.B2(n_260),
.Y(n_937)
);

NAND2x1_ASAP7_75t_L g938 ( 
.A(n_680),
.B(n_681),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_680),
.B(n_681),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_682),
.B(n_594),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_682),
.B(n_594),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_727),
.A2(n_311),
.B1(n_262),
.B2(n_264),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_741),
.B(n_578),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_772),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_683),
.B(n_594),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_683),
.B(n_594),
.Y(n_946)
);

OAI21xp33_ASAP7_75t_L g947 ( 
.A1(n_789),
.A2(n_699),
.B(n_675),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_847),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_789),
.B(n_638),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_798),
.A2(n_689),
.B(n_684),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_827),
.B(n_749),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_777),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_786),
.B(n_750),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_778),
.B(n_684),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_851),
.Y(n_955)
);

INVxp33_ASAP7_75t_SL g956 ( 
.A(n_876),
.Y(n_956)
);

CKINVDCx11_ASAP7_75t_R g957 ( 
.A(n_810),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_791),
.A2(n_689),
.B(n_691),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_794),
.A2(n_775),
.B(n_691),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_867),
.B(n_679),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_867),
.B(n_770),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_901),
.A2(n_775),
.B(n_720),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_801),
.A2(n_748),
.B(n_390),
.C(n_380),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_827),
.B(n_626),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_879),
.B(n_688),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_777),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_800),
.A2(n_688),
.B1(n_700),
.B2(n_764),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_939),
.A2(n_559),
.B(n_598),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_804),
.A2(n_598),
.B(n_390),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_939),
.A2(n_922),
.B(n_920),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_781),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_931),
.B(n_932),
.Y(n_972)
);

CKINVDCx8_ASAP7_75t_R g973 ( 
.A(n_782),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_940),
.A2(n_720),
.B(n_647),
.Y(n_974)
);

OAI321xp33_ASAP7_75t_L g975 ( 
.A1(n_869),
.A2(n_322),
.A3(n_325),
.B1(n_330),
.B2(n_331),
.C(n_403),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_781),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_858),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_941),
.A2(n_598),
.B(n_688),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_871),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_788),
.B(n_261),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_941),
.A2(n_700),
.B(n_688),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_785),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_781),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_879),
.B(n_688),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_815),
.A2(n_670),
.B1(n_289),
.B2(n_695),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_790),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_946),
.A2(n_700),
.B(n_631),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_851),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_836),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_796),
.B(n_334),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_813),
.A2(n_720),
.B(n_647),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_817),
.A2(n_647),
.B(n_695),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_811),
.B(n_824),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_946),
.A2(n_700),
.B(n_631),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_787),
.A2(n_712),
.B1(n_742),
.B2(n_695),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_823),
.B(n_334),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_917),
.A2(n_632),
.B(n_630),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_938),
.A2(n_742),
.B(n_712),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_829),
.B(n_700),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_945),
.A2(n_935),
.B(n_925),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_787),
.A2(n_742),
.B1(n_712),
.B2(n_274),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_851),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_913),
.A2(n_700),
.B1(n_764),
.B2(n_275),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_851),
.Y(n_1004)
);

OAI22x1_ASAP7_75t_L g1005 ( 
.A1(n_890),
.A2(n_806),
.B1(n_776),
.B2(n_784),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_803),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_854),
.B(n_558),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_842),
.B(n_892),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_829),
.B(n_700),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_913),
.A2(n_923),
.B(n_918),
.C(n_924),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_874),
.B(n_764),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_902),
.B(n_361),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_915),
.A2(n_672),
.B(n_669),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_906),
.B(n_558),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_820),
.B(n_368),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_874),
.B(n_764),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_918),
.A2(n_279),
.B1(n_281),
.B2(n_277),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_923),
.A2(n_928),
.B(n_924),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_SL g1019 ( 
.A1(n_895),
.A2(n_235),
.B(n_228),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_780),
.B(n_282),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_917),
.A2(n_632),
.B(n_630),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_928),
.B(n_764),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_943),
.B(n_764),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_943),
.B(n_764),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_898),
.B(n_564),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_L g1026 ( 
.A(n_898),
.B(n_283),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_808),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_916),
.A2(n_672),
.B(n_669),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_898),
.B(n_926),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_898),
.B(n_564),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_898),
.B(n_564),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_898),
.B(n_564),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_872),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_807),
.B(n_371),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_926),
.B(n_565),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_780),
.B(n_285),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_783),
.A2(n_863),
.B(n_914),
.C(n_933),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_919),
.A2(n_672),
.B(n_669),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_830),
.B(n_374),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_927),
.A2(n_566),
.B(n_565),
.C(n_593),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_834),
.B(n_290),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_868),
.B(n_375),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_843),
.B(n_565),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_818),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_921),
.A2(n_909),
.B(n_845),
.Y(n_1045)
);

BUFx4f_ASAP7_75t_L g1046 ( 
.A(n_858),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_868),
.B(n_376),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_818),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_934),
.A2(n_636),
.B(n_639),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_933),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_838),
.A2(n_672),
.B(n_669),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_934),
.A2(n_636),
.B(n_639),
.Y(n_1052)
);

CKINVDCx10_ASAP7_75t_R g1053 ( 
.A(n_825),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_838),
.A2(n_672),
.B(n_669),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_781),
.B(n_294),
.Y(n_1055)
);

NAND2x1_ASAP7_75t_L g1056 ( 
.A(n_903),
.B(n_643),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_858),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_845),
.A2(n_754),
.B(n_736),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_897),
.A2(n_298),
.B1(n_307),
.B2(n_314),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_856),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_914),
.A2(n_417),
.B1(n_317),
.B2(n_321),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_859),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_779),
.B(n_377),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_846),
.B(n_565),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_859),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_878),
.B(n_566),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_805),
.A2(n_566),
.B(n_593),
.C(n_588),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_853),
.A2(n_754),
.B(n_736),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_927),
.A2(n_566),
.B(n_593),
.C(n_588),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_854),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_888),
.B(n_569),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_853),
.A2(n_754),
.B(n_736),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_812),
.A2(n_649),
.B(n_643),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_872),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_795),
.B(n_235),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_792),
.B(n_315),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_850),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_881),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_857),
.A2(n_569),
.B(n_593),
.C(n_588),
.Y(n_1080)
);

O2A1O1Ixp5_ASAP7_75t_L g1081 ( 
.A1(n_822),
.A2(n_774),
.B(n_768),
.C(n_649),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_894),
.A2(n_686),
.B(n_677),
.Y(n_1082)
);

OAI21xp33_ASAP7_75t_L g1083 ( 
.A1(n_870),
.A2(n_383),
.B(n_378),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_844),
.B(n_569),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_872),
.B(n_327),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_872),
.B(n_332),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_795),
.B(n_333),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_866),
.A2(n_686),
.B(n_677),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_844),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_866),
.A2(n_698),
.B(n_687),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_825),
.B(n_896),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_797),
.A2(n_799),
.B1(n_816),
.B2(n_802),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_855),
.B(n_569),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_896),
.Y(n_1094)
);

O2A1O1Ixp5_ASAP7_75t_L g1095 ( 
.A1(n_822),
.A2(n_774),
.B(n_768),
.C(n_744),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_814),
.A2(n_353),
.B1(n_387),
.B2(n_389),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_833),
.A2(n_708),
.B(n_744),
.C(n_743),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_849),
.A2(n_852),
.B(n_833),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_809),
.B(n_354),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_855),
.B(n_583),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_861),
.B(n_365),
.Y(n_1101)
);

CKINVDCx10_ASAP7_75t_R g1102 ( 
.A(n_937),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_861),
.B(n_583),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_899),
.B(n_583),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_860),
.B(n_334),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_899),
.B(n_910),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_885),
.A2(n_369),
.B1(n_395),
.B2(n_396),
.Y(n_1107)
);

AO22x1_ASAP7_75t_L g1108 ( 
.A1(n_819),
.A2(n_398),
.B1(n_384),
.B2(n_385),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_942),
.B(n_386),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_826),
.A2(n_698),
.B(n_687),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_864),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_828),
.A2(n_703),
.B(n_701),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_910),
.A2(n_835),
.B(n_832),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_839),
.A2(n_703),
.B(n_701),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_896),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_886),
.A2(n_726),
.B(n_708),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_840),
.A2(n_735),
.B(n_726),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_864),
.B(n_865),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_841),
.A2(n_737),
.B(n_735),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_831),
.B(n_240),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_848),
.A2(n_738),
.B(n_737),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_862),
.A2(n_743),
.B(n_738),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_865),
.B(n_583),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_936),
.B(n_391),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_873),
.A2(n_757),
.B(n_754),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_880),
.A2(n_757),
.B(n_754),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_877),
.A2(n_402),
.B1(n_401),
.B2(n_418),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_882),
.A2(n_887),
.B(n_884),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_877),
.B(n_883),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_883),
.B(n_381),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_891),
.B(n_584),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_911),
.A2(n_584),
.B(n_587),
.C(n_588),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_889),
.A2(n_757),
.B(n_736),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_893),
.A2(n_757),
.B(n_736),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_951),
.A2(n_904),
.B1(n_930),
.B2(n_929),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_982),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_952),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_973),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_1010),
.A2(n_908),
.B(n_944),
.C(n_912),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_955),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_986),
.Y(n_1141)
);

INVx8_ASAP7_75t_L g1142 ( 
.A(n_1075),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_L g1143 ( 
.A1(n_947),
.A2(n_394),
.B(n_393),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1094),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_L g1145 ( 
.A(n_1094),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_966),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_989),
.Y(n_1147)
);

NOR2xp67_ASAP7_75t_SL g1148 ( 
.A(n_971),
.B(n_891),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_979),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1094),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1050),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1008),
.B(n_936),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_964),
.B(n_904),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1018),
.B(n_904),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_960),
.A2(n_908),
.B(n_875),
.C(n_900),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1039),
.A2(n_400),
.B(n_409),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_949),
.A2(n_821),
.B1(n_903),
.B2(n_241),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_961),
.B(n_821),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1026),
.A2(n_903),
.B(n_905),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1078),
.A2(n_397),
.B(n_241),
.C(n_253),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_956),
.B(n_903),
.Y(n_1161)
);

OR2x2_ASAP7_75t_SL g1162 ( 
.A(n_1102),
.B(n_240),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1109),
.A2(n_821),
.B1(n_793),
.B2(n_837),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_977),
.B(n_267),
.Y(n_1164)
);

AO32x1_ASAP7_75t_L g1165 ( 
.A1(n_985),
.A2(n_366),
.A3(n_259),
.B1(n_263),
.B2(n_268),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_955),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_972),
.B(n_392),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1015),
.B(n_412),
.C(n_413),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_954),
.A2(n_1000),
.B(n_1045),
.Y(n_1169)
);

AO21x1_ASAP7_75t_L g1170 ( 
.A1(n_963),
.A2(n_984),
.B(n_965),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1000),
.A2(n_907),
.B(n_905),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1042),
.B(n_907),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_988),
.Y(n_1173)
);

OAI22x1_ASAP7_75t_L g1174 ( 
.A1(n_1064),
.A2(n_421),
.B1(n_340),
.B2(n_359),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1025),
.A2(n_757),
.B(n_587),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1079),
.B(n_584),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1037),
.A2(n_403),
.B1(n_259),
.B2(n_263),
.Y(n_1177)
);

XOR2xp5_ASAP7_75t_L g1178 ( 
.A(n_1005),
.B(n_405),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1048),
.B(n_584),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1083),
.B(n_416),
.C(n_411),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1059),
.B(n_1061),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1063),
.B(n_587),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_999),
.A2(n_287),
.B(n_268),
.C(n_291),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1066),
.B(n_587),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1124),
.A2(n_373),
.B(n_287),
.C(n_291),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1071),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_957),
.Y(n_1187)
);

CKINVDCx14_ASAP7_75t_R g1188 ( 
.A(n_1034),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1006),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1027),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1012),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1030),
.A2(n_601),
.B(n_597),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1099),
.A2(n_300),
.B(n_414),
.C(n_253),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_990),
.B(n_334),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_971),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1031),
.A2(n_601),
.B(n_597),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1115),
.B(n_300),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1118),
.B(n_534),
.Y(n_1198)
);

CKINVDCx14_ASAP7_75t_R g1199 ( 
.A(n_948),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1032),
.A2(n_601),
.B(n_597),
.Y(n_1200)
);

BUFx8_ASAP7_75t_L g1201 ( 
.A(n_1053),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1044),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_972),
.B(n_407),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_953),
.A2(n_397),
.B(n_322),
.C(n_325),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1120),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_988),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1009),
.A2(n_414),
.B(n_340),
.C(n_342),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1111),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1043),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_948),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1065),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1089),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_996),
.B(n_267),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_988),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1067),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1029),
.A2(n_330),
.B1(n_331),
.B2(n_342),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_950),
.A2(n_601),
.B(n_597),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1047),
.B(n_408),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_997),
.A2(n_1052),
.B(n_1088),
.Y(n_1219)
);

AO32x1_ASAP7_75t_L g1220 ( 
.A1(n_1096),
.A2(n_406),
.A3(n_344),
.B1(n_346),
.B2(n_359),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1129),
.A2(n_344),
.B1(n_346),
.B2(n_366),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_SL g1222 ( 
.A1(n_1011),
.A2(n_367),
.B(n_373),
.C(n_406),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_970),
.B(n_534),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1089),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_970),
.A2(n_601),
.B(n_597),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_958),
.A2(n_555),
.B(n_544),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_993),
.B(n_367),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1076),
.B(n_540),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1007),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1014),
.B(n_267),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_971),
.B(n_537),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_971),
.B(n_594),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1105),
.B(n_560),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1088),
.A2(n_551),
.B(n_544),
.Y(n_1234)
);

CKINVDCx8_ASAP7_75t_R g1235 ( 
.A(n_1002),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1076),
.B(n_540),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_974),
.A2(n_959),
.B(n_958),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_959),
.A2(n_991),
.B(n_962),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1007),
.B(n_20),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1128),
.B(n_1113),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_991),
.A2(n_601),
.B(n_597),
.Y(n_1241)
);

AOI221xp5_ASAP7_75t_L g1242 ( 
.A1(n_975),
.A2(n_554),
.B1(n_546),
.B2(n_551),
.C(n_555),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1092),
.A2(n_554),
.B(n_546),
.C(n_560),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_980),
.B(n_23),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1104),
.Y(n_1245)
);

AOI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1128),
.A2(n_601),
.B1(n_597),
.B2(n_594),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1120),
.A2(n_1016),
.B(n_1017),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1019),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1002),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1106),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_977),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1113),
.B(n_560),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1123),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_976),
.B(n_560),
.Y(n_1254)
);

NAND2x1_ASAP7_75t_L g1255 ( 
.A(n_976),
.B(n_549),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1046),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1046),
.B(n_597),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1057),
.B(n_601),
.Y(n_1258)
);

AO21x1_ASAP7_75t_L g1259 ( 
.A1(n_1022),
.A2(n_25),
.B(n_26),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_SL g1260 ( 
.A(n_1057),
.B(n_537),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1131),
.B(n_537),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_1091),
.Y(n_1262)
);

INVx3_ASAP7_75t_SL g1263 ( 
.A(n_1077),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1072),
.B(n_209),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1035),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1041),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1004),
.B(n_205),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1004),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1108),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1004),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1084),
.B(n_200),
.Y(n_1271)
);

AOI221xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1062),
.A2(n_1036),
.B1(n_1020),
.B2(n_1060),
.C(n_1130),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_983),
.B(n_195),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1107),
.A2(n_1055),
.B(n_1086),
.C(n_1085),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1033),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1093),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_R g1277 ( 
.A(n_1033),
.B(n_983),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1033),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1100),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1023),
.A2(n_30),
.B(n_31),
.C(n_35),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_962),
.A2(n_194),
.B(n_189),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1024),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1103),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_967),
.A2(n_40),
.B(n_41),
.C(n_43),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1056),
.B(n_183),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1116),
.B(n_177),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_981),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_992),
.B(n_88),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1101),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_992),
.A2(n_95),
.B(n_171),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_969),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1110),
.B(n_93),
.Y(n_1293)
);

O2A1O1Ixp5_ASAP7_75t_L g1294 ( 
.A1(n_1087),
.A2(n_176),
.B(n_164),
.C(n_162),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_969),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1141),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1191),
.A2(n_1068),
.B(n_1132),
.C(n_1040),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1137),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1148),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1219),
.A2(n_1082),
.B(n_1090),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1172),
.A2(n_1003),
.B(n_1080),
.C(n_1070),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1181),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1169),
.A2(n_1082),
.B(n_1112),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1181),
.Y(n_1304)
);

AOI211x1_ASAP7_75t_L g1305 ( 
.A1(n_1259),
.A2(n_987),
.B(n_994),
.C(n_978),
.Y(n_1305)
);

AOI221x1_ASAP7_75t_L g1306 ( 
.A1(n_1238),
.A2(n_968),
.B1(n_1090),
.B2(n_1074),
.C(n_1112),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1250),
.B(n_1153),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1164),
.A2(n_1262),
.B1(n_1269),
.B2(n_1285),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1149),
.B(n_1001),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1170),
.A2(n_995),
.A3(n_1110),
.B(n_1122),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_SL g1311 ( 
.A1(n_1288),
.A2(n_1021),
.B(n_1049),
.C(n_998),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1189),
.Y(n_1312)
);

OAI222xp33_ASAP7_75t_L g1313 ( 
.A1(n_1282),
.A2(n_1098),
.B1(n_1114),
.B2(n_1117),
.C1(n_1119),
.C2(n_1122),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1152),
.B(n_1114),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1244),
.A2(n_1081),
.B(n_1095),
.C(n_1097),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_998),
.B1(n_1117),
.B2(n_1119),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1146),
.Y(n_1317)
);

OA22x2_ASAP7_75t_L g1318 ( 
.A1(n_1174),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1240),
.A2(n_1155),
.B(n_1237),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1240),
.A2(n_1013),
.B(n_1028),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_1121),
.B(n_1133),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1194),
.B(n_51),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1292),
.A2(n_1121),
.A3(n_1133),
.B(n_1126),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1159),
.A2(n_1223),
.B(n_1252),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1234),
.A2(n_1134),
.B(n_1126),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1195),
.B(n_1058),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1241),
.A2(n_1134),
.B(n_1125),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1225),
.A2(n_1125),
.B(n_1038),
.Y(n_1328)
);

NOR4xp25_ASAP7_75t_L g1329 ( 
.A(n_1282),
.B(n_52),
.C(n_55),
.D(n_56),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1190),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1223),
.A2(n_1069),
.B(n_1054),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1202),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1252),
.A2(n_1051),
.B(n_1073),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1152),
.B(n_57),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_SL g1335 ( 
.A1(n_1284),
.A2(n_106),
.B(n_146),
.C(n_145),
.Y(n_1335)
);

CKINVDCx12_ASAP7_75t_R g1336 ( 
.A(n_1142),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1209),
.B(n_63),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1211),
.B(n_65),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1171),
.A2(n_100),
.B(n_137),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1287),
.A2(n_151),
.B(n_99),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1289),
.A2(n_1287),
.B(n_1139),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1208),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1158),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1215),
.B(n_70),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1226),
.A2(n_1217),
.B(n_1289),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1176),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1213),
.B(n_71),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1210),
.B(n_116),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1177),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.C(n_74),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1293),
.A2(n_129),
.B(n_109),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1293),
.A2(n_118),
.B(n_127),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1177),
.A2(n_72),
.A3(n_73),
.B(n_128),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1147),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1176),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1228),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1276),
.B(n_1283),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1158),
.A2(n_1247),
.B(n_1175),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1247),
.A2(n_1271),
.B(n_1264),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1157),
.A2(n_1185),
.A3(n_1248),
.B(n_1216),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1229),
.B(n_1239),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1228),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1186),
.B(n_1236),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1233),
.Y(n_1363)
);

NOR4xp25_ASAP7_75t_L g1364 ( 
.A(n_1280),
.B(n_1290),
.C(n_1266),
.D(n_1160),
.Y(n_1364)
);

AOI31xp67_ASAP7_75t_L g1365 ( 
.A1(n_1271),
.A2(n_1264),
.A3(n_1135),
.B(n_1198),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1179),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1279),
.B(n_1265),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1157),
.A2(n_1216),
.A3(n_1243),
.B(n_1196),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_SL g1369 ( 
.A1(n_1267),
.A2(n_1257),
.B(n_1258),
.C(n_1274),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1236),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1246),
.A2(n_1200),
.B(n_1192),
.Y(n_1371)
);

AOI211x1_ASAP7_75t_L g1372 ( 
.A1(n_1143),
.A2(n_1156),
.B(n_1221),
.C(n_1168),
.Y(n_1372)
);

AOI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1179),
.A2(n_1184),
.B(n_1182),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1218),
.A2(n_1295),
.B(n_1230),
.C(n_1161),
.Y(n_1374)
);

AOI221xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1221),
.A2(n_1204),
.B1(n_1193),
.B2(n_1163),
.C(n_1242),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1182),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1198),
.A2(n_1261),
.B(n_1281),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1261),
.A2(n_1260),
.B(n_1253),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1256),
.B(n_1144),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1184),
.A2(n_1291),
.A3(n_1245),
.B(n_1227),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1136),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1235),
.A2(n_1278),
.B1(n_1145),
.B2(n_1180),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1232),
.A2(n_1222),
.B(n_1207),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1255),
.A2(n_1286),
.B(n_1231),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1138),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1294),
.A2(n_1183),
.B(n_1272),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1254),
.A2(n_1203),
.B(n_1167),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1242),
.A2(n_1224),
.B(n_1212),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1165),
.A2(n_1220),
.A3(n_1249),
.B(n_1286),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1254),
.A2(n_1197),
.B(n_1178),
.Y(n_1390)
);

AOI221xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1166),
.A2(n_1268),
.B1(n_1173),
.B2(n_1206),
.C(n_1165),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1231),
.A2(n_1273),
.B(n_1140),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1197),
.A2(n_1205),
.B1(n_1263),
.B2(n_1199),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1165),
.A2(n_1220),
.B(n_1251),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1145),
.A2(n_1273),
.B(n_1140),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1220),
.A2(n_1151),
.A3(n_1214),
.B(n_1270),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1144),
.B(n_1150),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1187),
.A2(n_1142),
.B1(n_1144),
.B2(n_1150),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1275),
.A2(n_1277),
.A3(n_1173),
.B(n_1268),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1136),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1275),
.A2(n_1162),
.B(n_1142),
.C(n_1150),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1166),
.A2(n_1173),
.B(n_1206),
.C(n_1268),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1166),
.Y(n_1403)
);

AO32x2_ASAP7_75t_L g1404 ( 
.A1(n_1206),
.A2(n_1157),
.A3(n_1177),
.B1(n_1282),
.B2(n_1216),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1201),
.A2(n_1259),
.B(n_1274),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1201),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_SL g1407 ( 
.A(n_1187),
.B(n_973),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1191),
.B(n_876),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1237),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1172),
.A2(n_1010),
.B(n_752),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1158),
.A2(n_1010),
.B1(n_960),
.B2(n_789),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1172),
.A2(n_951),
.B(n_1010),
.C(n_947),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1172),
.A2(n_951),
.B(n_1010),
.C(n_947),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1158),
.A2(n_1010),
.B1(n_960),
.B2(n_789),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1282),
.A2(n_1010),
.B1(n_927),
.B2(n_1018),
.C(n_947),
.Y(n_1416)
);

AO21x1_ASAP7_75t_L g1417 ( 
.A1(n_1177),
.A2(n_1018),
.B(n_949),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1170),
.A2(n_1292),
.A3(n_1240),
.B(n_1238),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1147),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1288),
.A2(n_1010),
.B(n_1018),
.C(n_960),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1191),
.B(n_876),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1141),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1425)
);

AOI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1174),
.A2(n_591),
.B1(n_947),
.B2(n_951),
.C(n_827),
.Y(n_1426)
);

AO21x1_ASAP7_75t_L g1427 ( 
.A1(n_1177),
.A2(n_1018),
.B(n_949),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1237),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1194),
.B(n_902),
.Y(n_1429)
);

O2A1O1Ixp5_ASAP7_75t_L g1430 ( 
.A1(n_1170),
.A2(n_1010),
.B(n_951),
.C(n_1018),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1285),
.A2(n_951),
.B1(n_947),
.B2(n_809),
.Y(n_1432)
);

AOI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1158),
.A2(n_1293),
.B(n_960),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1237),
.Y(n_1434)
);

AO31x2_ASAP7_75t_L g1435 ( 
.A1(n_1170),
.A2(n_1292),
.A3(n_1240),
.B(n_1238),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1172),
.A2(n_951),
.B(n_1010),
.C(n_947),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1237),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1201),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1145),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1172),
.A2(n_951),
.B(n_1010),
.C(n_947),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1147),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1154),
.A2(n_1226),
.B(n_1225),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1446)
);

AO32x2_ASAP7_75t_L g1447 ( 
.A1(n_1157),
.A2(n_1177),
.A3(n_1282),
.B1(n_1216),
.B2(n_1221),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1237),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1191),
.B(n_789),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_SL g1450 ( 
.A(n_1164),
.B(n_890),
.C(n_876),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1169),
.A2(n_1010),
.B(n_1018),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1169),
.A2(n_731),
.B(n_791),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1191),
.A2(n_1010),
.B(n_947),
.C(n_951),
.Y(n_1453)
);

NOR3xp33_ASAP7_75t_L g1454 ( 
.A(n_1168),
.B(n_951),
.C(n_947),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1147),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1195),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1250),
.B(n_789),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1195),
.Y(n_1458)
);

AOI221x1_ASAP7_75t_L g1459 ( 
.A1(n_1238),
.A2(n_1010),
.B1(n_947),
.B2(n_1018),
.C(n_951),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1169),
.A2(n_1010),
.B(n_1018),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_SL g1461 ( 
.A(n_1164),
.B(n_890),
.C(n_876),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1385),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1454),
.A2(n_1426),
.B1(n_1432),
.B2(n_1427),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1439),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_1439),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1296),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_1439),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1353),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1417),
.B1(n_1343),
.B2(n_1411),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1318),
.A2(n_1343),
.B1(n_1415),
.B2(n_1411),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1438),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1381),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1415),
.A2(n_1309),
.B1(n_1460),
.B2(n_1451),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1420),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1405),
.A2(n_1461),
.B1(n_1450),
.B2(n_1408),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1322),
.A2(n_1347),
.B1(n_1350),
.B2(n_1340),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1350),
.A2(n_1340),
.B1(n_1460),
.B2(n_1451),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1298),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1308),
.A2(n_1422),
.B(n_1349),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1455),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1355),
.A2(n_1370),
.B1(n_1361),
.B2(n_1449),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1379),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1400),
.Y(n_1484)
);

OAI21xp33_ASAP7_75t_L g1485 ( 
.A1(n_1412),
.A2(n_1436),
.B(n_1413),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1317),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1406),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1360),
.A2(n_1329),
.B1(n_1344),
.B2(n_1337),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1423),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1407),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1344),
.A2(n_1338),
.B1(n_1363),
.B2(n_1457),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1302),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1429),
.Y(n_1493)
);

BUFx2_ASAP7_75t_SL g1494 ( 
.A(n_1348),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1329),
.A2(n_1393),
.B1(n_1336),
.B2(n_1372),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1397),
.Y(n_1496)
);

CKINVDCx6p67_ASAP7_75t_R g1497 ( 
.A(n_1334),
.Y(n_1497)
);

CKINVDCx6p67_ASAP7_75t_R g1498 ( 
.A(n_1334),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1312),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_SL g1500 ( 
.A(n_1403),
.Y(n_1500)
);

BUFx2_ASAP7_75t_SL g1501 ( 
.A(n_1382),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1330),
.Y(n_1502)
);

CKINVDCx11_ASAP7_75t_R g1503 ( 
.A(n_1382),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1399),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1457),
.A2(n_1304),
.B1(n_1356),
.B2(n_1354),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1440),
.A2(n_1367),
.B1(n_1453),
.B2(n_1346),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1332),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1358),
.A2(n_1342),
.B1(n_1386),
.B2(n_1341),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1396),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1386),
.A2(n_1314),
.B1(n_1366),
.B2(n_1376),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1396),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1399),
.Y(n_1512)
);

BUFx8_ASAP7_75t_L g1513 ( 
.A(n_1404),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1316),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1314),
.A2(n_1351),
.B1(n_1357),
.B2(n_1387),
.Y(n_1515)
);

CKINVDCx11_ASAP7_75t_R g1516 ( 
.A(n_1398),
.Y(n_1516)
);

INVx6_ASAP7_75t_L g1517 ( 
.A(n_1399),
.Y(n_1517)
);

CKINVDCx11_ASAP7_75t_R g1518 ( 
.A(n_1390),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1326),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1396),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1456),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1459),
.A2(n_1388),
.B1(n_1447),
.B2(n_1299),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1402),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1401),
.A2(n_1339),
.B(n_1301),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1326),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1456),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1458),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1395),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1357),
.A2(n_1388),
.B1(n_1394),
.B2(n_1447),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1352),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1352),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1458),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1319),
.A2(n_1324),
.B1(n_1378),
.B2(n_1345),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1392),
.Y(n_1535)
);

BUFx5_ASAP7_75t_L g1536 ( 
.A(n_1313),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1352),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_L g1538 ( 
.A(n_1374),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1364),
.A2(n_1410),
.B(n_1297),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1419),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1384),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1305),
.A2(n_1383),
.B1(n_1315),
.B2(n_1377),
.Y(n_1542)
);

CKINVDCx6p67_ASAP7_75t_R g1543 ( 
.A(n_1335),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1404),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1414),
.A2(n_1444),
.B1(n_1418),
.B2(n_1452),
.Y(n_1545)
);

CKINVDCx11_ASAP7_75t_R g1546 ( 
.A(n_1364),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1375),
.A2(n_1303),
.B1(n_1430),
.B2(n_1404),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1435),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1433),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_SL g1550 ( 
.A(n_1369),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1424),
.A2(n_1431),
.B1(n_1446),
.B2(n_1445),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1375),
.A2(n_1311),
.B1(n_1320),
.B2(n_1331),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1333),
.A2(n_1425),
.B1(n_1443),
.B2(n_1359),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1373),
.A2(n_1306),
.B1(n_1442),
.B2(n_1321),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1365),
.A2(n_1380),
.B1(n_1368),
.B2(n_1391),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1409),
.A2(n_1448),
.B1(n_1437),
.B2(n_1434),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1428),
.A2(n_1327),
.B1(n_1328),
.B2(n_1325),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1391),
.A2(n_1368),
.B1(n_1371),
.B2(n_1300),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1380),
.B(n_1368),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1380),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1323),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1389),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1389),
.A2(n_604),
.B1(n_820),
.B2(n_1318),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1310),
.A2(n_1426),
.B1(n_951),
.B2(n_947),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1389),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1310),
.A2(n_1426),
.B1(n_951),
.B2(n_947),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_947),
.B2(n_1018),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1385),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1439),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_947),
.B2(n_1018),
.Y(n_1570)
);

BUFx4_ASAP7_75t_R g1571 ( 
.A(n_1400),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1419),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1439),
.Y(n_1574)
);

BUFx10_ASAP7_75t_L g1575 ( 
.A(n_1439),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1298),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_876),
.B2(n_890),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_947),
.B2(n_1018),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1432),
.A2(n_890),
.B1(n_876),
.B2(n_827),
.Y(n_1579)
);

BUFx8_ASAP7_75t_L g1580 ( 
.A(n_1438),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_947),
.B2(n_1018),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1298),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1439),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1298),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1296),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1296),
.Y(n_1588)
);

BUFx10_ASAP7_75t_L g1589 ( 
.A(n_1439),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1296),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1426),
.A2(n_951),
.B1(n_947),
.B2(n_1018),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1296),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1298),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1298),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1420),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1298),
.Y(n_1596)
);

OAI22x1_ASAP7_75t_L g1597 ( 
.A1(n_1390),
.A2(n_951),
.B1(n_876),
.B2(n_890),
.Y(n_1597)
);

BUFx8_ASAP7_75t_L g1598 ( 
.A(n_1438),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1420),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1439),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1412),
.A2(n_1436),
.B(n_1413),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1349),
.A2(n_1318),
.B1(n_820),
.B2(n_1426),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1385),
.Y(n_1605)
);

OAI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1349),
.A2(n_1318),
.B1(n_820),
.B2(n_1426),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1362),
.B(n_1307),
.Y(n_1607)
);

INVx6_ASAP7_75t_L g1608 ( 
.A(n_1439),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1318),
.A2(n_604),
.B1(n_820),
.B2(n_656),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1385),
.Y(n_1610)
);

CKINVDCx11_ASAP7_75t_R g1611 ( 
.A(n_1610),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1579),
.A2(n_1577),
.B1(n_1597),
.B2(n_1480),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1542),
.A2(n_1551),
.B(n_1545),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1556),
.A2(n_1557),
.B(n_1553),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1481),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1544),
.B(n_1531),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1466),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1544),
.B(n_1474),
.Y(n_1618)
);

BUFx12f_ASAP7_75t_L g1619 ( 
.A(n_1490),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1532),
.Y(n_1620)
);

AOI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1537),
.A2(n_1555),
.B(n_1559),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1544),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1504),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1489),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1544),
.B(n_1474),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1535),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1574),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1567),
.A2(n_1570),
.B(n_1578),
.C(n_1591),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1541),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1541),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1540),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1567),
.A2(n_1578),
.B(n_1570),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1556),
.A2(n_1553),
.B(n_1534),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1546),
.A2(n_1514),
.B1(n_1477),
.B2(n_1591),
.Y(n_1636)
);

OR2x6_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1519),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1468),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1512),
.B(n_1587),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1482),
.B(n_1491),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1548),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1472),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1534),
.A2(n_1508),
.B(n_1552),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1588),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1560),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1533),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1590),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1462),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1533),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1592),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1482),
.B(n_1491),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1499),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1547),
.B(n_1530),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1530),
.A2(n_1508),
.B(n_1547),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1470),
.B(n_1563),
.Y(n_1655)
);

OAI21xp33_ASAP7_75t_SL g1656 ( 
.A1(n_1581),
.A2(n_1492),
.B(n_1463),
.Y(n_1656)
);

BUFx12f_ASAP7_75t_L g1657 ( 
.A(n_1568),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1502),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1507),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1605),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1492),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1479),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1486),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1554),
.A2(n_1522),
.B(n_1539),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1517),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1571),
.Y(n_1666)
);

BUFx2_ASAP7_75t_SL g1667 ( 
.A(n_1528),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1509),
.A2(n_1520),
.B(n_1511),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1573),
.B(n_1529),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1576),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1573),
.B(n_1565),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1583),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1515),
.A2(n_1562),
.B(n_1510),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1561),
.Y(n_1674)
);

AOI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1506),
.A2(n_1523),
.B(n_1594),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1525),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1505),
.B(n_1581),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1477),
.A2(n_1478),
.B1(n_1485),
.B2(n_1495),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1517),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1585),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1593),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1596),
.Y(n_1682)
);

AO32x2_ASAP7_75t_L g1683 ( 
.A1(n_1488),
.A2(n_1513),
.A3(n_1522),
.B1(n_1536),
.B2(n_1604),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1561),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1470),
.B(n_1563),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1488),
.B(n_1469),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1513),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1518),
.A2(n_1498),
.B1(n_1497),
.B2(n_1501),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1505),
.B(n_1609),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1572),
.A2(n_1609),
.B1(n_1599),
.B2(n_1586),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1515),
.A2(n_1510),
.B(n_1524),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1572),
.B(n_1582),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1536),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1536),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1469),
.B(n_1536),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1517),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1536),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1483),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1582),
.B(n_1586),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1536),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1550),
.Y(n_1701)
);

AO31x2_ASAP7_75t_L g1702 ( 
.A1(n_1558),
.A2(n_1554),
.A3(n_1606),
.B(n_1604),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1550),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1549),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1493),
.Y(n_1705)
);

O2A1O1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1606),
.A2(n_1564),
.B(n_1566),
.C(n_1476),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1558),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1521),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1538),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1538),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1543),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1527),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1493),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1599),
.B(n_1601),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1608),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1595),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1496),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1526),
.A2(n_1601),
.B(n_1600),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1494),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1500),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1503),
.A2(n_1500),
.B(n_1487),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1487),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1580),
.Y(n_1723)
);

AO21x1_ASAP7_75t_SL g1724 ( 
.A1(n_1516),
.A2(n_1465),
.B(n_1467),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1635),
.A2(n_1569),
.B(n_1584),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1615),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1615),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1706),
.A2(n_1608),
.B(n_1465),
.C(n_1467),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1612),
.B(n_1464),
.Y(n_1729)
);

OR2x6_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1475),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1668),
.Y(n_1731)
);

OAI31xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1634),
.A2(n_1473),
.A3(n_1580),
.B(n_1598),
.Y(n_1732)
);

AND2x6_ASAP7_75t_L g1733 ( 
.A(n_1655),
.B(n_1685),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1629),
.A2(n_1471),
.B(n_1589),
.C(n_1575),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1692),
.A2(n_1602),
.B(n_1484),
.C(n_1598),
.Y(n_1735)
);

O2A1O1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1699),
.A2(n_1656),
.B(n_1677),
.C(n_1678),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_1611),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1689),
.B(n_1640),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1690),
.A2(n_1714),
.B(n_1636),
.C(n_1686),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1632),
.B(n_1713),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1651),
.B(n_1718),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1713),
.B(n_1618),
.Y(n_1743)
);

AO32x2_ASAP7_75t_L g1744 ( 
.A1(n_1665),
.A2(n_1696),
.A3(n_1683),
.B1(n_1664),
.B2(n_1616),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1618),
.B(n_1625),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_SL g1746 ( 
.A1(n_1711),
.A2(n_1703),
.B(n_1701),
.C(n_1710),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1625),
.B(n_1705),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1616),
.B(n_1669),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1637),
.A2(n_1643),
.B(n_1691),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1675),
.B(n_1688),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_SL g1751 ( 
.A1(n_1711),
.A2(n_1710),
.B(n_1709),
.C(n_1719),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1695),
.B(n_1687),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1676),
.Y(n_1753)
);

BUFx4f_ASAP7_75t_SL g1754 ( 
.A(n_1657),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1718),
.B(n_1714),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1686),
.A2(n_1643),
.B(n_1655),
.C(n_1685),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1718),
.B(n_1667),
.Y(n_1757)
);

INVx4_ASAP7_75t_L g1758 ( 
.A(n_1676),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1693),
.A2(n_1694),
.B(n_1697),
.C(n_1700),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1637),
.A2(n_1664),
.B(n_1693),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1695),
.B(n_1687),
.Y(n_1761)
);

BUFx8_ASAP7_75t_SL g1762 ( 
.A(n_1723),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1648),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1676),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1637),
.A2(n_1721),
.B(n_1718),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1668),
.Y(n_1766)
);

OAI21xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1709),
.A2(n_1719),
.B(n_1661),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1668),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1638),
.B(n_1642),
.Y(n_1769)
);

AO32x2_ASAP7_75t_L g1770 ( 
.A1(n_1665),
.A2(n_1696),
.A3(n_1683),
.B1(n_1664),
.B2(n_1668),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_R g1771 ( 
.A(n_1666),
.B(n_1723),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1720),
.A2(n_1717),
.B(n_1722),
.C(n_1698),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1673),
.A2(n_1614),
.B(n_1613),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1669),
.B(n_1694),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1666),
.A2(n_1704),
.B1(n_1717),
.B2(n_1721),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1644),
.B(n_1647),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1620),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1704),
.A2(n_1722),
.B(n_1716),
.C(n_1712),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1653),
.A2(n_1707),
.B1(n_1659),
.B2(n_1617),
.C(n_1658),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_1619),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_R g1782 ( 
.A(n_1721),
.B(n_1654),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1650),
.B(n_1652),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1675),
.B(n_1679),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1624),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1623),
.B(n_1627),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1620),
.Y(n_1787)
);

AO32x2_ASAP7_75t_L g1788 ( 
.A1(n_1683),
.A2(n_1698),
.A3(n_1702),
.B1(n_1649),
.B2(n_1646),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1662),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1633),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1627),
.B(n_1630),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1671),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1630),
.B(n_1631),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1671),
.B(n_1645),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1613),
.A2(n_1614),
.B(n_1621),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1641),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1787),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1791),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1745),
.B(n_1707),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1777),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1790),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1738),
.B(n_1672),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1796),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1738),
.B(n_1670),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1755),
.B(n_1683),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1755),
.B(n_1683),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1752),
.B(n_1673),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1761),
.B(n_1743),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1758),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1771),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1747),
.B(n_1621),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1767),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1744),
.B(n_1654),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1786),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1792),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1792),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_SL g1817 ( 
.A1(n_1733),
.A2(n_1721),
.B1(n_1619),
.B2(n_1654),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1731),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1748),
.B(n_1774),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1726),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1794),
.B(n_1742),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1791),
.Y(n_1822)
);

OAI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1736),
.A2(n_1680),
.B1(n_1682),
.B2(n_1681),
.C1(n_1663),
.C2(n_1708),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1769),
.B(n_1702),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1741),
.B(n_1742),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1766),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1766),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1744),
.B(n_1684),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1744),
.B(n_1739),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1789),
.B(n_1702),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1768),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1785),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1756),
.B(n_1702),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1770),
.B(n_1674),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1776),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1779),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1756),
.B(n_1702),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1781),
.B(n_1720),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1783),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1770),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1829),
.B(n_1770),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1812),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1834),
.B(n_1793),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1840),
.B(n_1821),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1829),
.B(n_1770),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1834),
.B(n_1725),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1821),
.B(n_1757),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1813),
.B(n_1773),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1818),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1833),
.A2(n_1837),
.B1(n_1733),
.B2(n_1806),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1818),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1826),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1828),
.B(n_1759),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1812),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1828),
.B(n_1759),
.Y(n_1855)
);

NAND2x1p5_ASAP7_75t_SL g1856 ( 
.A(n_1805),
.B(n_1750),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1795),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1827),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1806),
.A2(n_1733),
.B1(n_1729),
.B2(n_1757),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1831),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1807),
.B(n_1795),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1807),
.B(n_1760),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1811),
.B(n_1788),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_R g1864 ( 
.A(n_1810),
.B(n_1737),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1811),
.B(n_1788),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1815),
.B(n_1749),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1816),
.B(n_1780),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1797),
.Y(n_1868)
);

OAI31xp33_ASAP7_75t_L g1869 ( 
.A1(n_1823),
.A2(n_1740),
.A3(n_1734),
.B(n_1736),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1830),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1800),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1797),
.Y(n_1872)
);

NOR2x1_ASAP7_75t_SL g1873 ( 
.A(n_1800),
.B(n_1784),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1824),
.A2(n_1740),
.B1(n_1734),
.B2(n_1750),
.C(n_1729),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1870),
.B(n_1825),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1868),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1842),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1849),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1870),
.B(n_1835),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1851),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_R g1881 ( 
.A(n_1842),
.B(n_1754),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1851),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1841),
.B(n_1808),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1846),
.B(n_1808),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1867),
.B(n_1836),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1868),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1873),
.B(n_1798),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1842),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1842),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1841),
.B(n_1845),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1891)
);

INVx4_ASAP7_75t_L g1892 ( 
.A(n_1854),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1849),
.Y(n_1893)
);

OA21x2_ASAP7_75t_L g1894 ( 
.A1(n_1848),
.A2(n_1803),
.B(n_1801),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1873),
.B(n_1822),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1841),
.B(n_1814),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1874),
.B(n_1817),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1845),
.B(n_1814),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1854),
.Y(n_1899)
);

NAND2x1_ASAP7_75t_L g1900 ( 
.A(n_1860),
.B(n_1765),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1852),
.Y(n_1902)
);

AND2x4_ASAP7_75t_SL g1903 ( 
.A(n_1843),
.B(n_1730),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1845),
.B(n_1799),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1853),
.B(n_1799),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1867),
.B(n_1836),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1854),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1846),
.B(n_1839),
.Y(n_1908)
);

OR2x2_ASAP7_75t_SL g1909 ( 
.A(n_1847),
.B(n_1802),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1853),
.B(n_1839),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1872),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1858),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1871),
.B(n_1832),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1872),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1854),
.B(n_1804),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1880),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1877),
.B(n_1873),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_SL g1918 ( 
.A(n_1892),
.B(n_1869),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1880),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_L g1920 ( 
.A(n_1897),
.B(n_1881),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1882),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1882),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1883),
.B(n_1853),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1915),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1902),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1894),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1892),
.B(n_1730),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1877),
.B(n_1866),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1894),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1902),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1910),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1915),
.B(n_1874),
.Y(n_1932)
);

CKINVDCx16_ASAP7_75t_R g1933 ( 
.A(n_1881),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1910),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1910),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1885),
.B(n_1847),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1909),
.B(n_1875),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1892),
.B(n_1869),
.Y(n_1938)
);

OAI21xp33_ASAP7_75t_L g1939 ( 
.A1(n_1897),
.A2(n_1850),
.B(n_1859),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1913),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1913),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1905),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1905),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1892),
.B(n_1730),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1885),
.B(n_1850),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1905),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1889),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1909),
.B(n_1856),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1889),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1906),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1883),
.B(n_1855),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1889),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1883),
.B(n_1855),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1891),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1909),
.B(n_1856),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1906),
.B(n_1855),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1891),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1891),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1908),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1884),
.B(n_1862),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1884),
.B(n_1890),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1899),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1908),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1894),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1875),
.B(n_1856),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1920),
.A2(n_1900),
.B(n_1732),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1961),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1916),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1949),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1961),
.B(n_1877),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1932),
.B(n_1924),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1949),
.B(n_1877),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1916),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1939),
.B(n_1857),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1923),
.B(n_1892),
.Y(n_1975)
);

NAND2x1_ASAP7_75t_L g1976 ( 
.A(n_1917),
.B(n_1892),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1945),
.B(n_1857),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1956),
.B(n_1879),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1947),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1933),
.B(n_1762),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1923),
.B(n_1890),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1918),
.B(n_1762),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1938),
.B(n_1754),
.Y(n_1983)
);

OAI21xp33_ASAP7_75t_L g1984 ( 
.A1(n_1920),
.A2(n_1955),
.B(n_1948),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1965),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1951),
.B(n_1953),
.Y(n_1986)
);

NOR2xp67_ASAP7_75t_L g1987 ( 
.A(n_1917),
.B(n_1888),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1919),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1921),
.Y(n_1989)
);

NOR3xp33_ASAP7_75t_L g1990 ( 
.A(n_1952),
.B(n_1735),
.C(n_1838),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1951),
.B(n_1890),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1953),
.B(n_1899),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1928),
.Y(n_1993)
);

NAND4xp25_ASAP7_75t_L g1994 ( 
.A(n_1937),
.B(n_1859),
.C(n_1735),
.D(n_1907),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1942),
.B(n_1879),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1922),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1960),
.B(n_1899),
.Y(n_1997)
);

INVxp33_ASAP7_75t_L g1998 ( 
.A(n_1936),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1960),
.B(n_1899),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1928),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1950),
.B(n_1857),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1928),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1925),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1962),
.B(n_1861),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1954),
.B(n_1861),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1943),
.B(n_1856),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1972),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1982),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1983),
.A2(n_1958),
.B1(n_1957),
.B2(n_1946),
.Y(n_2009)
);

OAI32xp33_ASAP7_75t_L g2010 ( 
.A1(n_1984),
.A2(n_1965),
.A3(n_1907),
.B1(n_1930),
.B2(n_1888),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1981),
.B(n_1907),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1979),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1984),
.B(n_1940),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1981),
.B(n_1907),
.Y(n_2014)
);

OAI211xp5_ASAP7_75t_L g2015 ( 
.A1(n_1974),
.A2(n_1966),
.B(n_1994),
.C(n_1971),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1969),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1985),
.B(n_1941),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1980),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1990),
.A2(n_1888),
.B(n_1900),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1972),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1969),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1993),
.Y(n_2022)
);

OAI332xp33_ASAP7_75t_L g2023 ( 
.A1(n_1968),
.A2(n_1888),
.A3(n_1929),
.B1(n_1926),
.B2(n_1964),
.B3(n_1931),
.C1(n_1934),
.C2(n_1935),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1968),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1991),
.B(n_1917),
.Y(n_2025)
);

AOI222xp33_ASAP7_75t_L g2026 ( 
.A1(n_1998),
.A2(n_1733),
.B1(n_1963),
.B2(n_1959),
.C1(n_1865),
.C2(n_1863),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1973),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1988),
.B(n_1657),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1973),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1986),
.B(n_1862),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_1977),
.A2(n_1900),
.B1(n_1929),
.B2(n_1926),
.C(n_1964),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1988),
.B(n_1763),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_1989),
.A2(n_1861),
.B1(n_1862),
.B2(n_1895),
.C(n_1887),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1986),
.B(n_1884),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1991),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_L g2036 ( 
.A(n_1989),
.B(n_1775),
.C(n_1778),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2024),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2027),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_2007),
.Y(n_2039)
);

INVxp67_ASAP7_75t_L g2040 ( 
.A(n_2032),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2018),
.A2(n_1992),
.B1(n_1975),
.B2(n_1967),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2029),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2035),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2016),
.B(n_1992),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_2007),
.B(n_1987),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2021),
.B(n_2002),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2025),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2010),
.A2(n_2003),
.B(n_1996),
.C(n_1987),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_2010),
.A2(n_1996),
.B1(n_2003),
.B2(n_2001),
.C(n_1972),
.Y(n_2050)
);

AOI21xp33_ASAP7_75t_L g2051 ( 
.A1(n_2015),
.A2(n_1976),
.B(n_2000),
.Y(n_2051)
);

AOI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_2013),
.A2(n_1978),
.B1(n_2000),
.B2(n_2004),
.C(n_1967),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2008),
.B(n_1997),
.Y(n_2053)
);

CKINVDCx16_ASAP7_75t_R g2054 ( 
.A(n_2032),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2028),
.A2(n_1999),
.B1(n_1997),
.B2(n_1975),
.Y(n_2055)
);

INVxp67_ASAP7_75t_SL g2056 ( 
.A(n_2020),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_L g2057 ( 
.A(n_2036),
.B(n_1864),
.Y(n_2057)
);

NAND4xp25_ASAP7_75t_L g2058 ( 
.A(n_2009),
.B(n_1999),
.C(n_1978),
.D(n_2006),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2025),
.B(n_1970),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2028),
.A2(n_1976),
.B1(n_1970),
.B2(n_2006),
.Y(n_2060)
);

AOI21xp33_ASAP7_75t_L g2061 ( 
.A1(n_2049),
.A2(n_2017),
.B(n_2020),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2056),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_L g2063 ( 
.A(n_2050),
.B(n_2026),
.C(n_2019),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2048),
.B(n_2023),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2050),
.A2(n_2033),
.B1(n_2031),
.B2(n_2014),
.C(n_2011),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_2047),
.B(n_2034),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2049),
.A2(n_2057),
.B(n_2054),
.Y(n_2067)
);

OAI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2051),
.A2(n_2058),
.B(n_2041),
.C(n_2044),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2039),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2053),
.B(n_2011),
.Y(n_2070)
);

NAND5xp2_ASAP7_75t_L g2071 ( 
.A(n_2055),
.B(n_2014),
.C(n_2030),
.D(n_1778),
.E(n_1728),
.Y(n_2071)
);

AO22x2_ASAP7_75t_L g2072 ( 
.A1(n_2037),
.A2(n_1970),
.B1(n_1995),
.B2(n_2005),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2059),
.A2(n_1944),
.B1(n_1927),
.B2(n_1887),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2043),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2045),
.B(n_1995),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2040),
.B(n_1884),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_2062),
.B(n_2069),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2070),
.B(n_2046),
.Y(n_2078)
);

NAND3xp33_ASAP7_75t_L g2079 ( 
.A(n_2067),
.B(n_2068),
.C(n_2061),
.Y(n_2079)
);

NAND4xp25_ASAP7_75t_SL g2080 ( 
.A(n_2063),
.B(n_2052),
.C(n_2038),
.D(n_2042),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_2072),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_2074),
.Y(n_2082)
);

AOI322xp5_ASAP7_75t_L g2083 ( 
.A1(n_2064),
.A2(n_2052),
.A3(n_2046),
.B1(n_1865),
.B2(n_1863),
.C1(n_1896),
.C2(n_1898),
.Y(n_2083)
);

HAxp5_ASAP7_75t_SL g2084 ( 
.A(n_2073),
.B(n_2060),
.CON(n_2084),
.SN(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2066),
.B(n_1864),
.Y(n_2085)
);

NAND3xp33_ASAP7_75t_L g2086 ( 
.A(n_2065),
.B(n_1944),
.C(n_1927),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2076),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2075),
.B(n_1904),
.Y(n_2088)
);

NAND2xp33_ASAP7_75t_SL g2089 ( 
.A(n_2072),
.B(n_1771),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_SL g2090 ( 
.A(n_2071),
.B(n_1648),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_2067),
.B(n_1887),
.Y(n_2091)
);

AOI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2079),
.A2(n_1944),
.B1(n_1927),
.B2(n_1895),
.Y(n_2092)
);

XNOR2x1_ASAP7_75t_L g2093 ( 
.A(n_2078),
.B(n_1660),
.Y(n_2093)
);

AOI221x1_ASAP7_75t_L g2094 ( 
.A1(n_2077),
.A2(n_1887),
.B1(n_1895),
.B2(n_1876),
.C(n_1914),
.Y(n_2094)
);

O2A1O1Ixp33_ASAP7_75t_L g2095 ( 
.A1(n_2081),
.A2(n_1746),
.B(n_1927),
.C(n_1944),
.Y(n_2095)
);

AOI211xp5_ASAP7_75t_L g2096 ( 
.A1(n_2080),
.A2(n_2086),
.B(n_2089),
.C(n_2091),
.Y(n_2096)
);

AOI221x1_ASAP7_75t_L g2097 ( 
.A1(n_2077),
.A2(n_1887),
.B1(n_1895),
.B2(n_1911),
.C(n_1876),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2090),
.A2(n_1728),
.B1(n_1660),
.B2(n_1820),
.C(n_1758),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2093),
.B(n_2085),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_2092),
.Y(n_2100)
);

AOI221xp5_ASAP7_75t_SL g2101 ( 
.A1(n_2096),
.A2(n_2082),
.B1(n_2087),
.B2(n_2084),
.C(n_2088),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2098),
.A2(n_2082),
.B1(n_1887),
.B2(n_1895),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2095),
.A2(n_2090),
.B1(n_2083),
.B2(n_1895),
.Y(n_2103)
);

A2O1A1Ixp33_ASAP7_75t_L g2104 ( 
.A1(n_2094),
.A2(n_1903),
.B(n_1820),
.C(n_1753),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_2097),
.A2(n_1746),
.B1(n_1751),
.B2(n_1772),
.C(n_1863),
.Y(n_2105)
);

AOI221x1_ASAP7_75t_L g2106 ( 
.A1(n_2096),
.A2(n_1914),
.B1(n_1876),
.B2(n_1911),
.C(n_1886),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_2099),
.Y(n_2107)
);

INVxp67_ASAP7_75t_L g2108 ( 
.A(n_2100),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2101),
.B(n_1896),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2102),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2106),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2103),
.A2(n_1903),
.B1(n_1727),
.B2(n_1753),
.Y(n_2112)
);

O2A1O1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_2109),
.A2(n_2104),
.B(n_2105),
.C(n_1751),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2107),
.Y(n_2114)
);

NOR2x1p5_ASAP7_75t_L g2115 ( 
.A(n_2107),
.B(n_1676),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_L g2116 ( 
.A(n_2108),
.B(n_1764),
.C(n_1809),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_2114),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2115),
.B(n_2110),
.Y(n_2118)
);

AO22x2_ASAP7_75t_L g2119 ( 
.A1(n_2118),
.A2(n_2111),
.B1(n_2116),
.B2(n_2113),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2119),
.B(n_2117),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2119),
.A2(n_2112),
.B1(n_1901),
.B2(n_1912),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2121),
.B(n_1878),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_2120),
.A2(n_1878),
.B1(n_1912),
.B2(n_1893),
.Y(n_2123)
);

OAI21xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2122),
.A2(n_1676),
.B(n_1764),
.Y(n_2124)
);

XNOR2x1_ASAP7_75t_L g2125 ( 
.A(n_2124),
.B(n_2123),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2125),
.A2(n_1896),
.B1(n_1898),
.B2(n_1893),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_2126),
.Y(n_2127)
);

OAI221xp5_ASAP7_75t_R g2128 ( 
.A1(n_2127),
.A2(n_1782),
.B1(n_1724),
.B2(n_1772),
.C(n_1912),
.Y(n_2128)
);

AOI211xp5_ASAP7_75t_L g2129 ( 
.A1(n_2128),
.A2(n_1626),
.B(n_1628),
.C(n_1715),
.Y(n_2129)
);


endmodule