module fake_jpeg_9188_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_30),
.Y(n_64)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_46),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_27),
.B1(n_36),
.B2(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_42),
.B1(n_17),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_59),
.B1(n_65),
.B2(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_31),
.B(n_33),
.C(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_68),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_34),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_42),
.B1(n_22),
.B2(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_103),
.B1(n_7),
.B2(n_15),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_24),
.B1(n_8),
.B2(n_9),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_74),
.A2(n_98),
.B1(n_100),
.B2(n_80),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_134)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_40),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_87),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_57),
.B1(n_66),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_12),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_12),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_39),
.C(n_45),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_21),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_96),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_23),
.B(n_29),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_83),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_55),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_102),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_45),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_20),
.B1(n_23),
.B2(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_45),
.B1(n_23),
.B2(n_21),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_21),
.B1(n_23),
.B2(n_43),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_77),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_86),
.C(n_73),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_126),
.B1(n_134),
.B2(n_78),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_115),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_69),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_101),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_126)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_131),
.Y(n_149)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_1),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_90),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_104),
.B1(n_106),
.B2(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_72),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_138),
.B(n_153),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_146),
.B1(n_159),
.B2(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_141),
.B(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_154),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_151),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_88),
.B(n_94),
.C(n_93),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_92),
.Y(n_148)
);

NAND2x1p5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_112),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_157),
.C(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_135),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_97),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_69),
.B(n_95),
.C(n_76),
.D(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_108),
.A2(n_110),
.B(n_126),
.C(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_120),
.Y(n_160)
);

NAND4xp25_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_143),
.C(n_163),
.D(n_111),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_85),
.B1(n_80),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_85),
.B1(n_91),
.B2(n_95),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_117),
.B1(n_129),
.B2(n_118),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_85),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_121),
.C(n_107),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_175),
.C(n_151),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_121),
.C(n_116),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_105),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_145),
.B(n_146),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_128),
.A3(n_98),
.B1(n_122),
.B2(n_95),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_105),
.B1(n_91),
.B2(n_130),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_198),
.Y(n_219)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_157),
.B1(n_159),
.B2(n_150),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_194),
.A2(n_196),
.B1(n_197),
.B2(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_164),
.B1(n_140),
.B2(n_144),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_164),
.B1(n_142),
.B2(n_159),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_177),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_139),
.B(n_159),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_186),
.B(n_187),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_174),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_147),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_206),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_210),
.C(n_189),
.Y(n_212)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_224),
.B(n_225),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_223),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_199),
.C(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_186),
.B1(n_179),
.B2(n_182),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_204),
.B(n_198),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_167),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

OAI322xp33_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_171),
.A3(n_165),
.B1(n_172),
.B2(n_170),
.C1(n_168),
.C2(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_1),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_1),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_236),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_197),
.B1(n_196),
.B2(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_209),
.C(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_232),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_209),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_219),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_218),
.B1(n_217),
.B2(n_203),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_221),
.B(n_216),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_244),
.B(n_250),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_201),
.B(n_219),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_217),
.B1(n_212),
.B2(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_201),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_220),
.C(n_226),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_191),
.B1(n_214),
.B2(n_190),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_235),
.B1(n_239),
.B2(n_233),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_254),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_259),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_222),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_247),
.B1(n_245),
.B2(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_260),
.B(n_262),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_233),
.B1(n_240),
.B2(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_222),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_267),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_251),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_264),
.A3(n_261),
.B1(n_240),
.B2(n_253),
.C1(n_229),
.C2(n_228),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_2),
.A3(n_3),
.B1(n_16),
.B2(n_130),
.C1(n_268),
.C2(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_228),
.C(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_227),
.C(n_91),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_274),
.B(n_269),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_130),
.Y(n_276)
);


endmodule