module fake_jpeg_26833_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_0),
.B(n_7),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_76),
.Y(n_89)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_0),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_86),
.Y(n_97)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_65),
.B1(n_58),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_91),
.B1(n_62),
.B2(n_67),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_65),
.B1(n_50),
.B2(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_75),
.B1(n_60),
.B2(n_48),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_105),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_49),
.B1(n_69),
.B2(n_53),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_103),
.B1(n_104),
.B2(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_1),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_106),
.C(n_2),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_61),
.B1(n_57),
.B2(n_51),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_56),
.B1(n_53),
.B2(n_68),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_2),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_68),
.C(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_116),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_96),
.B1(n_95),
.B2(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_122),
.B1(n_9),
.B2(n_10),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_123),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_3),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_99),
.B(n_66),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_6),
.B(n_8),
.Y(n_137)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_23),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_20),
.B(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_18),
.C(n_43),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_17),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_9),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_35),
.B1(n_11),
.B2(n_25),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_142),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_144),
.B1(n_126),
.B2(n_139),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_134),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_145),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_129),
.B(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_128),
.C(n_147),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_28),
.B1(n_30),
.B2(n_37),
.C(n_39),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_41),
.Y(n_157)
);


endmodule