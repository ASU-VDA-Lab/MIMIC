module fake_jpeg_8826_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_16),
.Y(n_52)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_1),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_22),
.C(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_28),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_65),
.B1(n_29),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_30),
.B1(n_18),
.B2(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_30),
.B1(n_18),
.B2(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_30),
.B1(n_20),
.B2(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_26),
.B(n_31),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_16),
.C(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_79),
.B1(n_35),
.B2(n_27),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_76),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_60),
.B1(n_55),
.B2(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_112),
.B1(n_68),
.B2(n_86),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_61),
.C(n_52),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_36),
.B1(n_46),
.B2(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_32),
.B1(n_19),
.B2(n_23),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_23),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_39),
.B(n_41),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_23),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_27),
.B1(n_32),
.B2(n_19),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_46),
.B1(n_39),
.B2(n_19),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_14),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_134),
.B(n_136),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_39),
.B1(n_32),
.B2(n_41),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_51),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_51),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_103),
.B(n_96),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_94),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_153),
.C(n_157),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_104),
.B(n_101),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_157),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_108),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_101),
.B(n_27),
.C(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_132),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_41),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_113),
.C(n_91),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_91),
.C(n_51),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_32),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_129),
.B1(n_124),
.B2(n_126),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_172),
.B1(n_179),
.B2(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_171),
.Y(n_196)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_125),
.C(n_114),
.Y(n_173)
);

AOI31xp67_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_138),
.A3(n_155),
.B(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_116),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_131),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_149),
.B1(n_141),
.B2(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_174),
.B1(n_166),
.B2(n_172),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_156),
.B1(n_158),
.B2(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_2),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_147),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_190),
.C(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_195),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_153),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_98),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_107),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_98),
.Y(n_195)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_194),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_191),
.C(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_167),
.C(n_169),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_177),
.C(n_160),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_171),
.B(n_88),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_208),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_3),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_3),
.B(n_4),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_3),
.Y(n_222)
);

XOR2x2_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_181),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_200),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_107),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_198),
.B(n_5),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_13),
.C(n_10),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_13),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_224),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_204),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_225),
.B(n_228),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_201),
.B(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_203),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_215),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_4),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_6),
.C(n_7),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_217),
.B1(n_220),
.B2(n_7),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_6),
.B(n_7),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_232),
.C(n_231),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_6),
.B(n_8),
.Y(n_243)
);

AOI31xp33_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.A3(n_240),
.B(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_9),
.Y(n_246)
);


endmodule