module real_jpeg_10919_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_317, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_317;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_1),
.A2(n_32),
.B1(n_63),
.B2(n_64),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_3),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_50),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_50),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_4),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_87),
.B1(n_90),
.B2(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_4),
.B(n_102),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_25),
.B(n_27),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_176),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_50),
.B(n_61),
.C(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_69),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_35),
.B1(n_48),
.B2(n_50),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_11),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_13),
.A2(n_48),
.B1(n_50),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_167),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_167),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_14),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_158),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_158),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_158),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_15),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_140),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_140),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_140),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_103),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_83),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_21),
.A2(n_71),
.B1(n_72),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_21),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_22),
.A2(n_23),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_58),
.C(n_70),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_33),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.C(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_24),
.A2(n_29),
.B1(n_37),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_24),
.A2(n_37),
.B1(n_259),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_24),
.A2(n_37),
.B1(n_139),
.B2(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_44),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_27),
.B(n_176),
.CON(n_201),
.SN(n_201)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_28),
.A2(n_31),
.B(n_176),
.C(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_36),
.A2(n_102),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_37),
.A2(n_99),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_37),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_42),
.A2(n_57),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_42),
.A2(n_57),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_42),
.A2(n_112),
.B(n_255),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_47),
.B1(n_52),
.B2(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_43),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_43),
.A2(n_47),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_43),
.A2(n_55),
.B(n_113),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_44),
.B(n_50),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_46),
.A2(n_48),
.B1(n_201),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_75),
.B(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_57),
.B(n_176),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_59),
.B1(n_111),
.B2(n_116),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_67),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_60),
.A2(n_62),
.B1(n_94),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_60),
.A2(n_62),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_60),
.A2(n_62),
.B1(n_166),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_60),
.A2(n_62),
.B1(n_191),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_60),
.A2(n_77),
.B(n_199),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_62),
.B(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_62),
.A2(n_79),
.B(n_136),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_63),
.B(n_66),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_63),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_64),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_68),
.A2(n_82),
.B(n_96),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_97),
.B(n_98),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_85),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_97),
.B1(n_98),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_86),
.A2(n_93),
.B1(n_97),
.B2(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_87),
.A2(n_90),
.B1(n_157),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_87),
.A2(n_134),
.B(n_160),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_87),
.A2(n_91),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_87),
.A2(n_90),
.B1(n_223),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_87),
.A2(n_209),
.B(n_245),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_88),
.A2(n_89),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_92),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_89),
.B(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_90),
.B(n_176),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_90),
.A2(n_132),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_93),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_102),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_117),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_147),
.B(n_315),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_144),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_122),
.B(n_144),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_123),
.B(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_123),
.B(n_307),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.CI(n_129),
.CON(n_123),
.SN(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.C(n_142),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_130),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_131),
.B(n_135),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_143),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_294),
.A3(n_306),
.B1(n_308),
.B2(n_314),
.C(n_317),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_261),
.C(n_290),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_235),
.B(n_260),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_212),
.B(n_234),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_194),
.B(n_211),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_185),
.B(n_193),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_173),
.B(n_184),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_172),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_165),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_179),
.B(n_183),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_195),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.CI(n_192),
.CON(n_188),
.SN(n_188)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_205),
.B2(n_210),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_204),
.C(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_228),
.B2(n_229),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_231),
.C(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_227),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_236),
.B(n_237),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_249),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_248),
.C(n_249),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_253),
.C(n_256),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_277),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_277),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_271),
.C(n_275),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_286),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_286),
.C(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_282),
.C(n_285),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_309),
.B(n_313),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_297),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_303),
.C(n_305),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_309)
);


endmodule