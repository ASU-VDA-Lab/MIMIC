module real_aes_9148_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_0), .A2(n_239), .B(n_240), .C(n_244), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_1), .B(n_180), .Y(n_245) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_3), .B(n_152), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_4), .A2(n_138), .B(n_143), .C(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_5), .A2(n_133), .B(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_6), .A2(n_133), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_7), .B(n_180), .Y(n_546) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_168), .B(n_184), .Y(n_183) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_10), .A2(n_138), .B(n_143), .C(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g484 ( .A(n_11), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_41), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_13), .B(n_243), .Y(n_504) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_15), .B(n_152), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_16), .A2(n_153), .B(n_492), .C(n_494), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_17), .B(n_180), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_18), .A2(n_466), .B1(n_743), .B2(n_749), .C1(n_751), .C2(n_752), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_19), .B(n_217), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_20), .A2(n_143), .B(n_194), .C(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_21), .A2(n_192), .B(n_242), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_22), .B(n_243), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_23), .B(n_243), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_24), .Y(n_531) );
INVx1_ASAP7_75t_L g523 ( .A(n_25), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_26), .A2(n_143), .B(n_187), .C(n_194), .Y(n_186) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_28), .Y(n_500) );
INVx1_ASAP7_75t_L g580 ( .A(n_29), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_30), .A2(n_133), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_32), .A2(n_141), .B(n_156), .C(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_33), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_34), .A2(n_242), .B(n_543), .C(n_545), .Y(n_542) );
INVxp67_ASAP7_75t_L g581 ( .A(n_35), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_36), .A2(n_46), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_37), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_38), .A2(n_143), .B(n_194), .C(n_522), .Y(n_521) );
CKINVDCx14_ASAP7_75t_R g541 ( .A(n_39), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_40), .A2(n_45), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_40), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_42), .A2(n_244), .B(n_482), .C(n_483), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_43), .B(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_44), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_45), .Y(n_747) );
INVx1_ASAP7_75t_L g125 ( .A(n_46), .Y(n_125) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_47), .A2(n_122), .A3(n_456), .B1(n_459), .B2(n_460), .C(n_462), .Y(n_121) );
INVx1_ASAP7_75t_L g459 ( .A(n_47), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_48), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_49), .B(n_133), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_50), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_51), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_52), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
INVx1_ASAP7_75t_L g241 ( .A(n_53), .Y(n_241) );
INVx1_ASAP7_75t_L g147 ( .A(n_54), .Y(n_147) );
INVx1_ASAP7_75t_L g512 ( .A(n_55), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_56), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_57), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_58), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_59), .Y(n_480) );
INVx1_ASAP7_75t_L g139 ( .A(n_60), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_61), .B(n_133), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_62), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_63), .A2(n_174), .B(n_176), .C(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g161 ( .A(n_64), .Y(n_161) );
INVx1_ASAP7_75t_SL g544 ( .A(n_65), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_67), .B(n_152), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_68), .B(n_180), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_104), .B1(n_115), .B2(n_758), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_70), .B(n_153), .Y(n_255) );
INVx1_ASAP7_75t_L g534 ( .A(n_71), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_72), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_73), .B(n_149), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_74), .A2(n_143), .B(n_156), .C(n_226), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_75), .Y(n_172) );
INVx1_ASAP7_75t_L g107 ( .A(n_76), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_77), .A2(n_133), .B(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_78), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_79), .A2(n_133), .B(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_80), .A2(n_211), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g490 ( .A(n_81), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_82), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_83), .B(n_148), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_84), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_84), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_85), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_86), .A2(n_133), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g493 ( .A(n_87), .Y(n_493) );
INVx2_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
INVx1_ASAP7_75t_L g503 ( .A(n_89), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_90), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_91), .B(n_243), .Y(n_256) );
INVx2_ASAP7_75t_L g110 ( .A(n_92), .Y(n_110) );
OR2x2_ASAP7_75t_L g458 ( .A(n_92), .B(n_111), .Y(n_458) );
OR2x2_ASAP7_75t_L g742 ( .A(n_92), .B(n_112), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_93), .A2(n_143), .B(n_156), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_94), .B(n_133), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_95), .Y(n_203) );
INVxp67_ASAP7_75t_L g177 ( .A(n_96), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_97), .B(n_168), .Y(n_485) );
INVx2_ASAP7_75t_L g515 ( .A(n_98), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_99), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g227 ( .A(n_100), .Y(n_227) );
INVx1_ASAP7_75t_L g251 ( .A(n_101), .Y(n_251) );
AND2x2_ASAP7_75t_L g163 ( .A(n_102), .B(n_158), .Y(n_163) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g750 ( .A(n_109), .Y(n_750) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g471 ( .A(n_110), .B(n_112), .Y(n_471) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_464), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g757 ( .A(n_119), .Y(n_757) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_122), .B(n_461), .Y(n_460) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_126), .A2(n_468), .B1(n_472), .B2(n_739), .Y(n_467) );
INVx4_ASAP7_75t_L g755 ( .A(n_126), .Y(n_755) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR5x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_329), .C(n_407), .D(n_431), .E(n_448), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_195), .B(n_246), .C(n_306), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
AND2x2_ASAP7_75t_L g260 ( .A(n_130), .B(n_166), .Y(n_260) );
INVx5_ASAP7_75t_SL g288 ( .A(n_130), .Y(n_288) );
AND2x2_ASAP7_75t_L g324 ( .A(n_130), .B(n_309), .Y(n_324) );
OR2x2_ASAP7_75t_L g363 ( .A(n_130), .B(n_165), .Y(n_363) );
OR2x2_ASAP7_75t_L g394 ( .A(n_130), .B(n_285), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_130), .B(n_298), .Y(n_430) );
AND2x2_ASAP7_75t_L g442 ( .A(n_130), .B(n_285), .Y(n_442) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_158), .Y(n_131) );
BUFx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_134), .B(n_138), .Y(n_252) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_137), .Y(n_243) );
INVx4_ASAP7_75t_SL g157 ( .A(n_138), .Y(n_157) );
BUFx3_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_157), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_142), .A2(n_157), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_142), .A2(n_157), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_142), .A2(n_157), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_142), .A2(n_157), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_142), .A2(n_157), .B(n_541), .C(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_SL g576 ( .A1(n_142), .A2(n_157), .B(n_577), .C(n_578), .Y(n_576) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_148), .A2(n_154), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_L g502 ( .A1(n_148), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_148), .A2(n_505), .B(n_534), .C(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_152), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g239 ( .A(n_152), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_216), .B(n_523), .C(n_524), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_152), .A2(n_175), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_153), .B(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g244 ( .A(n_155), .Y(n_244) );
INVx1_ASAP7_75t_L g494 ( .A(n_155), .Y(n_494) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_158), .A2(n_478), .B(n_485), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_158), .A2(n_252), .B(n_520), .C(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g169 ( .A(n_159), .B(n_160), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g441 ( .A(n_164), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g304 ( .A(n_165), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_166), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
INVx3_ASAP7_75t_L g312 ( .A(n_166), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_166), .B(n_182), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_166), .B(n_288), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_166), .B(n_309), .Y(n_349) );
AND2x2_ASAP7_75t_L g355 ( .A(n_166), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g392 ( .A(n_166), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_166), .B(n_249), .Y(n_406) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_179), .Y(n_166) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_167), .A2(n_488), .B(n_495), .Y(n_487) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_167), .A2(n_510), .B(n_516), .Y(n_509) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_167), .A2(n_539), .B(n_546), .Y(n_538) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g181 ( .A(n_168), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_185), .B(n_186), .Y(n_184) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_175), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_175), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_178), .B(n_579), .Y(n_578) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_235), .B(n_245), .Y(n_234) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_224), .B(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_181), .B(n_233), .Y(n_232) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_181), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_181), .B(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_181), .A2(n_530), .B(n_536), .Y(n_529) );
OR2x2_ASAP7_75t_L g298 ( .A(n_182), .B(n_249), .Y(n_298) );
AND2x2_ASAP7_75t_L g309 ( .A(n_182), .B(n_285), .Y(n_309) );
AND2x2_ASAP7_75t_L g321 ( .A(n_182), .B(n_312), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_182), .B(n_249), .Y(n_344) );
INVx1_ASAP7_75t_SL g356 ( .A(n_182), .Y(n_356) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g248 ( .A(n_183), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_183), .B(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_191), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
AND2x2_ASAP7_75t_L g269 ( .A(n_197), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_197), .B(n_222), .Y(n_273) );
AND2x2_ASAP7_75t_L g276 ( .A(n_197), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g301 ( .A(n_197), .B(n_292), .Y(n_301) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_197), .Y(n_320) );
AND2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g351 ( .A(n_197), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g397 ( .A(n_197), .B(n_280), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_197), .B(n_303), .Y(n_424) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
AND2x2_ASAP7_75t_L g360 ( .A(n_198), .B(n_292), .Y(n_360) );
AND2x2_ASAP7_75t_L g444 ( .A(n_198), .B(n_312), .Y(n_444) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_207), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_207), .Y(n_433) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g263 ( .A(n_208), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g272 ( .A(n_208), .B(n_270), .Y(n_272) );
INVx5_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_234), .Y(n_303) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_212), .B(n_217), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_218), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_221), .A2(n_499), .B(n_506), .Y(n_498) );
INVx1_ASAP7_75t_L g381 ( .A(n_222), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_222), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g414 ( .A(n_222), .B(n_280), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_222), .A2(n_337), .B(n_444), .C(n_445), .Y(n_443) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
BUFx2_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_223), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g545 ( .A(n_230), .Y(n_545) );
INVx2_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_234), .B(n_268), .Y(n_277) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_280), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_242), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g482 ( .A(n_243), .Y(n_482) );
INVx2_ASAP7_75t_L g505 ( .A(n_244), .Y(n_505) );
AOI211x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_261), .B(n_274), .C(n_299), .Y(n_246) );
INVx1_ASAP7_75t_L g365 ( .A(n_247), .Y(n_365) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_260), .Y(n_247) );
INVx5_ASAP7_75t_SL g285 ( .A(n_249), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_249), .B(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g373 ( .A1(n_249), .A2(n_374), .A3(n_376), .B(n_377), .C(n_383), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_249), .A2(n_321), .B(n_409), .C(n_412), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_252), .A2(n_500), .B(n_501), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_252), .A2(n_531), .B(n_532), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g573 ( .A(n_259), .Y(n_573) );
INVxp67_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
NAND4xp25_ASAP7_75t_SL g261 ( .A(n_262), .B(n_265), .C(n_271), .D(n_273), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_262), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g319 ( .A(n_263), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_266), .B(n_272), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_266), .B(n_279), .Y(n_399) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_267), .B(n_280), .Y(n_417) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVxp67_ASAP7_75t_L g327 ( .A(n_269), .Y(n_327) );
AND2x4_ASAP7_75t_L g279 ( .A(n_270), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g353 ( .A(n_270), .B(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g380 ( .A(n_270), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_270), .B(n_367), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_271), .B(n_341), .Y(n_361) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_272), .B(n_294), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_272), .B(n_341), .Y(n_440) );
INVx1_ASAP7_75t_L g451 ( .A(n_273), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B(n_281), .C(n_289), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_277), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g290 ( .A(n_279), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_279), .B(n_341), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_279), .B(n_360), .Y(n_384) );
OR2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g404 ( .A(n_280), .B(n_360), .Y(n_404) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_282), .A2(n_294), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_415) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g305 ( .A(n_285), .B(n_288), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_285), .B(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_285), .B(n_312), .Y(n_420) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g419 ( .A(n_287), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_288), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g386 ( .A(n_288), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_288), .B(n_335), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_288), .B(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_295), .Y(n_289) );
INVx2_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
OR2x2_ASAP7_75t_L g346 ( .A(n_294), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g449 ( .A(n_294), .B(n_417), .Y(n_449) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g453 ( .A(n_300), .Y(n_453) );
INVx2_ASAP7_75t_SL g367 ( .A(n_301), .Y(n_367) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_304), .A2(n_385), .B(n_449), .C(n_450), .Y(n_448) );
OAI322xp33_ASAP7_75t_SL g317 ( .A1(n_305), .A2(n_318), .A3(n_321), .B1(n_322), .B2(n_323), .C1(n_325), .C2(n_328), .Y(n_317) );
INVx2_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_314), .B2(n_316), .C(n_317), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_SL g383 ( .A1(n_308), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_309), .B(n_312), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_309), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g382 ( .A(n_311), .B(n_344), .Y(n_382) );
INVx1_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_316), .A2(n_426), .B(n_428), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp67_ASAP7_75t_SL g379 ( .A(n_320), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_320), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g436 ( .A(n_321), .Y(n_436) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_330), .B(n_357), .C(n_373), .D(n_389), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_338), .C(n_350), .Y(n_330) );
INVx1_ASAP7_75t_L g422 ( .A(n_331), .Y(n_422) );
AND2x2_ASAP7_75t_L g370 ( .A(n_332), .B(n_353), .Y(n_370) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_337), .B(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_346), .B2(n_348), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_340), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_380), .B(n_403), .C(n_405), .Y(n_402) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g447 ( .A(n_345), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g437 ( .A(n_346), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g376 ( .A(n_355), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B(n_362), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_369), .B2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_367), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_372), .B(n_393), .Y(n_455) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_381), .B(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B1(n_398), .B2(n_400), .C(n_402), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_415), .C(n_425), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .C(n_443), .Y(n_431) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_439), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g461 ( .A(n_458), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_461), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_462), .B(n_465), .C(n_756), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI22x1_ASAP7_75t_SL g753 ( .A1(n_468), .A2(n_739), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g754 ( .A(n_472), .Y(n_754) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_669), .Y(n_472) );
NAND5xp2_ASAP7_75t_L g473 ( .A(n_474), .B(n_584), .C(n_616), .D(n_633), .E(n_656), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_517), .B1(n_547), .B2(n_551), .C(n_555), .Y(n_474) );
INVx1_ASAP7_75t_L g696 ( .A(n_475), .Y(n_696) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_496), .Y(n_475) );
AND3x2_ASAP7_75t_L g671 ( .A(n_476), .B(n_498), .C(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_477), .B(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g562 ( .A(n_477), .Y(n_562) );
AND2x2_ASAP7_75t_L g566 ( .A(n_477), .B(n_508), .Y(n_566) );
INVx2_ASAP7_75t_L g593 ( .A(n_477), .Y(n_593) );
OR2x2_ASAP7_75t_L g604 ( .A(n_477), .B(n_509), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_477), .B(n_497), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_477), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g683 ( .A(n_477), .B(n_509), .Y(n_683) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
AND2x2_ASAP7_75t_L g624 ( .A(n_486), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_486), .B(n_497), .Y(n_643) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g554 ( .A(n_487), .B(n_497), .Y(n_554) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
AND2x2_ASAP7_75t_L g610 ( .A(n_487), .B(n_509), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_487), .B(n_496), .C(n_593), .Y(n_635) );
AND2x2_ASAP7_75t_L g700 ( .A(n_487), .B(n_498), .Y(n_700) );
AND2x2_ASAP7_75t_L g734 ( .A(n_487), .B(n_497), .Y(n_734) );
INVxp67_ASAP7_75t_L g563 ( .A(n_496), .Y(n_563) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_497), .B(n_593), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_497), .B(n_624), .Y(n_632) );
AND2x2_ASAP7_75t_L g682 ( .A(n_497), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g710 ( .A(n_497), .Y(n_710) );
INVx4_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g617 ( .A(n_498), .B(n_610), .Y(n_617) );
BUFx3_ASAP7_75t_L g649 ( .A(n_498), .Y(n_649) );
INVx2_ASAP7_75t_L g625 ( .A(n_508), .Y(n_625) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_509), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_517), .A2(n_685), .B1(n_687), .B2(n_688), .Y(n_684) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
AND2x2_ASAP7_75t_L g547 ( .A(n_518), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_SL g558 ( .A(n_518), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_518), .B(n_588), .Y(n_620) );
OR2x2_ASAP7_75t_L g639 ( .A(n_518), .B(n_528), .Y(n_639) );
AND2x2_ASAP7_75t_L g644 ( .A(n_518), .B(n_596), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_518), .B(n_589), .Y(n_647) );
AND2x2_ASAP7_75t_L g659 ( .A(n_518), .B(n_538), .Y(n_659) );
AND2x2_ASAP7_75t_L g675 ( .A(n_518), .B(n_529), .Y(n_675) );
AND2x4_ASAP7_75t_L g678 ( .A(n_518), .B(n_549), .Y(n_678) );
OR2x2_ASAP7_75t_L g695 ( .A(n_518), .B(n_631), .Y(n_695) );
OR2x2_ASAP7_75t_L g726 ( .A(n_518), .B(n_571), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_518), .B(n_654), .Y(n_728) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g602 ( .A(n_527), .B(n_569), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_527), .B(n_589), .Y(n_721) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_538), .Y(n_527) );
AND2x2_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g588 ( .A(n_528), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g596 ( .A(n_528), .B(n_571), .Y(n_596) );
AND2x2_ASAP7_75t_L g614 ( .A(n_528), .B(n_549), .Y(n_614) );
OR2x2_ASAP7_75t_L g631 ( .A(n_528), .B(n_589), .Y(n_631) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g550 ( .A(n_529), .Y(n_550) );
AND2x2_ASAP7_75t_L g654 ( .A(n_529), .B(n_538), .Y(n_654) );
INVx2_ASAP7_75t_L g549 ( .A(n_538), .Y(n_549) );
INVx1_ASAP7_75t_L g666 ( .A(n_538), .Y(n_666) );
AND2x2_ASAP7_75t_L g716 ( .A(n_538), .B(n_558), .Y(n_716) );
AND2x2_ASAP7_75t_L g568 ( .A(n_548), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g600 ( .A(n_548), .B(n_558), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_548), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x2_ASAP7_75t_L g587 ( .A(n_549), .B(n_558), .Y(n_587) );
OR2x2_ASAP7_75t_L g703 ( .A(n_550), .B(n_677), .Y(n_703) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_553), .B(n_683), .Y(n_689) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OAI32xp33_ASAP7_75t_L g645 ( .A1(n_554), .A2(n_646), .A3(n_648), .B1(n_650), .B2(n_651), .Y(n_645) );
OR2x2_ASAP7_75t_L g662 ( .A(n_554), .B(n_604), .Y(n_662) );
OAI21xp33_ASAP7_75t_SL g687 ( .A1(n_554), .A2(n_564), .B(n_592), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B1(n_564), .B2(n_567), .Y(n_555) );
INVxp33_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_557), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_558), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g613 ( .A(n_558), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g713 ( .A(n_558), .B(n_654), .Y(n_713) );
OR2x2_ASAP7_75t_L g737 ( .A(n_558), .B(n_631), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g720 ( .A1(n_559), .A2(n_619), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_561), .B(n_566), .Y(n_615) );
AND2x2_ASAP7_75t_L g637 ( .A(n_562), .B(n_610), .Y(n_637) );
INVx1_ASAP7_75t_L g650 ( .A(n_562), .Y(n_650) );
OR2x2_ASAP7_75t_L g655 ( .A(n_562), .B(n_589), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_565), .B(n_604), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g585 ( .A1(n_566), .A2(n_586), .B1(n_591), .B2(n_595), .Y(n_585) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_569), .A2(n_628), .B1(n_635), .B2(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g712 ( .A(n_569), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_571), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g731 ( .A(n_571), .B(n_614), .Y(n_731) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_582), .Y(n_571) );
INVx1_ASAP7_75t_L g590 ( .A(n_572), .Y(n_590) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_575), .A2(n_583), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_597), .B1(n_598), .B2(n_603), .C(n_605), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_587), .B(n_589), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g606 ( .A(n_588), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_588), .A2(n_694), .B(n_695), .C(n_696), .Y(n_693) );
AND2x2_ASAP7_75t_L g698 ( .A(n_588), .B(n_678), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_SL g736 ( .A1(n_588), .A2(n_677), .B(n_737), .C(n_738), .Y(n_736) );
BUFx3_ASAP7_75t_L g628 ( .A(n_589), .Y(n_628) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_592), .B(n_649), .Y(n_692) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_592), .A2(n_712), .B(n_714), .C(n_720), .Y(n_711) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVxp67_ASAP7_75t_L g672 ( .A(n_594), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_596), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_600), .A2(n_617), .B(n_618), .C(n_626), .Y(n_616) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g701 ( .A(n_604), .Y(n_701) );
OR2x2_ASAP7_75t_L g718 ( .A(n_604), .B(n_648), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_612), .B2(n_615), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_607), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
OR2x2_ASAP7_75t_L g705 ( .A(n_609), .B(n_649), .Y(n_705) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g660 ( .A(n_610), .B(n_650), .Y(n_660) );
INVx1_ASAP7_75t_L g668 ( .A(n_611), .Y(n_668) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_614), .B(n_628), .Y(n_676) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_624), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g733 ( .A(n_625), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_632), .Y(n_626) );
INVx1_ASAP7_75t_L g663 ( .A(n_627), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_628), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_628), .B(n_659), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_628), .B(n_654), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_628), .B(n_675), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_628), .A2(n_638), .B(n_678), .C(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_638), .B1(n_640), .B2(n_644), .C(n_645), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_642), .B(n_650), .Y(n_724) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_644), .A2(n_659), .B(n_661), .C(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_647), .B(n_654), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_648), .B(n_701), .Y(n_738) );
CKINVDCx16_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
INVxp33_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
AOI21xp33_ASAP7_75t_SL g664 ( .A1(n_653), .A2(n_665), .B(n_667), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_653), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_654), .B(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_660), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g694 ( .A(n_666), .Y(n_694) );
NAND5xp2_ASAP7_75t_L g669 ( .A(n_670), .B(n_697), .C(n_711), .D(n_722), .E(n_735), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B(n_680), .C(n_693), .Y(n_670) );
INVx2_ASAP7_75t_SL g717 ( .A(n_671), .Y(n_717) );
NAND4xp25_ASAP7_75t_SL g673 ( .A(n_674), .B(n_676), .C(n_677), .D(n_679), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_679), .A2(n_681), .B(n_684), .C(n_690), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_682), .A2(n_723), .B1(n_725), .B2(n_727), .C(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_699), .B1(n_702), .B2(n_704), .C(n_706), .Y(n_697) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_705), .A2(n_728), .B1(n_730), .B2(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_743), .Y(n_751) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
endmodule