module real_jpeg_25931_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_36),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_0),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_2),
.B(n_43),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_2),
.B(n_40),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_2),
.B(n_50),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_2),
.B(n_387),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_6),
.B(n_43),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_50),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_6),
.B(n_131),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_6),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_7),
.B(n_43),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_7),
.B(n_40),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_50),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_7),
.B(n_327),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_8),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_8),
.B(n_40),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_8),
.B(n_50),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_8),
.B(n_205),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_10),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_10),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_10),
.B(n_43),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_10),
.B(n_36),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_10),
.B(n_40),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_10),
.B(n_50),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_10),
.B(n_131),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_10),
.B(n_327),
.Y(n_363)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_12),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_12),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_36),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_12),
.B(n_40),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_50),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_12),
.B(n_205),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_13),
.B(n_61),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_13),
.B(n_43),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_13),
.B(n_36),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_13),
.B(n_40),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_13),
.B(n_50),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_13),
.B(n_131),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_13),
.B(n_327),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_50),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_14),
.B(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_16),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_16),
.B(n_50),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_16),
.B(n_131),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_16),
.B(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_382),
.B(n_383),
.C(n_388),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_372),
.C(n_381),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_357),
.C(n_358),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_335),
.C(n_336),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_302),
.C(n_303),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_277),
.C(n_278),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_245),
.C(n_246),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_207),
.C(n_208),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_170),
.C(n_171),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_138),
.C(n_139),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_112),
.C(n_113),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_72),
.C(n_84),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_36),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_64),
.C(n_65),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_71),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_83),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_108),
.C(n_109),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.C(n_98),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.C(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.C(n_103),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_107),
.B(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_127),
.C(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_122),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.CI(n_125),
.CON(n_122),
.SN(n_122)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_136),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_154),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.C(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_150),
.C(n_153),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_145),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.CI(n_148),
.CON(n_145),
.SN(n_145)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_147),
.C(n_148),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_162),
.C(n_168),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_162),
.B1(n_168),
.B2(n_169),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_160),
.B(n_161),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_196),
.C(n_197),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_191)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_164),
.Y(n_329)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_164),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_192),
.B2(n_206),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_193),
.C(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_176),
.C(n_185),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_181),
.C(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_179),
.B(n_231),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_190),
.C(n_191),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_189),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_241),
.C(n_242),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_202),
.CI(n_204),
.CON(n_198),
.SN(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_243),
.B2(n_244),
.Y(n_208)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_235),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_235),
.C(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_222),
.C(n_223),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_214),
.B(n_220),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_220),
.B(n_231),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_234),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_229),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_233),
.C(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_252),
.C(n_255),
.Y(n_300)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_249),
.C(n_276),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_263),
.B2(n_276),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_258),
.C(n_259),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_256),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g317 ( 
.A(n_255),
.B(n_282),
.C(n_285),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_259),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.CI(n_262),
.CON(n_259),
.SN(n_259)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_275),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_271),
.C(n_273),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_273),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_299),
.C(n_300),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_301),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_292),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_292),
.C(n_301),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_287),
.C(n_288),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_285),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_SL g346 ( 
.A(n_285),
.B(n_310),
.C(n_312),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_288),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.CI(n_291),
.CON(n_288),
.SN(n_288)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_306),
.C(n_319),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_319),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_316),
.C(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_313),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_351),
.C(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_322),
.C(n_325),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_331),
.C(n_334),
.Y(n_344)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_336)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_339),
.C(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_345),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_346),
.C(n_347),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_359),
.C(n_361),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.CI(n_344),
.CON(n_341),
.SN(n_341)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_348),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_349),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_350),
.A2(n_351),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_368),
.C(n_371),
.Y(n_374)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_364),
.C(n_365),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_368),
.A2(n_369),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_SL g389 ( 
.A(n_369),
.B(n_376),
.C(n_379),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_370),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_375),
.C(n_380),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_378),
.A2(n_379),
.B1(n_386),
.B2(n_388),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_379),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_386),
.Y(n_388)
);


endmodule