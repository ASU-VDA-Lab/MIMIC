module fake_aes_9389_n_645 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_645);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_645;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_36), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_20), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_53), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_1), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_8), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_37), .Y(n_80) );
BUFx2_ASAP7_75t_SL g81 ( .A(n_56), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_28), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_58), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_70), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_5), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_49), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_46), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_69), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_13), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_14), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_21), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_27), .Y(n_94) );
NOR2xp67_ASAP7_75t_L g95 ( .A(n_63), .B(n_40), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_38), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_48), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_4), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_21), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_66), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_59), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_15), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_5), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_23), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_4), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_7), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_61), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_72), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_43), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_102), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_112), .B(n_0), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_113), .B(n_3), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_104), .B(n_3), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_93), .B(n_6), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_120), .B(n_6), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_76), .B(n_7), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_76), .B(n_8), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_98), .B(n_9), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_102), .B(n_78), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_78), .B(n_9), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_82), .B(n_10), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_85), .B(n_10), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_100), .B(n_11), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_79), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_85), .B(n_12), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_83), .B(n_12), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_88), .B(n_16), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
XNOR2xp5_ASAP7_75t_L g156 ( .A(n_107), .B(n_16), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
AND3x1_ASAP7_75t_L g160 ( .A(n_90), .B(n_17), .C(n_18), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_160), .A2(n_103), .B1(n_89), .B2(n_109), .Y(n_161) );
OAI221xp5_ASAP7_75t_L g162 ( .A1(n_152), .A2(n_91), .B1(n_118), .B2(n_90), .C(n_116), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_121), .B(n_118), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_139), .B(n_119), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_139), .B(n_91), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_139), .B(n_92), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_139), .B(n_92), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_121), .B(n_94), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_157), .B(n_105), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_157), .B(n_110), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_142), .B(n_105), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_158), .B(n_117), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_127), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_146), .B(n_116), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_111), .B1(n_114), .B2(n_117), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_147), .B(n_111), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_128), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_122), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_124), .B(n_114), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_128), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_122), .B(n_81), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_124), .B(n_106), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_129), .B(n_86), .Y(n_200) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_129), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_130), .B(n_106), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_130), .B(n_81), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_128), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_131), .B(n_159), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_131), .B(n_97), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
AND3x4_ASAP7_75t_L g210 ( .A(n_156), .B(n_95), .C(n_18), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_132), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_132), .B(n_97), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_136), .B(n_96), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_123), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_205), .Y(n_217) );
INVx5_ASAP7_75t_L g218 ( .A(n_163), .Y(n_218) );
AND3x1_ASAP7_75t_L g219 ( .A(n_161), .B(n_125), .C(n_126), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_203), .B(n_159), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_192), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_192), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_184), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_205), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_205), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_175), .B(n_155), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_182), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_182), .Y(n_228) );
OR2x4_ASAP7_75t_L g229 ( .A(n_183), .B(n_133), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
AND3x1_ASAP7_75t_SL g231 ( .A(n_162), .B(n_126), .C(n_156), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_203), .B(n_155), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_163), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_201), .B(n_150), .Y(n_234) );
BUFx12f_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_211), .B(n_153), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_201), .A2(n_136), .B(n_137), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_186), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_197), .B(n_140), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_163), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_197), .A2(n_153), .B1(n_137), .B2(n_141), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_182), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_211), .B(n_140), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_163), .B(n_151), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_173), .B(n_151), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_182), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_182), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_168), .B(n_135), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_186), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_214), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_214), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_168), .B(n_135), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_190), .B(n_165), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_161), .Y(n_255) );
INVx5_ASAP7_75t_L g256 ( .A(n_187), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_182), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_174), .B(n_134), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_200), .B(n_134), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_208), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_168), .B(n_144), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_208), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_174), .A2(n_138), .B1(n_149), .B2(n_20), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_168), .B(n_149), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_208), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_201), .Y(n_269) );
NOR2x1p5_ASAP7_75t_L g270 ( .A(n_190), .B(n_149), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_201), .B(n_42), .Y(n_271) );
BUFx4f_ASAP7_75t_L g272 ( .A(n_180), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_169), .B(n_17), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_189), .A2(n_19), .B1(n_22), .B2(n_24), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_164), .Y(n_275) );
BUFx8_ASAP7_75t_L g276 ( .A(n_221), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_224), .A2(n_196), .B1(n_177), .B2(n_198), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_239), .A2(n_187), .B1(n_196), .B2(n_188), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_239), .B(n_165), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_238), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_217), .Y(n_282) );
INVx8_ASAP7_75t_L g283 ( .A(n_235), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_239), .B(n_213), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_238), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g286 ( .A1(n_224), .A2(n_196), .B(n_213), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_249), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_221), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_235), .B(n_169), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_248), .B(n_213), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_275), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_249), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_225), .B(n_187), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_227), .A2(n_164), .B(n_198), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_225), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_256), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_222), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_230), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_248), .B(n_213), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_248), .B(n_206), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_258), .A2(n_215), .B(n_166), .C(n_212), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_250), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_251), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_251), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_226), .B(n_189), .C(n_194), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_223), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_252), .A2(n_210), .B1(n_180), .B2(n_188), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_272), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_264), .Y(n_315) );
NOR2x1_ASAP7_75t_R g316 ( .A(n_255), .B(n_210), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_264), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_256), .B(n_164), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_233), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_258), .B(n_206), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_244), .B(n_169), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_320), .B(n_252), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_309), .A2(n_273), .B(n_274), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_276), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_312), .A2(n_252), .B1(n_210), .B2(n_270), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_279), .B(n_229), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_320), .A2(n_270), .B1(n_263), .B2(n_267), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_276), .A2(n_255), .B1(n_253), .B2(n_219), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_288), .B(n_220), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_303), .A2(n_263), .B1(n_267), .B2(n_180), .Y(n_332) );
AO21x1_ASAP7_75t_L g333 ( .A1(n_281), .A2(n_271), .B(n_179), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_313), .A2(n_263), .B1(n_267), .B2(n_188), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_285), .B(n_253), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_313), .B(n_232), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_285), .A2(n_244), .B1(n_206), .B2(n_272), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_299), .B(n_229), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_296), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_287), .A2(n_188), .B1(n_169), .B2(n_170), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_296), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_237), .B(n_247), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_287), .A2(n_244), .B1(n_206), .B2(n_272), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_293), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_293), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_291), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_276), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_305), .A2(n_170), .B1(n_241), .B2(n_164), .Y(n_350) );
AOI21x1_ASAP7_75t_SL g351 ( .A1(n_321), .A2(n_202), .B(n_236), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_326), .Y(n_352) );
NAND2x1_ASAP7_75t_L g353 ( .A(n_325), .B(n_306), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_328), .A2(n_304), .B1(n_298), .B2(n_300), .C(n_245), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
BUFx2_ASAP7_75t_SL g356 ( .A(n_325), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_330), .B(n_298), .C(n_266), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_330), .A2(n_321), .B1(n_289), .B2(n_311), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g359 ( .A1(n_327), .A2(n_259), .B(n_283), .C(n_199), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_349), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_337), .A2(n_283), .B1(n_321), .B2(n_316), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_328), .A2(n_338), .B1(n_327), .B2(n_324), .C(n_335), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_331), .B(n_284), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_170), .B1(n_290), .B2(n_302), .C(n_301), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_342), .A2(n_286), .B(n_306), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_336), .B(n_308), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_324), .A2(n_321), .B1(n_289), .B2(n_283), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_331), .B(n_283), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_329), .A2(n_283), .B(n_286), .C(n_278), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_289), .B1(n_244), .B2(n_317), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_331), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_347), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_346), .B(n_308), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_329), .A2(n_243), .B(n_282), .C(n_234), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_373), .B(n_347), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_357), .A2(n_344), .B1(n_336), .B2(n_323), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_372), .B(n_229), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_358), .A2(n_350), .B1(n_335), .B2(n_289), .C(n_332), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_377), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_377), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_344), .B1(n_336), .B2(n_323), .Y(n_388) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_322), .B1(n_345), .B2(n_348), .C1(n_347), .C2(n_350), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_371), .A2(n_332), .B1(n_334), .B2(n_340), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_359), .A2(n_323), .B1(n_334), .B2(n_348), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_355), .B(n_347), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_363), .B1(n_375), .B2(n_353), .Y(n_393) );
OAI31xp33_ASAP7_75t_L g394 ( .A1(n_370), .A2(n_340), .A3(n_345), .B(n_322), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_375), .A2(n_317), .B1(n_310), .B2(n_315), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_368), .Y(n_396) );
AOI33xp33_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_170), .A3(n_231), .B1(n_191), .B2(n_185), .B3(n_204), .Y(n_397) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_367), .A2(n_204), .B(n_181), .C(n_185), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_315), .B1(n_310), .B2(n_296), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_356), .A2(n_296), .B1(n_280), .B2(n_291), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_365), .B(n_296), .C(n_339), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_356), .A2(n_314), .B1(n_339), .B2(n_280), .Y(n_403) );
AOI33xp33_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_195), .A3(n_181), .B1(n_191), .B2(n_209), .B3(n_179), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_352), .B(n_314), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_318), .B1(n_294), .B2(n_277), .C(n_319), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_353), .A2(n_342), .B1(n_341), .B2(n_339), .C1(n_351), .C2(n_318), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_352), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_360), .B(n_339), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_401), .Y(n_411) );
INVx3_ASAP7_75t_SL g412 ( .A(n_409), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_394), .A2(n_360), .B1(n_297), .B2(n_198), .C(n_177), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_394), .A2(n_342), .B(n_341), .C(n_339), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_383), .B(n_195), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_380), .B(n_208), .C(n_171), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_409), .B(n_280), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_395), .A2(n_341), .B(n_333), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_409), .B(n_280), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_177), .B1(n_198), .B2(n_208), .C(n_209), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_382), .A2(n_280), .B1(n_333), .B2(n_292), .Y(n_424) );
OAI31xp33_ASAP7_75t_L g425 ( .A1(n_389), .A2(n_294), .A3(n_318), .B(n_177), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_386), .B(n_207), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_392), .B(n_207), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_397), .B(n_171), .C(n_207), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_396), .Y(n_432) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_378), .B(n_351), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_379), .B(n_167), .C(n_172), .D(n_176), .Y(n_434) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_393), .A2(n_294), .A3(n_307), .B(n_297), .Y(n_435) );
OAI33xp33_ASAP7_75t_L g436 ( .A1(n_395), .A2(n_167), .A3(n_172), .B1(n_176), .B2(n_178), .B3(n_19), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_409), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_396), .B(n_343), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_381), .B(n_171), .C(n_207), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_384), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_384), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_385), .B(n_22), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_385), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_402), .B(n_343), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_388), .B(n_207), .Y(n_447) );
OAI221xp5_ASAP7_75t_SL g448 ( .A1(n_391), .A2(n_319), .B1(n_292), .B2(n_297), .C(n_307), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_391), .B(n_207), .Y(n_449) );
AND3x1_ASAP7_75t_L g450 ( .A(n_406), .B(n_178), .C(n_26), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_410), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_399), .A2(n_218), .B(n_256), .C(n_171), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_408), .A2(n_240), .A3(n_233), .B(n_262), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_409), .A2(n_333), .B1(n_171), .B2(n_233), .C(n_240), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_343), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_407), .A2(n_398), .B1(n_403), .B2(n_218), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_441), .B(n_404), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_429), .B(n_171), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_453), .A2(n_269), .B(n_218), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_439), .B(n_25), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_431), .B(n_29), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_431), .B(n_30), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
OR2x6_ASAP7_75t_L g468 ( .A(n_443), .B(n_268), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_452), .A2(n_268), .B1(n_246), .B2(n_260), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_439), .B(n_31), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_443), .B(n_33), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_448), .A2(n_269), .B(n_257), .C(n_265), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_455), .B(n_34), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_437), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_426), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_439), .B(n_426), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_432), .B(n_35), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_39), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_455), .B(n_41), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_44), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_437), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_416), .B(n_45), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_442), .B(n_47), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_415), .B(n_51), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_438), .B(n_54), .Y(n_488) );
OAI21xp33_ASAP7_75t_SL g489 ( .A1(n_435), .A2(n_55), .B(n_57), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_438), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_452), .B(n_60), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g494 ( .A1(n_444), .A2(n_242), .A3(n_265), .B1(n_261), .B2(n_257), .B3(n_247), .Y(n_494) );
AOI221x1_ASAP7_75t_L g495 ( .A1(n_418), .A2(n_268), .B1(n_260), .B2(n_246), .C(n_228), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_424), .B(n_262), .C(n_240), .D(n_261), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_452), .B(n_62), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_444), .B(n_64), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_446), .B(n_67), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_433), .B(n_68), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_457), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_412), .B(n_71), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_433), .B(n_74), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_457), .B(n_246), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_412), .B(n_227), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_428), .B(n_228), .Y(n_508) );
NAND3xp33_ASAP7_75t_SL g509 ( .A(n_425), .B(n_242), .C(n_218), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_421), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_428), .B(n_414), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_420), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_414), .B(n_246), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_469), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_478), .B(n_447), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_486), .B(n_447), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
AOI22x1_ASAP7_75t_L g519 ( .A1(n_505), .A2(n_450), .B1(n_436), .B2(n_420), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_478), .B(n_456), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_476), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_486), .B(n_417), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_477), .B(n_449), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_509), .A2(n_440), .B(n_422), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_491), .B(n_427), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_477), .B(n_423), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_459), .B(n_458), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_492), .B(n_434), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_491), .B(n_413), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_489), .B(n_430), .C(n_262), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_475), .B(n_246), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_493), .B(n_260), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_493), .B(n_260), .Y(n_533) );
INVx3_ASAP7_75t_SL g534 ( .A(n_475), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_490), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_483), .B(n_260), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_503), .B(n_454), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_500), .B(n_268), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_483), .Y(n_540) );
AOI21xp33_ASAP7_75t_L g541 ( .A1(n_502), .A2(n_268), .B(n_218), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_503), .B(n_256), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_500), .B(n_256), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_465), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_463), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_463), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_466), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_466), .Y(n_548) );
AOI21xp33_ASAP7_75t_SL g549 ( .A1(n_464), .A2(n_505), .B(n_499), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g550 ( .A1(n_511), .A2(n_510), .B1(n_501), .B2(n_462), .C1(n_471), .C2(n_485), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_464), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_511), .B(n_497), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_467), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_497), .B(n_510), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_462), .B(n_471), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_472), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_506), .B(n_501), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_512), .B(n_499), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_468), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_468), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_479), .B(n_485), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_515), .B(n_479), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_525), .B(n_468), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_552), .B(n_506), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_552), .B(n_513), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_515), .B(n_460), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_554), .B(n_513), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_525), .B(n_482), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_534), .B(n_482), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_468), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_534), .B(n_480), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_527), .B(n_473), .C(n_496), .D(n_504), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_540), .B(n_494), .Y(n_576) );
AND3x1_ASAP7_75t_L g577 ( .A(n_558), .B(n_498), .C(n_487), .Y(n_577) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_519), .B(n_492), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_521), .Y(n_579) );
NAND5xp2_ASAP7_75t_SL g580 ( .A(n_550), .B(n_498), .C(n_470), .D(n_488), .E(n_487), .Y(n_580) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_524), .B(n_480), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_530), .A2(n_472), .B(n_507), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_554), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_520), .B(n_488), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_538), .Y(n_586) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_546), .A2(n_474), .B(n_481), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_544), .Y(n_588) );
AOI211xp5_ASAP7_75t_SL g589 ( .A1(n_551), .A2(n_507), .B(n_508), .C(n_484), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_520), .B(n_495), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_547), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_549), .A2(n_461), .B(n_495), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_545), .B(n_523), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_529), .A2(n_522), .B(n_526), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_559), .Y(n_595) );
NAND4xp75_ASAP7_75t_L g596 ( .A(n_537), .B(n_557), .C(n_555), .D(n_559), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_548), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_537), .B(n_553), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_528), .A2(n_519), .B1(n_556), .B2(n_560), .C(n_561), .Y(n_599) );
AND3x1_ASAP7_75t_L g600 ( .A(n_557), .B(n_560), .C(n_528), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_553), .B(n_543), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_543), .B(n_541), .C(n_536), .Y(n_602) );
OAI21x1_ASAP7_75t_SL g603 ( .A1(n_528), .A2(n_539), .B(n_542), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_542), .Y(n_604) );
XNOR2xp5_ASAP7_75t_L g605 ( .A(n_532), .B(n_533), .Y(n_605) );
XOR2xp5_ASAP7_75t_L g606 ( .A(n_533), .B(n_532), .Y(n_606) );
NAND4xp25_ASAP7_75t_SL g607 ( .A(n_531), .B(n_550), .C(n_549), .D(n_489), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_532), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_533), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_552), .B(n_554), .Y(n_610) );
NAND2xp33_ASAP7_75t_SL g611 ( .A(n_534), .B(n_551), .Y(n_611) );
XNOR2x1_ASAP7_75t_L g612 ( .A(n_528), .B(n_219), .Y(n_612) );
NAND4xp75_ASAP7_75t_L g613 ( .A(n_600), .B(n_581), .C(n_576), .D(n_577), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_607), .A2(n_611), .B(n_599), .Y(n_614) );
AO22x2_ASAP7_75t_L g615 ( .A1(n_612), .A2(n_603), .B1(n_596), .B2(n_595), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_598), .Y(n_616) );
NAND3x1_ASAP7_75t_SL g617 ( .A(n_582), .B(n_611), .C(n_580), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_584), .B(n_593), .Y(n_618) );
OAI211xp5_ASAP7_75t_SL g619 ( .A1(n_594), .A2(n_589), .B(n_590), .C(n_576), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_612), .A2(n_578), .B1(n_574), .B2(n_592), .C(n_570), .Y(n_620) );
NOR4xp75_ASAP7_75t_L g621 ( .A(n_573), .B(n_585), .C(n_587), .D(n_566), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_578), .A2(n_584), .B1(n_563), .B2(n_571), .Y(n_622) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_602), .B(n_584), .Y(n_623) );
XNOR2xp5_ASAP7_75t_L g624 ( .A(n_606), .B(n_605), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_569), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_620), .A2(n_578), .B(n_580), .C(n_595), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_614), .A2(n_568), .B(n_579), .C(n_575), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_616), .B(n_565), .Y(n_628) );
AOI211xp5_ASAP7_75t_SL g629 ( .A1(n_619), .A2(n_563), .B(n_571), .C(n_609), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_615), .A2(n_565), .B1(n_567), .B2(n_608), .Y(n_630) );
OAI221xp5_ASAP7_75t_SL g631 ( .A1(n_622), .A2(n_605), .B1(n_562), .B2(n_567), .C(n_604), .Y(n_631) );
NOR3x1_ASAP7_75t_L g632 ( .A(n_613), .B(n_601), .C(n_583), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_626), .B(n_617), .C(n_623), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_630), .A2(n_615), .B1(n_624), .B2(n_618), .Y(n_634) );
OA22x2_ASAP7_75t_L g635 ( .A1(n_632), .A2(n_621), .B1(n_625), .B2(n_610), .Y(n_635) );
AO22x2_ASAP7_75t_L g636 ( .A1(n_629), .A2(n_586), .B1(n_572), .B2(n_610), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_636), .Y(n_637) );
AOI31xp33_ASAP7_75t_L g638 ( .A1(n_634), .A2(n_627), .A3(n_628), .B(n_631), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_635), .B(n_564), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_639), .B(n_633), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_637), .A2(n_588), .B1(n_597), .B2(n_591), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_641), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_642), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_643), .Y(n_644) );
NAND3x2_ASAP7_75t_L g645 ( .A(n_644), .B(n_640), .C(n_638), .Y(n_645) );
endmodule