module fake_netlist_6_488_n_1802 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1802);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1802;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_82),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_33),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_44),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_40),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_90),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_21),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_107),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_35),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g201 ( 
.A(n_2),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_121),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_94),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_105),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_55),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_103),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_73),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_34),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_101),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_46),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_60),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_65),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_66),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

BUFx2_ASAP7_75t_SL g233 ( 
.A(n_35),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_29),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_53),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_70),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_165),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_119),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_52),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_64),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_11),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_112),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_4),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_160),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_151),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_125),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_62),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_142),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_123),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_59),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_115),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_117),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_122),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_16),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_99),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_88),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_133),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_36),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_75),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_162),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_53),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_126),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_72),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_51),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_39),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_19),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_51),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_50),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_16),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_109),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_71),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_18),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_50),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_159),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_30),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_45),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_14),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_25),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_26),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_139),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_95),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_78),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_34),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_13),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_45),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_118),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_22),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_52),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_22),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_98),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_9),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_49),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_110),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_136),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_87),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_124),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_42),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_214),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_203),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_205),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_206),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_170),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_208),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_210),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_308),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_226),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_232),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_216),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_264),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_215),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_279),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_204),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_204),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_173),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_217),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_265),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_234),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_225),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_168),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_237),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_238),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_181),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_177),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_240),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_241),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_262),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_190),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_219),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_228),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_235),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_244),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_295),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_243),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_292),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_293),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_294),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_245),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_252),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_173),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_286),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_239),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_169),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_169),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_291),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_257),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_291),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_171),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_258),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_260),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_183),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_334),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_352),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_359),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_353),
.B(n_175),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_218),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_406),
.A2(n_187),
.B(n_172),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_335),
.B(n_248),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_336),
.B(n_224),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_354),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_357),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_337),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_342),
.A2(n_275),
.B1(n_333),
.B2(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_196),
.B(n_192),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_248),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_383),
.B(n_175),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_266),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_348),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_361),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_372),
.B(n_266),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_345),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_414),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_347),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_341),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_343),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_368),
.B(n_313),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_343),
.B(n_239),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_371),
.B(n_313),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_346),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_373),
.B(n_198),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_351),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_376),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_344),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_351),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_378),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_362),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_382),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_391),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_396),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_362),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_SL g488 ( 
.A(n_402),
.B(n_176),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_486),
.B(n_399),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_422),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_438),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_441),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_486),
.B(n_410),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_424),
.B(n_402),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_239),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_451),
.B(n_366),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_451),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_435),
.B(n_413),
.Y(n_504)
);

CKINVDCx11_ASAP7_75t_R g505 ( 
.A(n_416),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_455),
.A2(n_355),
.B1(n_390),
.B2(n_349),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_198),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_434),
.B(n_377),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_467),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_456),
.B(n_379),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_202),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_425),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_473),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_488),
.A2(n_324),
.B1(n_287),
.B2(n_278),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_202),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_464),
.B(n_247),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_441),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_239),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_452),
.A2(n_212),
.B(n_207),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_R g532 ( 
.A(n_477),
.B(n_167),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

BUFx6f_ASAP7_75t_SL g537 ( 
.A(n_456),
.Y(n_537)
);

AOI21x1_ASAP7_75t_L g538 ( 
.A1(n_461),
.A2(n_411),
.B(n_222),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_456),
.B(n_175),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

CKINVDCx11_ASAP7_75t_R g543 ( 
.A(n_436),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_477),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_417),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_456),
.B(n_191),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

BUFx6f_ASAP7_75t_SL g551 ( 
.A(n_460),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_454),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_441),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_483),
.B(n_253),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_454),
.B(n_364),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_429),
.B(n_247),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_417),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_431),
.B(n_395),
.C(n_394),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_418),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_459),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_431),
.B(n_398),
.C(n_397),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_449),
.B(n_263),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_460),
.B(n_191),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_167),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_420),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_446),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_449),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_460),
.B(n_403),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_442),
.A2(n_193),
.B1(n_221),
.B2(n_272),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_440),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_446),
.A2(n_233),
.B1(n_401),
.B2(n_400),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_420),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_421),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_430),
.B(n_447),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_421),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_432),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_432),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_446),
.B(n_213),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_433),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_459),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_459),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_458),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_446),
.B(n_178),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_465),
.B(n_268),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_453),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_364),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_465),
.B(n_277),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_418),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_450),
.B(n_404),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_465),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_469),
.B(n_283),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_478),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_418),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_478),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_469),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_469),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_450),
.B(n_404),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_484),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_450),
.A2(n_431),
.B1(n_444),
.B2(n_485),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_418),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_469),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_474),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_481),
.B(n_174),
.C(n_209),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_474),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_475),
.A2(n_270),
.B1(n_230),
.B2(n_298),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_418),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_418),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_485),
.B(n_178),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_480),
.B(n_179),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_423),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_482),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_423),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_481),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_580),
.B(n_176),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_495),
.B(n_431),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_495),
.B(n_444),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_502),
.B(n_444),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_493),
.B(n_439),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_592),
.B(n_375),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_502),
.B(n_444),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_597),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_509),
.A2(n_290),
.B1(n_186),
.B2(n_323),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_508),
.B(n_474),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_552),
.A2(n_305),
.B1(n_184),
.B2(n_182),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_490),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_597),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_552),
.B(n_179),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_569),
.A2(n_375),
.B(n_387),
.C(n_380),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_544),
.B(n_380),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_503),
.B(n_180),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_474),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_556),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_556),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_637),
.B(n_180),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_510),
.B(n_474),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_510),
.B(n_489),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_573),
.B(n_182),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_507),
.A2(n_296),
.B1(n_271),
.B2(n_269),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_577),
.B(n_184),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_511),
.B(n_489),
.Y(n_672)
);

INVxp33_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_625),
.B(n_523),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_520),
.A2(n_304),
.B1(n_197),
.B2(n_189),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_625),
.B(n_185),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_598),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_587),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_572),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_544),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_625),
.B(n_185),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_489),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_514),
.B(n_489),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_628),
.B(n_632),
.C(n_499),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_525),
.A2(n_303),
.B1(n_261),
.B2(n_259),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_504),
.B(n_186),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_554),
.B(n_491),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_584),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_584),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_555),
.B(n_223),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_532),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_514),
.B(n_489),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_496),
.B(n_188),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_594),
.A2(n_423),
.B(n_427),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_572),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_588),
.B(n_188),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_517),
.B(n_489),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_519),
.B(n_463),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_519),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_601),
.A2(n_328),
.B(n_227),
.C(n_229),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_522),
.B(n_463),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_506),
.B(n_194),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_512),
.B(n_194),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_587),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_522),
.B(n_463),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_606),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_609),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_550),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_540),
.B(n_201),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_618),
.B(n_463),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_555),
.B(n_463),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_503),
.B(n_195),
.Y(n_720)
);

INVx8_ASAP7_75t_L g721 ( 
.A(n_537),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_557),
.B(n_463),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_546),
.B(n_195),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_550),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_609),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_557),
.B(n_231),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_568),
.B(n_423),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_568),
.B(n_423),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_524),
.B(n_423),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_598),
.B(n_384),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_613),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_587),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_537),
.A2(n_329),
.B1(n_200),
.B2(n_305),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_566),
.B(n_199),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_593),
.B(n_200),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_624),
.B(n_314),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_524),
.B(n_427),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_537),
.A2(n_332),
.B1(n_314),
.B2(n_318),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_501),
.B(n_318),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_526),
.B(n_427),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_613),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_565),
.B(n_427),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_614),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_561),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_612),
.B(n_631),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_505),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_526),
.B(n_427),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_545),
.B(n_559),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_574),
.B(n_323),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_560),
.B(n_564),
.Y(n_752)
);

INVx6_ASAP7_75t_L g753 ( 
.A(n_587),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_529),
.B(n_427),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_614),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_529),
.B(n_439),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_327),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_545),
.B(n_251),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_559),
.B(n_274),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_615),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_562),
.B(n_567),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_515),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_520),
.B(n_384),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_560),
.B(n_327),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_537),
.B(n_329),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_562),
.Y(n_766)
);

INVx8_ASAP7_75t_L g767 ( 
.A(n_551),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_567),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_561),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_564),
.B(n_332),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_551),
.B(n_599),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_551),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_615),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_570),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_551),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_534),
.B(n_443),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_543),
.B(n_386),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_578),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_616),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_635),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_534),
.B(n_443),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_535),
.B(n_487),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_588),
.B(n_605),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_535),
.A2(n_276),
.B(n_281),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_588),
.B(n_312),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_211),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_588),
.A2(n_319),
.B1(n_487),
.B2(n_309),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_547),
.B(n_386),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_588),
.B(n_181),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_578),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_585),
.Y(n_791)
);

INVxp33_ASAP7_75t_L g792 ( 
.A(n_558),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_588),
.A2(n_307),
.B1(n_197),
.B2(n_302),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_547),
.B(n_242),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_585),
.B(n_387),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_616),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_539),
.B(n_388),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_586),
.B(n_230),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_530),
.B(n_388),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_589),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_539),
.B(n_389),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_617),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_790),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_778),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_669),
.B(n_675),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_647),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_778),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_686),
.B(n_589),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_677),
.B(n_590),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_766),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_697),
.B(n_591),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_673),
.Y(n_812)
);

HB1xp67_ASAP7_75t_SL g813 ( 
.A(n_748),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_764),
.A2(n_770),
.B(n_664),
.C(n_663),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_647),
.Y(n_815)
);

CKINVDCx8_ASAP7_75t_R g816 ( 
.A(n_681),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_768),
.Y(n_817)
);

BUFx8_ASAP7_75t_L g818 ( 
.A(n_682),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_752),
.B(n_547),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_774),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_660),
.B(n_798),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_678),
.B(n_591),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_648),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_648),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_SL g825 ( 
.A(n_679),
.B(n_302),
.C(n_189),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_752),
.A2(n_531),
.B1(n_617),
.B2(n_619),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_743),
.A2(n_603),
.B(n_608),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_651),
.A2(n_602),
.B1(n_604),
.B2(n_610),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_791),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_800),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_792),
.B(n_602),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_657),
.B(n_230),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_647),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_731),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_641),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_638),
.B(n_604),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_747),
.A2(n_610),
.B1(n_621),
.B2(n_622),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_780),
.B(n_298),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_643),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_751),
.A2(n_541),
.B(n_401),
.C(n_393),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_646),
.B(n_389),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_683),
.B(n_553),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_683),
.B(n_553),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_392),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_746),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_679),
.B(n_393),
.C(n_392),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_648),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_695),
.B(n_703),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_730),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_650),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_707),
.B(n_400),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_762),
.B(n_621),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_750),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_730),
.B(n_298),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_690),
.A2(n_531),
.B1(n_619),
.B2(n_626),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_730),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_674),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_676),
.A2(n_622),
.B1(n_611),
.B2(n_608),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_744),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_763),
.B(n_365),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_R g862 ( 
.A(n_721),
.B(n_304),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_642),
.A2(n_531),
.B1(n_626),
.B2(n_541),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_683),
.B(n_553),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_693),
.A2(n_710),
.B1(n_740),
.B2(n_733),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_661),
.B(n_494),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_761),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_681),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_718),
.A2(n_563),
.B(n_583),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_782),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_782),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_702),
.B(n_718),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_658),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_702),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_684),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_702),
.B(n_789),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_746),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_716),
.B(n_563),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_769),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_724),
.B(n_494),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_786),
.B(n_494),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_681),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_769),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_756),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_769),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_642),
.A2(n_516),
.B1(n_518),
.B2(n_521),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_685),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_SL g888 ( 
.A(n_639),
.B(n_310),
.C(n_307),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_720),
.B(n_513),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_682),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_736),
.B(n_513),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_756),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_776),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_668),
.B(n_513),
.Y(n_894)
);

BUFx12f_ASAP7_75t_L g895 ( 
.A(n_777),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_784),
.A2(n_518),
.B(n_516),
.C(n_492),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_712),
.B(n_563),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_644),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_644),
.A2(n_498),
.B1(n_497),
.B2(n_521),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_781),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_706),
.B(n_527),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_709),
.B(n_527),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_665),
.B(n_365),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_735),
.A2(n_320),
.B(n_309),
.C(n_310),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_645),
.A2(n_498),
.B1(n_497),
.B2(n_492),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_654),
.B(n_527),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_645),
.A2(n_331),
.B(n_330),
.C(n_326),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_640),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_783),
.A2(n_603),
.B(n_611),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_652),
.B(n_527),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_R g911 ( 
.A(n_721),
.B(n_316),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_781),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_713),
.B(n_528),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_655),
.B(n_528),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_753),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_795),
.B(n_608),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_797),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_721),
.B(n_561),
.Y(n_918)
);

NOR2x1p5_ASAP7_75t_L g919 ( 
.A(n_797),
.B(n_316),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_777),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_680),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_649),
.A2(n_575),
.B(n_528),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_767),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_654),
.B(n_528),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_777),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_793),
.A2(n_331),
.B(n_326),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_649),
.A2(n_603),
.B(n_611),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_753),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_662),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_784),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_753),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_788),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_687),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_692),
.B(n_575),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_794),
.A2(n_596),
.B1(n_583),
.B2(n_581),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_723),
.B(n_575),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_662),
.B(n_575),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_788),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_688),
.B(n_581),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_SL g940 ( 
.A(n_737),
.B(n_322),
.C(n_321),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_788),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_717),
.B(n_367),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_767),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_671),
.B(n_246),
.C(n_249),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_688),
.B(n_689),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_653),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_767),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_700),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_801),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_711),
.B(n_581),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_689),
.B(n_581),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_765),
.A2(n_771),
.B1(n_757),
.B2(n_704),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_SL g953 ( 
.A(n_699),
.B(n_250),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_698),
.B(n_583),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_698),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_801),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_656),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_734),
.B(n_583),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_772),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_714),
.B(n_802),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_739),
.B(n_596),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_715),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_725),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_719),
.B(n_596),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_696),
.Y(n_965)
);

BUFx8_ASAP7_75t_SL g966 ( 
.A(n_758),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_732),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_708),
.A2(n_634),
.B(n_623),
.C(n_627),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_742),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_745),
.B(n_596),
.Y(n_970)
);

INVx3_ASAP7_75t_SL g971 ( 
.A(n_772),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_755),
.B(n_623),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_759),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_772),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_760),
.B(n_627),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_775),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_799),
.B(n_367),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_773),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_666),
.B(n_603),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_779),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_696),
.B(n_629),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_667),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_796),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_672),
.Y(n_984)
);

OR2x6_ASAP7_75t_L g985 ( 
.A(n_775),
.B(n_369),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_908),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_923),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_812),
.B(n_705),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_821),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_873),
.B(n_719),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_945),
.A2(n_898),
.B(n_841),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_835),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_873),
.B(n_727),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_SL g994 ( 
.A1(n_865),
.A2(n_933),
.B1(n_855),
.B2(n_842),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_803),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_898),
.A2(n_785),
.B(n_701),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_839),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_814),
.A2(n_659),
.B(n_787),
.C(n_722),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_946),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_917),
.B(n_949),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_921),
.B(n_727),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_957),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_SL g1003 ( 
.A(n_920),
.B(n_254),
.C(n_255),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_904),
.A2(n_670),
.B(n_691),
.C(n_728),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_917),
.B(n_728),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_923),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_SL g1007 ( 
.A(n_925),
.B(n_256),
.C(n_267),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_870),
.B(n_696),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_861),
.B(n_369),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_930),
.A2(n_273),
.B(n_285),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_910),
.A2(n_754),
.B(n_749),
.C(n_741),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_876),
.A2(n_749),
.B(n_741),
.C(n_738),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_910),
.A2(n_738),
.B(n_729),
.C(n_634),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_914),
.A2(n_630),
.B(n_629),
.C(n_636),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_923),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_860),
.A2(n_288),
.B1(n_289),
.B2(n_299),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_871),
.B(n_726),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_884),
.A2(n_300),
.B1(n_370),
.B2(n_636),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_948),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_928),
.B(n_726),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_914),
.A2(n_630),
.B(n_633),
.C(n_370),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_915),
.B(n_931),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_923),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_813),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_921),
.B(n_633),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_851),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_907),
.A2(n_633),
.B(n_726),
.C(n_696),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_892),
.B(n_726),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_930),
.A2(n_633),
.B1(n_600),
.B2(n_607),
.C(n_620),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_838),
.Y(n_1030)
);

CKINVDCx6p67_ASAP7_75t_R g1031 ( 
.A(n_971),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_842),
.A2(n_726),
.B1(n_696),
.B2(n_620),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_948),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_979),
.A2(n_620),
.B(n_607),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_810),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_808),
.B(n_620),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_956),
.B(n_607),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_979),
.A2(n_607),
.B(n_600),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_909),
.A2(n_538),
.B(n_600),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_907),
.A2(n_0),
.B(n_6),
.C(n_7),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_922),
.A2(n_607),
.B(n_600),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_893),
.B(n_600),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_840),
.A2(n_0),
.B(n_8),
.C(n_10),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_813),
.B(n_890),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_953),
.B(n_10),
.C(n_12),
.Y(n_1045)
);

AND2x2_ASAP7_75t_SL g1046 ( 
.A(n_947),
.B(n_959),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_832),
.B(n_14),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_820),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_900),
.A2(n_912),
.B(n_934),
.C(n_867),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_982),
.B(n_854),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_881),
.A2(n_561),
.B(n_538),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_891),
.A2(n_561),
.B(n_500),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_876),
.A2(n_500),
.B(n_561),
.C(n_74),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_840),
.A2(n_17),
.B(n_19),
.C(n_20),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_831),
.B(n_21),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_973),
.B(n_93),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_882),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_826),
.A2(n_863),
.B1(n_805),
.B2(n_849),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_868),
.B(n_96),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_826),
.A2(n_863),
.B1(n_856),
.B2(n_929),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_915),
.B(n_80),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_882),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_927),
.A2(n_500),
.B(n_100),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_831),
.B(n_23),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_834),
.B(n_823),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_955),
.B(n_500),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_848),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_SL g1068 ( 
.A(n_947),
.B(n_959),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_934),
.A2(n_27),
.B(n_28),
.C(n_32),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_811),
.B(n_500),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_830),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_817),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_824),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_984),
.B(n_68),
.Y(n_1074)
);

AND2x2_ASAP7_75t_SL g1075 ( 
.A(n_943),
.B(n_28),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_819),
.A2(n_827),
.B(n_906),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_819),
.A2(n_106),
.B(n_161),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_943),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_811),
.B(n_32),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_883),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_845),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_883),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_SL g1084 ( 
.A(n_926),
.B(n_33),
.C(n_37),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_942),
.B(n_108),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_866),
.A2(n_67),
.B(n_156),
.C(n_152),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_865),
.A2(n_63),
.B1(n_150),
.B2(n_147),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_850),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_853),
.B(n_37),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_974),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_977),
.A2(n_38),
.B(n_41),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_847),
.A2(n_38),
.B(n_41),
.C(n_44),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_966),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_974),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_924),
.A2(n_113),
.B(n_130),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_816),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_974),
.B(n_61),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_866),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_937),
.A2(n_954),
.B(n_939),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_857),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_883),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_919),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_971),
.B(n_116),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_825),
.B(n_47),
.C(n_48),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_818),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_852),
.B(n_129),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_852),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_951),
.A2(n_163),
.B(n_869),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_903),
.B(n_825),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_836),
.B(n_983),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_847),
.B(n_940),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_836),
.B(n_865),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_918),
.A2(n_872),
.B(n_846),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_895),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_976),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_889),
.A2(n_944),
.B(n_952),
.C(n_968),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_889),
.B(n_897),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_958),
.A2(n_961),
.B1(n_950),
.B2(n_936),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_976),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_872),
.B(n_829),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_962),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_958),
.A2(n_961),
.B1(n_950),
.B2(n_936),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_856),
.A2(n_886),
.B1(n_899),
.B2(n_905),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_858),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_886),
.A2(n_899),
.B1(n_905),
.B2(n_828),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_894),
.A2(n_896),
.B(n_837),
.C(n_980),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_875),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_897),
.B(n_815),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1120),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_996),
.A2(n_877),
.B(n_809),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1099),
.A2(n_822),
.B(n_864),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_989),
.B(n_911),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1065),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1050),
.B(n_940),
.Y(n_1136)
);

CKINVDCx11_ASAP7_75t_R g1137 ( 
.A(n_1105),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1006),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1009),
.B(n_874),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1011),
.A2(n_1013),
.B(n_1117),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_989),
.B(n_874),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1055),
.B(n_888),
.C(n_969),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1024),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1000),
.B(n_833),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1076),
.A2(n_991),
.B(n_1125),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1064),
.A2(n_888),
.B(n_965),
.C(n_941),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1060),
.A2(n_932),
.A3(n_938),
.B(n_880),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1114),
.Y(n_1149)
);

OAI22x1_ASAP7_75t_L g1150 ( 
.A1(n_1087),
.A2(n_1112),
.B1(n_1124),
.B2(n_1119),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_995),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1030),
.B(n_862),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1111),
.A2(n_833),
.B1(n_806),
.B2(n_815),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_1044),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1034),
.A2(n_901),
.B(n_902),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1067),
.B(n_967),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1125),
.A2(n_985),
.B1(n_941),
.B2(n_885),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1060),
.A2(n_975),
.A3(n_972),
.B(n_970),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1038),
.A2(n_902),
.B(n_913),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1049),
.A2(n_844),
.B(n_843),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1022),
.B(n_985),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1071),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1006),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1123),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1128),
.A2(n_913),
.B(n_901),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1081),
.B(n_963),
.Y(n_1166)
);

BUFx8_ASAP7_75t_L g1167 ( 
.A(n_1115),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1109),
.A2(n_964),
.B(n_916),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1057),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_993),
.B(n_806),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1127),
.A2(n_964),
.B(n_916),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1027),
.A2(n_859),
.B(n_935),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1012),
.A2(n_960),
.B(n_878),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_997),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_988),
.B(n_804),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1127),
.A2(n_985),
.B1(n_885),
.B2(n_883),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1058),
.A2(n_885),
.B1(n_807),
.B2(n_879),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_887),
.B(n_978),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1058),
.A2(n_885),
.B(n_981),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_SL g1180 ( 
.A(n_1010),
.B(n_862),
.C(n_911),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1006),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1014),
.A2(n_878),
.B(n_981),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1108),
.B(n_879),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1015),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_SL g1186 ( 
.A1(n_1074),
.A2(n_1054),
.B(n_1043),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1062),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1026),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1091),
.A2(n_1016),
.B1(n_1092),
.B2(n_1040),
.C(n_1104),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1035),
.Y(n_1191)
);

NOR4xp25_ASAP7_75t_L g1192 ( 
.A(n_1098),
.B(n_1069),
.C(n_1091),
.D(n_1079),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1004),
.A2(n_1089),
.B(n_990),
.C(n_1122),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1072),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1073),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1074),
.C(n_1017),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1037),
.A2(n_1042),
.B(n_1063),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1118),
.A2(n_1008),
.B(n_1028),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_998),
.A2(n_1029),
.B(n_1042),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1021),
.A2(n_1086),
.B(n_1053),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1047),
.A2(n_994),
.B(n_1102),
.Y(n_1201)
);

NOR4xp25_ASAP7_75t_L g1202 ( 
.A(n_1018),
.B(n_1085),
.C(n_1106),
.D(n_1056),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_SL g1203 ( 
.A1(n_1077),
.A2(n_1095),
.B(n_1037),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1088),
.Y(n_1204)
);

AO32x2_ASAP7_75t_L g1205 ( 
.A1(n_1018),
.A2(n_1084),
.A3(n_987),
.B1(n_1121),
.B2(n_1116),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_987),
.B(n_1023),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1015),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1075),
.B(n_1046),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1045),
.B(n_1003),
.C(n_1007),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1036),
.B(n_1129),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1101),
.A2(n_1070),
.B(n_1066),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1068),
.B(n_1061),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1126),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1025),
.B(n_986),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_999),
.B(n_1002),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1130),
.A2(n_1032),
.B(n_1083),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1019),
.B(n_1033),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1096),
.Y(n_1218)
);

INVx3_ASAP7_75t_SL g1219 ( 
.A(n_1031),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1061),
.A2(n_1068),
.B(n_1022),
.C(n_1100),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1097),
.A2(n_1059),
.B(n_1080),
.Y(n_1221)
);

AND2x4_ASAP7_75t_SL g1222 ( 
.A(n_1023),
.B(n_1121),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1078),
.Y(n_1223)
);

AOI31xp67_ASAP7_75t_L g1224 ( 
.A1(n_1097),
.A2(n_1101),
.A3(n_1059),
.B(n_1020),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1059),
.B(n_1097),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1078),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_1107),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1078),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1093),
.B(n_1082),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1082),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1082),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1103),
.A2(n_1051),
.B(n_1109),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_R g1233 ( 
.A(n_1024),
.B(n_576),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_989),
.B(n_697),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_989),
.B(n_821),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1050),
.B(n_949),
.Y(n_1236)
);

CKINVDCx8_ASAP7_75t_R g1237 ( 
.A(n_1024),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1055),
.B(n_690),
.C(n_1064),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1039),
.A2(n_1076),
.B(n_1041),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_1011),
.B(n_1013),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_992),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_992),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_SL g1243 ( 
.A(n_1024),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_995),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_992),
.Y(n_1245)
);

AND3x1_ASAP7_75t_L g1246 ( 
.A(n_1084),
.B(n_825),
.C(n_690),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1099),
.A2(n_1011),
.B(n_1013),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_996),
.A2(n_898),
.B(n_1099),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1022),
.B(n_1081),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_690),
.C(n_736),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1076),
.A2(n_1117),
.B(n_1051),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1050),
.B(n_334),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_987),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_690),
.C(n_736),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1039),
.A2(n_1076),
.B(n_1041),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1125),
.A2(n_1127),
.B1(n_1060),
.B2(n_898),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_992),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1111),
.A2(n_1050),
.B1(n_1124),
.B2(n_1119),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1050),
.B(n_949),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1125),
.A2(n_1127),
.B1(n_1060),
.B2(n_898),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_690),
.C(n_736),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_989),
.B(n_1000),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1050),
.B(n_334),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_996),
.A2(n_898),
.B(n_1099),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1050),
.B(n_949),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_996),
.A2(n_898),
.B(n_1099),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1050),
.B(n_949),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1099),
.A2(n_1011),
.B(n_1013),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_989),
.B(n_1000),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_989),
.B(n_697),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1022),
.B(n_1081),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_992),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_987),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_996),
.A2(n_898),
.B(n_1099),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1050),
.B(n_949),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1076),
.A2(n_1117),
.B(n_1051),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1238),
.B(n_1250),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1254),
.A2(n_1261),
.B(n_1238),
.C(n_1193),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1208),
.A2(n_1187),
.B1(n_1212),
.B2(n_1234),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1169),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1179),
.B(n_1221),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1196),
.A2(n_1147),
.B(n_1220),
.C(n_1190),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1256),
.A2(n_1260),
.A3(n_1146),
.B(n_1264),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1195),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1149),
.A2(n_1255),
.B(n_1239),
.Y(n_1285)
);

INVx6_ASAP7_75t_L g1286 ( 
.A(n_1181),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1137),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1252),
.A2(n_1263),
.B1(n_1246),
.B2(n_1201),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1132),
.A2(n_1266),
.B(n_1248),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1148),
.Y(n_1291)
);

OAI211xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1136),
.A2(n_1141),
.B(n_1270),
.C(n_1236),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1181),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1235),
.B(n_1246),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1155),
.A2(n_1159),
.B(n_1197),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1186),
.A2(n_1201),
.B(n_1172),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1259),
.B(n_1265),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1151),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1267),
.B(n_1275),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1185),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1192),
.A2(n_1141),
.B1(n_1256),
.B2(n_1260),
.C(n_1258),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1140),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_L g1303 ( 
.A(n_1209),
.B(n_1143),
.C(n_1192),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1178),
.A2(n_1168),
.B(n_1133),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1162),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1244),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1183),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1224),
.B(n_1225),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1237),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1175),
.B(n_1249),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1241),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1240),
.A2(n_1247),
.B(n_1268),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1199),
.A2(n_1157),
.B(n_1214),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1200),
.A2(n_1203),
.B(n_1232),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1209),
.A2(n_1180),
.B1(n_1134),
.B2(n_1150),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1183),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1204),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1139),
.B(n_1145),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1251),
.A2(n_1276),
.B(n_1171),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1143),
.B(n_1142),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1271),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1211),
.A2(n_1160),
.B(n_1216),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1242),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1251),
.A2(n_1276),
.B(n_1165),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1185),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1152),
.A2(n_1161),
.B1(n_1218),
.B2(n_1271),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1198),
.A2(n_1173),
.B(n_1177),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1156),
.B(n_1166),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1153),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1257),
.Y(n_1331)
);

AOI21xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1219),
.A2(n_1144),
.B(n_1229),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1188),
.A2(n_1170),
.B1(n_1164),
.B2(n_1272),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1210),
.A2(n_1189),
.B(n_1174),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1138),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1194),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1202),
.B(n_1191),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1148),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1138),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1215),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1213),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1217),
.A2(n_1184),
.B(n_1227),
.C(n_1206),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1228),
.B(n_1230),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1243),
.B(n_1154),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1182),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1138),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1253),
.A2(n_1273),
.B(n_1158),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1226),
.B(n_1223),
.Y(n_1349)
);

NOR2x1_ASAP7_75t_SL g1350 ( 
.A(n_1163),
.B(n_1207),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1131),
.B(n_1273),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1131),
.B(n_1253),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1205),
.A2(n_1222),
.B(n_1163),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1205),
.A2(n_1163),
.B(n_1207),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1207),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1167),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1223),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1238),
.A2(n_1075),
.B1(n_554),
.B2(n_354),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1220),
.B(n_1212),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1220),
.B(n_1212),
.Y(n_1360)
);

OAI222xp33_ASAP7_75t_L g1361 ( 
.A1(n_1256),
.A2(n_1260),
.B1(n_1092),
.B2(n_1087),
.C1(n_1040),
.C2(n_1054),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1245),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1245),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1187),
.B(n_1235),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1245),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1149),
.A2(n_1255),
.B(n_1239),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_L g1367 ( 
.A(n_1135),
.B(n_744),
.Y(n_1367)
);

NAND2x1p5_ASAP7_75t_L g1368 ( 
.A(n_1181),
.B(n_1101),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1245),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1181),
.B(n_1101),
.Y(n_1370)
);

BUFx2_ASAP7_75t_R g1371 ( 
.A(n_1237),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1256),
.A2(n_1260),
.A3(n_1146),
.B(n_1248),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1238),
.A2(n_1190),
.B1(n_1091),
.B2(n_1104),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1149),
.A2(n_1255),
.B(n_1239),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1183),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1248),
.A2(n_1274),
.B(n_1266),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1235),
.B(n_989),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1238),
.B(n_1250),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1248),
.A2(n_1274),
.B(n_1266),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_SL g1380 ( 
.A(n_1238),
.B(n_928),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1181),
.B(n_1101),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1187),
.B(n_1235),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1261),
.C(n_1238),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1238),
.A2(n_457),
.B1(n_354),
.B2(n_357),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1181),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1245),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1233),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1245),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1161),
.B(n_1271),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1256),
.A2(n_1260),
.A3(n_1146),
.B(n_1248),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1245),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1187),
.B(n_1235),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1245),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1219),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1135),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1238),
.A2(n_1190),
.B1(n_1091),
.B2(n_1104),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1149),
.A2(n_1255),
.B(n_1239),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1261),
.C(n_1238),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1262),
.B(n_1269),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1381),
.B(n_1394),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1294),
.B(n_1311),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1377),
.B(n_1306),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1278),
.A2(n_1400),
.B(n_1384),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1346),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1384),
.A2(n_1277),
.B(n_1378),
.C(n_1400),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1364),
.B(n_1383),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1393),
.B(n_1277),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_L g1411 ( 
.A1(n_1361),
.A2(n_1278),
.B(n_1378),
.C(n_1337),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1346),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1291),
.Y(n_1413)
);

O2A1O1Ixp5_ASAP7_75t_L g1414 ( 
.A1(n_1361),
.A2(n_1337),
.B(n_1380),
.C(n_1303),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1358),
.A2(n_1288),
.B1(n_1373),
.B2(n_1398),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1289),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1359),
.A2(n_1360),
.B(n_1338),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1319),
.B(n_1401),
.Y(n_1418)
);

NOR2x1_ASAP7_75t_L g1419 ( 
.A(n_1292),
.B(n_1321),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1358),
.A2(n_1373),
.B1(n_1398),
.B2(n_1316),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1376),
.A2(n_1379),
.B(n_1320),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1280),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1292),
.B(n_1279),
.Y(n_1423)
);

O2A1O1Ixp5_ASAP7_75t_L g1424 ( 
.A1(n_1359),
.A2(n_1360),
.B(n_1325),
.C(n_1320),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1385),
.A2(n_1327),
.B1(n_1301),
.B2(n_1367),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1329),
.B(n_1321),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1388),
.B(n_1343),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1390),
.B(n_1322),
.Y(n_1430)
);

OR2x2_ASAP7_75t_SL g1431 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1431)
);

AOI211xp5_ASAP7_75t_L g1432 ( 
.A1(n_1282),
.A2(n_1332),
.B(n_1333),
.C(n_1307),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1286),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1298),
.A2(n_1388),
.B1(n_1397),
.B2(n_1284),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1298),
.A2(n_1318),
.B1(n_1281),
.B2(n_1302),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1348),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1281),
.A2(n_1324),
.B1(n_1312),
.B2(n_1331),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1362),
.B(n_1365),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1368),
.A2(n_1382),
.B(n_1370),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1309),
.B(n_1362),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1340),
.B(n_1363),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1334),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1290),
.A2(n_1323),
.B(n_1304),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1334),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1281),
.A2(n_1371),
.B1(n_1309),
.B2(n_1387),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1330),
.A2(n_1313),
.B(n_1353),
.C(n_1354),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1287),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1365),
.B(n_1395),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1369),
.A2(n_1392),
.B1(n_1313),
.B2(n_1342),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1336),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1296),
.A2(n_1314),
.B(n_1342),
.C(n_1356),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1300),
.A2(n_1396),
.B1(n_1395),
.B2(n_1389),
.Y(n_1452)
);

CKINVDCx14_ASAP7_75t_R g1453 ( 
.A(n_1287),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1300),
.A2(n_1345),
.B1(n_1386),
.B2(n_1326),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1341),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1293),
.A2(n_1386),
.B(n_1326),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1293),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1344),
.B(n_1283),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1349),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1310),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1357),
.B(n_1347),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1357),
.B(n_1339),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1283),
.B(n_1372),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1339),
.B(n_1355),
.Y(n_1465)
);

INVxp33_ASAP7_75t_L g1466 ( 
.A(n_1335),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1335),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1335),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1283),
.B(n_1391),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1355),
.B(n_1375),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1315),
.A2(n_1328),
.B(n_1317),
.C(n_1308),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1283),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1308),
.B(n_1350),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1295),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1372),
.A2(n_1391),
.B(n_1366),
.C(n_1374),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1372),
.B(n_1391),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1372),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1391),
.B(n_1285),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1399),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1358),
.A2(n_1238),
.B1(n_1288),
.B2(n_1254),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1376),
.A2(n_1379),
.B(n_1320),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1294),
.B(n_1311),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1358),
.A2(n_1238),
.B1(n_1288),
.B2(n_1254),
.Y(n_1484)
);

AND2x2_ASAP7_75t_SL g1485 ( 
.A(n_1313),
.B(n_1301),
.Y(n_1485)
);

O2A1O1Ixp5_ASAP7_75t_L g1486 ( 
.A1(n_1361),
.A2(n_1250),
.B(n_1261),
.C(n_1254),
.Y(n_1486)
);

O2A1O1Ixp5_ASAP7_75t_L g1487 ( 
.A1(n_1361),
.A2(n_1250),
.B(n_1261),
.C(n_1254),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1294),
.B(n_1311),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1400),
.A2(n_1254),
.B(n_1261),
.C(n_1250),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1400),
.A2(n_1254),
.B(n_1261),
.C(n_1250),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1459),
.B(n_1464),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1485),
.B(n_1428),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1475),
.A2(n_1446),
.B(n_1424),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1469),
.B(n_1406),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1485),
.B(n_1428),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1442),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1444),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1428),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1406),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1476),
.B(n_1440),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1479),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1412),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1410),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1479),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1436),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1426),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1486),
.A2(n_1487),
.B(n_1411),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1415),
.B(n_1420),
.C(n_1480),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1477),
.A2(n_1472),
.B(n_1474),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1421),
.A2(n_1481),
.B(n_1443),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1477),
.A2(n_1414),
.B(n_1478),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1405),
.B(n_1471),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1403),
.B(n_1483),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1450),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1413),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1484),
.A2(n_1419),
.B1(n_1423),
.B2(n_1425),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1481),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1451),
.B(n_1445),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1448),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1407),
.B(n_1427),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1449),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1409),
.B(n_1423),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1402),
.B(n_1418),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1426),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1441),
.B(n_1437),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1443),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1431),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1457),
.B(n_1482),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1438),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1441),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1482),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1489),
.A2(n_1490),
.B1(n_1432),
.B2(n_1422),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1496),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1500),
.B(n_1488),
.Y(n_1538)
);

AOI322xp5_ASAP7_75t_L g1539 ( 
.A1(n_1517),
.A2(n_1453),
.A3(n_1482),
.B1(n_1447),
.B2(n_1461),
.C1(n_1404),
.C2(n_1460),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1493),
.B(n_1473),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1533),
.B(n_1435),
.Y(n_1541)
);

NOR2x1_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1458),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1434),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1506),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1509),
.A2(n_1453),
.B1(n_1468),
.B2(n_1456),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1509),
.A2(n_1447),
.B1(n_1429),
.B2(n_1454),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1416),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1533),
.B(n_1462),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1496),
.Y(n_1552)
);

INVx3_ASAP7_75t_SL g1553 ( 
.A(n_1519),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1494),
.B(n_1416),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1521),
.B(n_1452),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1497),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1529),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1521),
.B(n_1465),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1515),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1506),
.B(n_1470),
.Y(n_1560)
);

NAND2x1_ASAP7_75t_L g1561 ( 
.A(n_1513),
.B(n_1439),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1499),
.B(n_1458),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1508),
.A2(n_1468),
.B1(n_1417),
.B2(n_1430),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1492),
.B(n_1466),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1516),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1510),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1502),
.B(n_1433),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_R g1568 ( 
.A(n_1543),
.B(n_1525),
.Y(n_1568)
);

OAI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1546),
.A2(n_1535),
.B1(n_1508),
.B2(n_1522),
.C(n_1524),
.Y(n_1569)
);

OAI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1563),
.A2(n_1535),
.B1(n_1522),
.B2(n_1524),
.C(n_1519),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1492),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1545),
.A2(n_1519),
.B1(n_1513),
.B2(n_1525),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1545),
.A2(n_1523),
.B1(n_1555),
.B2(n_1541),
.C(n_1528),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1557),
.A2(n_1511),
.B(n_1518),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1552),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1552),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1512),
.Y(n_1577)
);

OAI211xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1539),
.A2(n_1528),
.B(n_1526),
.C(n_1534),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1536),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1538),
.B(n_1495),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1563),
.A2(n_1519),
.B1(n_1513),
.B2(n_1530),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1550),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1495),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_R g1584 ( 
.A(n_1543),
.B(n_1501),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1553),
.A2(n_1519),
.B1(n_1513),
.B2(n_1530),
.Y(n_1585)
);

NAND5xp2_ASAP7_75t_SL g1586 ( 
.A(n_1539),
.B(n_1467),
.C(n_1503),
.D(n_1513),
.E(n_1519),
.Y(n_1586)
);

OAI33xp33_ASAP7_75t_L g1587 ( 
.A1(n_1541),
.A2(n_1555),
.A3(n_1565),
.B1(n_1567),
.B2(n_1558),
.B3(n_1559),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1536),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1558),
.A2(n_1530),
.B1(n_1514),
.B2(n_1534),
.C(n_1503),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1551),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1553),
.A2(n_1527),
.B1(n_1507),
.B2(n_1531),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_SL g1593 ( 
.A(n_1566),
.B(n_1531),
.Y(n_1593)
);

NAND4xp25_ASAP7_75t_L g1594 ( 
.A(n_1542),
.B(n_1520),
.C(n_1514),
.D(n_1501),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1549),
.B(n_1498),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1551),
.Y(n_1597)
);

AND2x2_ASAP7_75t_SL g1598 ( 
.A(n_1566),
.B(n_1493),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1548),
.B(n_1554),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1553),
.A2(n_1531),
.B1(n_1507),
.B2(n_1527),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1565),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1579),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1574),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1603),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1591),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1575),
.Y(n_1608)
);

INVx4_ASAP7_75t_SL g1609 ( 
.A(n_1591),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

AO21x1_ASAP7_75t_L g1611 ( 
.A1(n_1568),
.A2(n_1561),
.B(n_1540),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1588),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1575),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1590),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1597),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1597),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1572),
.B(n_1581),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1596),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1594),
.B(n_1561),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1602),
.B(n_1531),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1571),
.B(n_1544),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1596),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1627)
);

INVx4_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1576),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1576),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1606),
.Y(n_1631)
);

NOR3xp33_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1569),
.C(n_1570),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1606),
.B(n_1589),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1623),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1604),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1608),
.B(n_1600),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1610),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1608),
.B(n_1599),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1607),
.Y(n_1642)
);

OAI33xp33_ASAP7_75t_L g1643 ( 
.A1(n_1629),
.A2(n_1578),
.A3(n_1577),
.B1(n_1547),
.B2(n_1567),
.B3(n_1562),
.Y(n_1643)
);

INVx5_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1615),
.B(n_1580),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1620),
.A2(n_1572),
.B(n_1598),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1628),
.B(n_1583),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1610),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1583),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1613),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1607),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1628),
.B(n_1601),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1605),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1610),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1616),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1605),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1625),
.B(n_1595),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1587),
.C(n_1618),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1610),
.B(n_1598),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1647),
.B(n_1628),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1625),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1607),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1657),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1645),
.B(n_1631),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1662),
.B(n_1627),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1547),
.Y(n_1672)
);

AOI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1646),
.A2(n_1611),
.B(n_1622),
.C(n_1619),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1642),
.B(n_1627),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1635),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1646),
.B(n_1598),
.C(n_1585),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1651),
.B(n_1618),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1637),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1634),
.A2(n_1592),
.B(n_1626),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1630),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1637),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1638),
.B(n_1636),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1638),
.B(n_1636),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1639),
.B(n_1626),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1609),
.Y(n_1691)
);

CKINVDCx16_ASAP7_75t_R g1692 ( 
.A(n_1636),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1650),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1663),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1660),
.B(n_1609),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1655),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1624),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1641),
.B(n_1617),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1668),
.B(n_1641),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1697),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1684),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1664),
.Y(n_1703)
);

NAND3x1_ASAP7_75t_SL g1704 ( 
.A(n_1689),
.B(n_1586),
.C(n_1611),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1677),
.A2(n_1586),
.B1(n_1644),
.B2(n_1624),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1668),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1678),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1697),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1690),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1666),
.B(n_1652),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1673),
.B(n_1666),
.C(n_1671),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1667),
.B(n_1652),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1654),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1694),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1664),
.B(n_1663),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1679),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1680),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1670),
.B(n_1663),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1672),
.B(n_1654),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1694),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1655),
.B(n_1659),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1682),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1702),
.B(n_1708),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1702),
.B(n_1674),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1703),
.B(n_1670),
.Y(n_1729)
);

OAI32xp33_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1692),
.A3(n_1694),
.B1(n_1696),
.B2(n_1698),
.Y(n_1730)
);

OAI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1713),
.A2(n_1584),
.B1(n_1644),
.B2(n_1624),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1703),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1707),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1703),
.B(n_1676),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1706),
.A2(n_1687),
.B1(n_1688),
.B2(n_1676),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1701),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1688),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1711),
.A2(n_1718),
.B1(n_1721),
.B2(n_1714),
.Y(n_1741)
);

XNOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1719),
.B(n_1691),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1717),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1701),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1726),
.B(n_1719),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1743),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1733),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1721),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1743),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1732),
.B(n_1711),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1734),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1728),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1740),
.B(n_1705),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1741),
.B(n_1710),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1733),
.B(n_1710),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1755),
.A2(n_1730),
.B(n_1756),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1727),
.C(n_1737),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1747),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1749),
.B(n_1742),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1748),
.A2(n_1731),
.B1(n_1724),
.B2(n_1716),
.C(n_1735),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1757),
.A2(n_1731),
.B(n_1724),
.C(n_1716),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1752),
.A2(n_1724),
.B1(n_1644),
.B2(n_1718),
.Y(n_1764)
);

OAI21xp33_ASAP7_75t_L g1765 ( 
.A1(n_1752),
.A2(n_1721),
.B(n_1718),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1751),
.B(n_1700),
.C(n_1715),
.D(n_1720),
.Y(n_1766)
);

AOI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1757),
.A2(n_1715),
.B1(n_1722),
.B2(n_1720),
.C1(n_1712),
.C2(n_1725),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1753),
.B(n_1717),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1758),
.A2(n_1750),
.B1(n_1724),
.B2(n_1754),
.C(n_1725),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1762),
.A2(n_1761),
.B1(n_1764),
.B2(n_1765),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1763),
.A2(n_1738),
.B(n_1736),
.Y(n_1771)
);

AOI21xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1759),
.A2(n_1700),
.B(n_1744),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1717),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1767),
.C(n_1766),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1773),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1774),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1772),
.B(n_1745),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1770),
.A2(n_1691),
.B(n_1712),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1771),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1775),
.A2(n_1723),
.B1(n_1709),
.B2(n_1722),
.Y(n_1781)
);

NOR2x1_ASAP7_75t_R g1782 ( 
.A(n_1776),
.B(n_1644),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1778),
.B(n_1681),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1777),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1723),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1785),
.B(n_1779),
.Y(n_1786)
);

NOR2x1_ASAP7_75t_L g1787 ( 
.A(n_1784),
.B(n_1723),
.Y(n_1787)
);

NOR3xp33_ASAP7_75t_L g1788 ( 
.A(n_1782),
.B(n_1723),
.C(n_1704),
.Y(n_1788)
);

XNOR2xp5_ASAP7_75t_L g1789 ( 
.A(n_1786),
.B(n_1781),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1789),
.A2(n_1787),
.B1(n_1783),
.B2(n_1788),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1709),
.B1(n_1648),
.B2(n_1640),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1790),
.Y(n_1792)
);

AO221x1_ASAP7_75t_L g1793 ( 
.A1(n_1792),
.A2(n_1648),
.B1(n_1640),
.B2(n_1695),
.C(n_1693),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1791),
.Y(n_1794)
);

AOI22x1_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1640),
.B1(n_1648),
.B2(n_1686),
.Y(n_1795)
);

XNOR2xp5_ASAP7_75t_L g1796 ( 
.A(n_1793),
.B(n_1704),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1796),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1797),
.B(n_1795),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1699),
.B(n_1659),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1699),
.B(n_1659),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1648),
.B1(n_1640),
.B2(n_1656),
.C(n_1655),
.Y(n_1801)
);

AOI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1656),
.B(n_1685),
.C(n_1658),
.Y(n_1802)
);


endmodule