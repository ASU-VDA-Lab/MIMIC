module fake_netlist_6_2603_n_19810 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_19810);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_19810;

wire n_5643;
wire n_18652;
wire n_2817;
wire n_18318;
wire n_2576;
wire n_1674;
wire n_16664;
wire n_19057;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_4251;
wire n_11111;
wire n_7933;
wire n_578;
wire n_4395;
wire n_19613;
wire n_1061;
wire n_16335;
wire n_5653;
wire n_4978;
wire n_13125;
wire n_3088;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_17647;
wire n_8899;
wire n_5345;
wire n_17634;
wire n_10053;
wire n_1930;
wire n_19785;
wire n_8534;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_19715;
wire n_17991;
wire n_15665;
wire n_19382;
wire n_1555;
wire n_17735;
wire n_19161;
wire n_7161;
wire n_19232;
wire n_830;
wire n_7868;
wire n_15764;
wire n_5725;
wire n_447;
wire n_5229;
wire n_3427;
wire n_18903;
wire n_18105;
wire n_5101;
wire n_3071;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_19220;
wire n_14341;
wire n_10392;
wire n_15074;
wire n_5545;
wire n_2321;
wire n_15253;
wire n_4501;
wire n_9626;
wire n_5598;
wire n_19097;
wire n_15898;
wire n_18013;
wire n_7389;
wire n_10719;
wire n_5259;
wire n_6913;
wire n_10015;
wire n_6948;
wire n_3929;
wire n_3048;
wire n_9362;
wire n_7401;
wire n_7516;
wire n_12767;
wire n_16095;
wire n_18502;
wire n_5930;
wire n_9658;
wire n_1971;
wire n_5354;
wire n_8426;
wire n_5908;
wire n_953;
wire n_19755;
wire n_3664;
wire n_13681;
wire n_5420;
wire n_17209;
wire n_6243;
wire n_4414;
wire n_6585;
wire n_16553;
wire n_18122;
wire n_2625;
wire n_11543;
wire n_4646;
wire n_7651;
wire n_2843;
wire n_3760;
wire n_14662;
wire n_13247;
wire n_16286;
wire n_7956;
wire n_7369;
wire n_16549;
wire n_15421;
wire n_5136;
wire n_15964;
wire n_5638;
wire n_9100;
wire n_6784;
wire n_18310;
wire n_10868;
wire n_9067;
wire n_6323;
wire n_17847;
wire n_14431;
wire n_17478;
wire n_13515;
wire n_6110;
wire n_1967;
wire n_11684;
wire n_16324;
wire n_14410;
wire n_15800;
wire n_9400;
wire n_1911;
wire n_13139;
wire n_7774;
wire n_15600;
wire n_16267;
wire n_6951;
wire n_15899;
wire n_279;
wire n_18317;
wire n_2735;
wire n_13729;
wire n_4671;
wire n_18709;
wire n_14813;
wire n_4314;
wire n_18002;
wire n_323;
wire n_14628;
wire n_8421;
wire n_1381;
wire n_331;
wire n_2093;
wire n_18863;
wire n_17854;
wire n_10114;
wire n_10357;
wire n_15762;
wire n_2770;
wire n_16351;
wire n_15883;
wire n_17706;
wire n_8389;
wire n_2917;
wire n_13711;
wire n_16721;
wire n_12742;
wire n_3923;
wire n_11768;
wire n_9267;
wire n_939;
wire n_19401;
wire n_9652;
wire n_5493;
wire n_8849;
wire n_9059;
wire n_15332;
wire n_5346;
wire n_5252;
wire n_3446;
wire n_18445;
wire n_5309;
wire n_1895;
wire n_4698;
wire n_16254;
wire n_7564;
wire n_3859;
wire n_14989;
wire n_17564;
wire n_10204;
wire n_6383;
wire n_3397;
wire n_18669;
wire n_11637;
wire n_3575;
wire n_8151;
wire n_2469;
wire n_9038;
wire n_16004;
wire n_8748;
wire n_13984;
wire n_5452;
wire n_6794;
wire n_18608;
wire n_8718;
wire n_2764;
wire n_9935;
wire n_6990;
wire n_14288;
wire n_14824;
wire n_18699;
wire n_8223;
wire n_4856;
wire n_3492;
wire n_9135;
wire n_16800;
wire n_13771;
wire n_18644;
wire n_11295;
wire n_4291;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_2434;
wire n_9070;
wire n_11708;
wire n_15629;
wire n_14401;
wire n_10827;
wire n_3247;
wire n_5922;
wire n_14922;
wire n_12158;
wire n_7823;
wire n_9477;
wire n_7062;
wire n_7569;
wire n_14769;
wire n_355;
wire n_14961;
wire n_8577;
wire n_8594;
wire n_8428;
wire n_9829;
wire n_13341;
wire n_2254;
wire n_5058;
wire n_10685;
wire n_1926;
wire n_17139;
wire n_15185;
wire n_12083;
wire n_12014;
wire n_14803;
wire n_19270;
wire n_1747;
wire n_16035;
wire n_10607;
wire n_15490;
wire n_18033;
wire n_5042;
wire n_19569;
wire n_8164;
wire n_4072;
wire n_835;
wire n_928;
wire n_15100;
wire n_10368;
wire n_19137;
wire n_9088;
wire n_10183;
wire n_17161;
wire n_6952;
wire n_11464;
wire n_19421;
wire n_3997;
wire n_14878;
wire n_15046;
wire n_2468;
wire n_5144;
wire n_10383;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_13550;
wire n_17601;
wire n_13348;
wire n_2812;
wire n_10724;
wire n_16398;
wire n_19396;
wire n_9988;
wire n_7009;
wire n_2136;
wire n_2409;
wire n_3834;
wire n_11553;
wire n_12795;
wire n_2075;
wire n_10876;
wire n_18780;
wire n_9137;
wire n_14043;
wire n_11180;
wire n_18820;
wire n_3192;
wire n_8995;
wire n_1546;
wire n_4394;
wire n_6010;
wire n_3352;
wire n_8711;
wire n_12505;
wire n_18602;
wire n_2150;
wire n_4082;
wire n_1420;
wire n_13721;
wire n_18430;
wire n_10820;
wire n_13514;
wire n_8306;
wire n_7488;
wire n_2558;
wire n_13194;
wire n_8887;
wire n_18677;
wire n_16183;
wire n_4289;
wire n_11866;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_15659;
wire n_1487;
wire n_9578;
wire n_13109;
wire n_7438;
wire n_16631;
wire n_14355;
wire n_7337;
wire n_9489;
wire n_14123;
wire n_5957;
wire n_10728;
wire n_6357;
wire n_925;
wire n_6800;
wire n_18962;
wire n_4322;
wire n_10655;
wire n_9797;
wire n_1249;
wire n_2693;
wire n_8332;
wire n_9478;
wire n_2767;
wire n_11379;
wire n_16627;
wire n_19571;
wire n_19659;
wire n_10670;
wire n_5929;
wire n_5787;
wire n_11981;
wire n_19181;
wire n_9351;
wire n_5445;
wire n_14556;
wire n_6839;
wire n_532;
wire n_173;
wire n_9189;
wire n_413;
wire n_18888;
wire n_16528;
wire n_2170;
wire n_4156;
wire n_14701;
wire n_7098;
wire n_16587;
wire n_18936;
wire n_3158;
wire n_1788;
wire n_8921;
wire n_9356;
wire n_15880;
wire n_16499;
wire n_1835;
wire n_5076;
wire n_18328;
wire n_5870;
wire n_9175;
wire n_6508;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_4310;
wire n_7782;
wire n_5212;
wire n_13385;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_16339;
wire n_1246;
wire n_4528;
wire n_899;
wire n_13992;
wire n_17429;
wire n_19103;
wire n_13790;
wire n_4914;
wire n_499;
wire n_3418;
wire n_705;
wire n_1004;
wire n_10624;
wire n_13304;
wire n_14633;
wire n_15699;
wire n_11900;
wire n_2297;
wire n_5901;
wire n_6538;
wire n_5599;
wire n_12883;
wire n_5324;
wire n_2103;
wire n_8983;
wire n_10422;
wire n_3770;
wire n_9818;
wire n_4402;
wire n_927;
wire n_16503;
wire n_18974;
wire n_12367;
wire n_17360;
wire n_5009;
wire n_13526;
wire n_12563;
wire n_7243;
wire n_13321;
wire n_15042;
wire n_15519;
wire n_14722;
wire n_13427;
wire n_4627;
wire n_4079;
wire n_9909;
wire n_19607;
wire n_8620;
wire n_19204;
wire n_15264;
wire n_13270;
wire n_10052;
wire n_10109;
wire n_18151;
wire n_3390;
wire n_19582;
wire n_10448;
wire n_11196;
wire n_16239;
wire n_11963;
wire n_16334;
wire n_9571;
wire n_8424;
wire n_2137;
wire n_16003;
wire n_4798;
wire n_2532;
wire n_12655;
wire n_7941;
wire n_16096;
wire n_18628;
wire n_11483;
wire n_15067;
wire n_19591;
wire n_19345;
wire n_5089;
wire n_13356;
wire n_2849;
wire n_14912;
wire n_1398;
wire n_884;
wire n_19177;
wire n_731;
wire n_8907;
wire n_11080;
wire n_958;
wire n_5137;
wire n_17557;
wire n_14079;
wire n_15168;
wire n_9894;
wire n_8324;
wire n_15411;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7913;
wire n_15144;
wire n_5288;
wire n_3606;
wire n_819;
wire n_14224;
wire n_2788;
wire n_10380;
wire n_6449;
wire n_18687;
wire n_18273;
wire n_3892;
wire n_6461;
wire n_4069;
wire n_14682;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_9033;
wire n_2331;
wire n_15031;
wire n_12933;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_17076;
wire n_13893;
wire n_5947;
wire n_1877;
wire n_2030;
wire n_11946;
wire n_9443;
wire n_9996;
wire n_14950;
wire n_7800;
wire n_13795;
wire n_3026;
wire n_17501;
wire n_14547;
wire n_15416;
wire n_221;
wire n_3847;
wire n_2552;
wire n_17942;
wire n_18735;
wire n_9938;
wire n_7261;
wire n_9023;
wire n_14415;
wire n_11818;
wire n_16298;
wire n_18739;
wire n_6773;
wire n_13569;
wire n_7455;
wire n_18042;
wire n_19105;
wire n_2160;
wire n_9201;
wire n_6531;
wire n_10952;
wire n_2131;
wire n_13628;
wire n_18958;
wire n_9559;
wire n_11803;
wire n_15738;
wire n_16301;
wire n_8015;
wire n_18507;
wire n_1933;
wire n_19102;
wire n_15613;
wire n_14786;
wire n_4411;
wire n_9184;
wire n_13585;
wire n_18418;
wire n_18472;
wire n_8024;
wire n_12562;
wire n_18396;
wire n_4180;
wire n_16531;
wire n_3354;
wire n_11090;
wire n_19035;
wire n_5740;
wire n_5820;
wire n_13266;
wire n_13957;
wire n_9403;
wire n_9875;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_11561;
wire n_5534;
wire n_8003;
wire n_8785;
wire n_3566;
wire n_17826;
wire n_2829;
wire n_8692;
wire n_6889;
wire n_16142;
wire n_9183;
wire n_3804;
wire n_4207;
wire n_14326;
wire n_5196;
wire n_16381;
wire n_10852;
wire n_4470;
wire n_9529;
wire n_3901;
wire n_465;
wire n_11425;
wire n_4704;
wire n_2142;
wire n_4596;
wire n_6478;
wire n_820;
wire n_6100;
wire n_6516;
wire n_17845;
wire n_6977;
wire n_16854;
wire n_17542;
wire n_7660;
wire n_2263;
wire n_6911;
wire n_6599;
wire n_6522;
wire n_17189;
wire n_5660;
wire n_2756;
wire n_5334;
wire n_9347;
wire n_807;
wire n_4761;
wire n_18879;
wire n_16395;
wire n_13603;
wire n_6207;
wire n_6931;
wire n_7948;
wire n_238;
wire n_9082;
wire n_1595;
wire n_8685;
wire n_6963;
wire n_16252;
wire n_4932;
wire n_19358;
wire n_5456;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_19531;
wire n_9445;
wire n_7627;
wire n_9803;
wire n_16698;
wire n_17041;
wire n_7601;
wire n_3195;
wire n_6346;
wire n_4274;
wire n_15729;
wire n_17519;
wire n_5386;
wire n_14737;
wire n_11676;
wire n_12266;
wire n_2595;
wire n_16949;
wire n_12287;
wire n_19713;
wire n_13485;
wire n_12991;
wire n_11134;
wire n_13735;
wire n_8886;
wire n_7211;
wire n_10933;
wire n_5618;
wire n_8506;
wire n_2264;
wire n_6494;
wire n_16365;
wire n_11548;
wire n_13041;
wire n_17037;
wire n_13154;
wire n_7822;
wire n_6453;
wire n_9307;
wire n_10762;
wire n_11342;
wire n_7785;
wire n_1891;
wire n_1213;
wire n_2235;
wire n_11266;
wire n_19706;
wire n_5082;
wire n_5338;
wire n_12479;
wire n_8352;
wire n_18941;
wire n_10360;
wire n_9450;
wire n_2298;
wire n_490;
wire n_3594;
wire n_5689;
wire n_16777;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_4144;
wire n_12537;
wire n_17183;
wire n_9693;
wire n_17582;
wire n_12921;
wire n_2169;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_13686;
wire n_13645;
wire n_16753;
wire n_12215;
wire n_18473;
wire n_9880;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_11546;
wire n_15259;
wire n_16946;
wire n_15460;
wire n_330;
wire n_7158;
wire n_1406;
wire n_13400;
wire n_9905;
wire n_18717;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_13331;
wire n_9456;
wire n_7044;
wire n_9710;
wire n_8623;
wire n_11113;
wire n_18593;
wire n_2518;
wire n_17769;
wire n_19193;
wire n_13812;
wire n_14970;
wire n_7838;
wire n_4842;
wire n_204;
wire n_482;
wire n_4135;
wire n_16969;
wire n_1845;
wire n_12731;
wire n_7518;
wire n_2798;
wire n_6147;
wire n_9199;
wire n_13544;
wire n_7791;
wire n_2753;
wire n_2007;
wire n_2039;
wire n_18172;
wire n_12616;
wire n_1544;
wire n_18333;
wire n_3437;
wire n_4111;
wire n_14375;
wire n_12653;
wire n_533;
wire n_7146;
wire n_18081;
wire n_16580;
wire n_18498;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12587;
wire n_10747;
wire n_13110;
wire n_16628;
wire n_2973;
wire n_9422;
wire n_18344;
wire n_5218;
wire n_12348;
wire n_3665;
wire n_16929;
wire n_273;
wire n_16099;
wire n_15590;
wire n_10843;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_16869;
wire n_3174;
wire n_10997;
wire n_1948;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_19640;
wire n_6073;
wire n_19157;
wire n_6331;
wire n_13498;
wire n_2283;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_18289;
wire n_11408;
wire n_4196;
wire n_2056;
wire n_13183;
wire n_12519;
wire n_17184;
wire n_4902;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_13007;
wire n_2680;
wire n_10112;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_502;
wire n_1257;
wire n_3197;
wire n_7223;
wire n_7833;
wire n_14868;
wire n_5512;
wire n_9297;
wire n_2398;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_18534;
wire n_2695;
wire n_4035;
wire n_7445;
wire n_11086;
wire n_6529;
wire n_1949;
wire n_3759;
wire n_4516;
wire n_1804;
wire n_11710;
wire n_251;
wire n_6290;
wire n_10253;
wire n_6025;
wire n_1337;
wire n_6455;
wire n_15277;
wire n_18435;
wire n_13804;
wire n_12455;
wire n_13099;
wire n_4492;
wire n_19524;
wire n_18516;
wire n_5607;
wire n_7695;
wire n_7179;
wire n_7122;
wire n_12157;
wire n_5999;
wire n_19676;
wire n_6203;
wire n_15806;
wire n_13064;
wire n_7630;
wire n_16246;
wire n_8643;
wire n_15660;
wire n_15357;
wire n_8565;
wire n_10821;
wire n_19784;
wire n_13648;
wire n_4542;
wire n_6892;
wire n_4462;
wire n_15722;
wire n_14181;
wire n_15278;
wire n_18054;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_4931;
wire n_14213;
wire n_17320;
wire n_17885;
wire n_7051;
wire n_8477;
wire n_19766;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_14842;
wire n_13115;
wire n_1291;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_5911;
wire n_11601;
wire n_11971;
wire n_2122;
wire n_12314;
wire n_3503;
wire n_1065;
wire n_11116;
wire n_12604;
wire n_13305;
wire n_1255;
wire n_8876;
wire n_5124;
wire n_19017;
wire n_3951;
wire n_9359;
wire n_14189;
wire n_3874;
wire n_15761;
wire n_5123;
wire n_8060;
wire n_3027;
wire n_4083;
wire n_11124;
wire n_6392;
wire n_182;
wire n_17470;
wire n_15301;
wire n_7351;
wire n_9352;
wire n_2746;
wire n_389;
wire n_7608;
wire n_17053;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_13202;
wire n_15350;
wire n_13638;
wire n_4171;
wire n_17948;
wire n_14392;
wire n_19347;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_10330;
wire n_1461;
wire n_8276;
wire n_2076;
wire n_3567;
wire n_11465;
wire n_8027;
wire n_4705;
wire n_3807;
wire n_17808;
wire n_11265;
wire n_11125;
wire n_1114;
wire n_17244;
wire n_7783;
wire n_13220;
wire n_10276;
wire n_191;
wire n_10594;
wire n_8978;
wire n_8245;
wire n_15072;
wire n_12910;
wire n_18725;
wire n_18215;
wire n_8454;
wire n_2881;
wire n_1116;
wire n_8891;
wire n_1219;
wire n_11690;
wire n_18719;
wire n_19142;
wire n_16194;
wire n_3897;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_6403;
wire n_7947;
wire n_1221;
wire n_16826;
wire n_6491;
wire n_19519;
wire n_16321;
wire n_14072;
wire n_17120;
wire n_11412;
wire n_13039;
wire n_13130;
wire n_10441;
wire n_19500;
wire n_17237;
wire n_5518;
wire n_15671;
wire n_9124;
wire n_6661;
wire n_13719;
wire n_8847;
wire n_14548;
wire n_19099;
wire n_4068;
wire n_10841;
wire n_16076;
wire n_12313;
wire n_18071;
wire n_2743;
wire n_4766;
wire n_14661;
wire n_8356;
wire n_6136;
wire n_16384;
wire n_16416;
wire n_3378;
wire n_15305;
wire n_15588;
wire n_3745;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_5357;
wire n_3523;
wire n_2222;
wire n_13062;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_14130;
wire n_14930;
wire n_5541;
wire n_10576;
wire n_16596;
wire n_334;
wire n_6668;
wire n_2999;
wire n_15548;
wire n_1239;
wire n_3697;
wire n_16714;
wire n_19168;
wire n_2408;
wire n_6859;
wire n_18752;
wire n_13752;
wire n_10237;
wire n_19484;
wire n_13596;
wire n_12889;
wire n_18092;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_9515;
wire n_6971;
wire n_17957;
wire n_9642;
wire n_393;
wire n_14231;
wire n_12385;
wire n_13219;
wire n_5673;
wire n_17449;
wire n_5443;
wire n_6351;
wire n_9382;
wire n_16392;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_19207;
wire n_13295;
wire n_3936;
wire n_1349;
wire n_16906;
wire n_18194;
wire n_17693;
wire n_6829;
wire n_2723;
wire n_17981;
wire n_3496;
wire n_13160;
wire n_15249;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_17337;
wire n_10708;
wire n_13818;
wire n_15024;
wire n_8803;
wire n_3239;
wire n_3902;
wire n_4062;
wire n_18478;
wire n_4396;
wire n_9706;
wire n_3101;
wire n_15174;
wire n_17904;
wire n_3374;
wire n_10387;
wire n_13764;
wire n_19408;
wire n_1552;
wire n_11224;
wire n_8790;
wire n_15569;
wire n_4293;
wire n_10219;
wire n_1031;
wire n_11924;
wire n_15193;
wire n_9591;
wire n_6137;
wire n_14833;
wire n_10364;
wire n_11422;
wire n_8338;
wire n_4412;
wire n_14480;
wire n_12489;
wire n_8491;
wire n_2217;
wire n_4781;
wire n_16610;
wire n_9283;
wire n_19299;
wire n_12030;
wire n_206;
wire n_633;
wire n_12565;
wire n_15236;
wire n_1040;
wire n_3059;
wire n_9468;
wire n_14098;
wire n_14482;
wire n_17174;
wire n_14223;
wire n_15962;
wire n_5424;
wire n_12415;
wire n_3017;
wire n_1805;
wire n_17332;
wire n_10559;
wire n_13173;
wire n_15355;
wire n_15945;
wire n_14848;
wire n_18548;
wire n_7154;
wire n_16232;
wire n_8304;
wire n_19644;
wire n_19012;
wire n_11418;
wire n_6655;
wire n_19694;
wire n_19187;
wire n_3274;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_16122;
wire n_722;
wire n_5613;
wire n_18852;
wire n_14604;
wire n_14735;
wire n_2223;
wire n_1621;
wire n_19572;
wire n_19688;
wire n_13101;
wire n_6786;
wire n_8315;
wire n_16446;
wire n_15885;
wire n_17528;
wire n_18964;
wire n_11040;
wire n_11754;
wire n_14916;
wire n_9756;
wire n_4762;
wire n_192;
wire n_13748;
wire n_11672;
wire n_3113;
wire n_10353;
wire n_10847;
wire n_10451;
wire n_1458;
wire n_15801;
wire n_17778;
wire n_5303;
wire n_12240;
wire n_12003;
wire n_7496;
wire n_223;
wire n_4154;
wire n_12165;
wire n_10866;
wire n_18127;
wire n_9940;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_3844;
wire n_1237;
wire n_11763;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_18730;
wire n_8535;
wire n_10653;
wire n_11587;
wire n_12280;
wire n_13461;
wire n_6373;
wire n_12492;
wire n_19535;
wire n_16282;
wire n_17011;
wire n_2243;
wire n_4898;
wire n_5601;
wire n_13188;
wire n_4819;
wire n_17639;
wire n_7131;
wire n_9586;
wire n_8909;
wire n_3332;
wire n_18977;
wire n_16356;
wire n_11843;
wire n_2570;
wire n_14614;
wire n_4645;
wire n_11629;
wire n_15147;
wire n_9554;
wire n_18246;
wire n_5635;
wire n_17180;
wire n_5091;
wire n_6546;
wire n_4302;
wire n_15927;
wire n_3395;
wire n_7060;
wire n_19439;
wire n_13217;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_16332;
wire n_1711;
wire n_14397;
wire n_17971;
wire n_10853;
wire n_13802;
wire n_18559;
wire n_7761;
wire n_10338;
wire n_12978;
wire n_1422;
wire n_15668;
wire n_15137;
wire n_8496;
wire n_1842;
wire n_12476;
wire n_8568;
wire n_516;
wire n_8852;
wire n_18423;
wire n_12023;
wire n_17655;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_16225;
wire n_16677;
wire n_4606;
wire n_13413;
wire n_6450;
wire n_15153;
wire n_13203;
wire n_2058;
wire n_2660;
wire n_19128;
wire n_14462;
wire n_8456;
wire n_7137;
wire n_4563;
wire n_4962;
wire n_14933;
wire n_5056;
wire n_9920;
wire n_12598;
wire n_9039;
wire n_11854;
wire n_8573;
wire n_2124;
wire n_19070;
wire n_5336;
wire n_5447;
wire n_18623;
wire n_17389;
wire n_13230;
wire n_7743;
wire n_6179;
wire n_19230;
wire n_9125;
wire n_9139;
wire n_17941;
wire n_5747;
wire n_12733;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_808;
wire n_18695;
wire n_14684;
wire n_5753;
wire n_12245;
wire n_15713;
wire n_1193;
wire n_18124;
wire n_14572;
wire n_9972;
wire n_6083;
wire n_12909;
wire n_6434;
wire n_551;
wire n_9157;
wire n_16417;
wire n_3884;
wire n_17880;
wire n_9324;
wire n_5808;
wire n_8807;
wire n_6933;
wire n_8521;
wire n_6547;
wire n_5193;
wire n_9442;
wire n_1481;
wire n_19374;
wire n_6984;
wire n_18394;
wire n_17392;
wire n_10763;
wire n_9957;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_17586;
wire n_5961;
wire n_18757;
wire n_6507;
wire n_9313;
wire n_6687;
wire n_9173;
wire n_6690;
wire n_7412;
wire n_12144;
wire n_9160;
wire n_219;
wire n_9974;
wire n_19365;
wire n_12129;
wire n_14753;
wire n_13658;
wire n_5533;
wire n_14671;
wire n_4257;
wire n_16454;
wire n_17977;
wire n_18441;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_4720;
wire n_14674;
wire n_3857;
wire n_243;
wire n_1873;
wire n_19496;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_12835;
wire n_10129;
wire n_16089;
wire n_1330;
wire n_7523;
wire n_8654;
wire n_2876;
wire n_14229;
wire n_15060;
wire n_11241;
wire n_15520;
wire n_5953;
wire n_14188;
wire n_11508;
wire n_7141;
wire n_5198;
wire n_16139;
wire n_5718;
wire n_6505;
wire n_1663;
wire n_12636;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_1107;
wire n_3294;
wire n_6001;
wire n_11218;
wire n_4502;
wire n_318;
wire n_10195;
wire n_13722;
wire n_3490;
wire n_4849;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_12938;
wire n_13057;
wire n_8367;
wire n_7367;
wire n_3581;
wire n_16439;
wire n_6023;
wire n_14897;
wire n_19251;
wire n_12173;
wire n_6905;
wire n_17520;
wire n_15925;
wire n_18255;
wire n_19275;
wire n_7368;
wire n_429;
wire n_5553;
wire n_8011;
wire n_4066;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_15141;
wire n_12411;
wire n_10280;
wire n_4004;
wire n_5404;
wire n_18634;
wire n_4292;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_9074;
wire n_5549;
wire n_9408;
wire n_267;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_19190;
wire n_12568;
wire n_3280;
wire n_16163;
wire n_13478;
wire n_18256;
wire n_12970;
wire n_1515;
wire n_14295;
wire n_8902;
wire n_7557;
wire n_593;
wire n_7128;
wire n_14367;
wire n_637;
wire n_13915;
wire n_7594;
wire n_15057;
wire n_19479;
wire n_16300;
wire n_19236;
wire n_18288;
wire n_10504;
wire n_2525;
wire n_7788;
wire n_13783;
wire n_5154;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_3889;
wire n_2687;
wire n_2887;
wire n_2194;
wire n_5637;
wire n_1987;
wire n_7586;
wire n_968;
wire n_7767;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_16402;
wire n_13705;
wire n_17986;
wire n_17771;
wire n_9277;
wire n_9257;
wire n_17773;
wire n_2391;
wire n_2431;
wire n_17070;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_18515;
wire n_7744;
wire n_10595;
wire n_7748;
wire n_6827;
wire n_18914;
wire n_11073;
wire n_1208;
wire n_1072;
wire n_815;
wire n_7485;
wire n_18867;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8671;
wire n_19196;
wire n_15313;
wire n_284;
wire n_3436;
wire n_9671;
wire n_1026;
wire n_289;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_12929;
wire n_16065;
wire n_685;
wire n_3240;
wire n_15075;
wire n_12261;
wire n_18007;
wire n_12106;
wire n_5333;
wire n_5594;
wire n_12291;
wire n_14510;
wire n_12124;
wire n_11755;
wire n_9510;
wire n_18055;
wire n_13497;
wire n_15406;
wire n_19529;
wire n_14396;
wire n_2517;
wire n_2713;
wire n_11918;
wire n_11748;
wire n_12433;
wire n_5000;
wire n_5551;
wire n_8701;
wire n_16810;
wire n_6499;
wire n_19678;
wire n_18158;
wire n_12217;
wire n_15922;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_13851;
wire n_9679;
wire n_8645;
wire n_13272;
wire n_18954;
wire n_4688;
wire n_4058;
wire n_3082;
wire n_4848;
wire n_16411;
wire n_19507;
wire n_156;
wire n_16717;
wire n_8824;
wire n_11673;
wire n_2407;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_6276;
wire n_10499;
wire n_8340;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_2667;
wire n_18425;
wire n_1571;
wire n_2948;
wire n_8455;
wire n_7208;
wire n_13613;
wire n_947;
wire n_12185;
wire n_9770;
wire n_1992;
wire n_8681;
wire n_7406;
wire n_11417;
wire n_16044;
wire n_18656;
wire n_3140;
wire n_4749;
wire n_9592;
wire n_5155;
wire n_17507;
wire n_9180;
wire n_10922;
wire n_926;
wire n_19013;
wire n_10718;
wire n_1698;
wire n_4100;
wire n_13821;
wire n_19198;
wire n_13712;
wire n_9625;
wire n_777;
wire n_15041;
wire n_4085;
wire n_15393;
wire n_4464;
wire n_14144;
wire n_6851;
wire n_6460;
wire n_19429;
wire n_4659;
wire n_5217;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_15595;
wire n_8255;
wire n_15081;
wire n_8461;
wire n_6368;
wire n_1857;
wire n_16474;
wire n_6583;
wire n_4866;
wire n_4889;
wire n_3638;
wire n_16940;
wire n_4816;
wire n_17419;
wire n_12520;
wire n_2110;
wire n_1659;
wire n_3393;
wire n_17134;
wire n_3451;
wire n_11459;
wire n_4937;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_16344;
wire n_2053;
wire n_12808;
wire n_4222;
wire n_18275;
wire n_2710;
wire n_6064;
wire n_1966;
wire n_13801;
wire n_5793;
wire n_19286;
wire n_8523;
wire n_12143;
wire n_4976;
wire n_13879;
wire n_5578;
wire n_18064;
wire n_231;
wire n_1457;
wire n_1993;
wire n_11806;
wire n_2617;
wire n_19682;
wire n_1466;
wire n_11050;
wire n_5207;
wire n_17714;
wire n_5676;
wire n_1893;
wire n_4665;
wire n_11484;
wire n_2387;
wire n_19483;
wire n_2846;
wire n_19183;
wire n_10295;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_10336;
wire n_4362;
wire n_7716;
wire n_17903;
wire n_8954;
wire n_12212;
wire n_7540;
wire n_775;
wire n_13231;
wire n_12624;
wire n_1531;
wire n_453;
wire n_8552;
wire n_17412;
wire n_7558;
wire n_4261;
wire n_8373;
wire n_13165;
wire n_426;
wire n_3986;
wire n_12151;
wire n_17407;
wire n_15204;
wire n_2556;
wire n_4747;
wire n_5251;
wire n_18284;
wire n_9970;
wire n_11365;
wire n_18138;
wire n_3175;
wire n_17016;
wire n_16081;
wire n_5475;
wire n_15341;
wire n_4448;
wire n_1096;
wire n_15477;
wire n_6233;
wire n_6377;
wire n_12402;
wire n_17959;
wire n_18782;
wire n_688;
wire n_1077;
wire n_4132;
wire n_10361;
wire n_1437;
wire n_7143;
wire n_10424;
wire n_8965;
wire n_4355;
wire n_18454;
wire n_2276;
wire n_13476;
wire n_2803;
wire n_379;
wire n_18399;
wire n_12162;
wire n_3202;
wire n_602;
wire n_17087;
wire n_7497;
wire n_4655;
wire n_11829;
wire n_11517;
wire n_7793;
wire n_16102;
wire n_587;
wire n_16274;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_13776;
wire n_7248;
wire n_7204;
wire n_15835;
wire n_12852;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_13343;
wire n_7654;
wire n_5132;
wire n_17339;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_5774;
wire n_13907;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_12821;
wire n_14782;
wire n_4024;
wire n_18756;
wire n_7120;
wire n_6335;
wire n_12837;
wire n_8728;
wire n_8386;
wire n_14070;
wire n_14330;
wire n_13491;
wire n_4860;
wire n_18654;
wire n_15748;
wire n_3414;
wire n_17995;
wire n_14235;
wire n_6173;
wire n_14851;
wire n_18012;
wire n_10058;
wire n_16471;
wire n_2563;
wire n_19434;
wire n_4989;
wire n_7757;
wire n_1683;
wire n_17539;
wire n_280;
wire n_6630;
wire n_1187;
wire n_4558;
wire n_8396;
wire n_16560;
wire n_6612;
wire n_6606;
wire n_13450;
wire n_3550;
wire n_19533;
wire n_14178;
wire n_5508;
wire n_12907;
wire n_15500;
wire n_14891;
wire n_17051;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_9028;
wire n_17217;
wire n_4328;
wire n_8020;
wire n_1057;
wire n_9374;
wire n_2785;
wire n_2636;
wire n_13634;
wire n_18027;
wire n_10413;
wire n_3399;
wire n_19268;
wire n_1611;
wire n_2740;
wire n_17786;
wire n_4808;
wire n_5767;
wire n_1589;
wire n_12708;
wire n_4712;
wire n_10369;
wire n_2309;
wire n_6821;
wire n_5462;
wire n_9983;
wire n_6688;
wire n_8580;
wire n_9993;
wire n_3533;
wire n_13622;
wire n_4725;
wire n_11207;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3132;
wire n_16951;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_14794;
wire n_17684;
wire n_9237;
wire n_13931;
wire n_14404;
wire n_6557;
wire n_18302;
wire n_6753;
wire n_18164;
wire n_17151;
wire n_7341;
wire n_4908;
wire n_12088;
wire n_15423;
wire n_14377;
wire n_6639;
wire n_12508;
wire n_12096;
wire n_5150;
wire n_8832;
wire n_3819;
wire n_2050;
wire n_19412;
wire n_19399;
wire n_2164;
wire n_11098;
wire n_15815;
wire n_5179;
wire n_7957;
wire n_10938;
wire n_6627;
wire n_17147;
wire n_3544;
wire n_2904;
wire n_18019;
wire n_10927;
wire n_4616;
wire n_4982;
wire n_370;
wire n_8592;
wire n_11204;
wire n_6190;
wire n_1979;
wire n_2738;
wire n_16920;
wire n_12701;
wire n_10578;
wire n_4323;
wire n_16199;
wire n_19113;
wire n_6615;
wire n_17331;
wire n_2342;
wire n_2167;
wire n_7294;
wire n_4017;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_4739;
wire n_15367;
wire n_19095;
wire n_8104;
wire n_2768;
wire n_18511;
wire n_17428;
wire n_4298;
wire n_2314;
wire n_10746;
wire n_9188;
wire n_16407;
wire n_18009;
wire n_4644;
wire n_19002;
wire n_8779;
wire n_5503;
wire n_5945;
wire n_10697;
wire n_11714;
wire n_16179;
wire n_2390;
wire n_15070;
wire n_1343;
wire n_2734;
wire n_7250;
wire n_8762;
wire n_17503;
wire n_18365;
wire n_17358;
wire n_1900;
wire n_3381;
wire n_13419;
wire n_9207;
wire n_11860;
wire n_17057;
wire n_10926;
wire n_8897;
wire n_11503;
wire n_17104;
wire n_4672;
wire n_8376;
wire n_18271;
wire n_2939;
wire n_18998;
wire n_5749;
wire n_1672;
wire n_15640;
wire n_6271;
wire n_15683;
wire n_16202;
wire n_4598;
wire n_8599;
wire n_13460;
wire n_15451;
wire n_5993;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_13105;
wire n_14467;
wire n_14789;
wire n_13076;
wire n_15526;
wire n_12950;
wire n_8628;
wire n_15150;
wire n_13028;
wire n_8547;
wire n_4424;
wire n_7113;
wire n_1751;
wire n_10433;
wire n_285;
wire n_9116;
wire n_14096;
wire n_11983;
wire n_10839;
wire n_11813;
wire n_3506;
wire n_1928;
wire n_14583;
wire n_4317;
wire n_14893;
wire n_8275;
wire n_6198;
wire n_5418;
wire n_18270;
wire n_6762;
wire n_4088;
wire n_3711;
wire n_9035;
wire n_729;
wire n_16960;
wire n_3642;
wire n_14915;
wire n_4650;
wire n_17780;
wire n_438;
wire n_17075;
wire n_2874;
wire n_1200;
wire n_4967;
wire n_9678;
wire n_8247;
wire n_6577;
wire n_12956;
wire n_17373;
wire n_14856;
wire n_15235;
wire n_4912;
wire n_9284;
wire n_5086;
wire n_4735;
wire n_187;
wire n_3300;
wire n_2978;
wire n_15711;
wire n_1050;
wire n_5170;
wire n_7604;
wire n_3515;
wire n_1150;
wire n_9606;
wire n_17018;
wire n_13459;
wire n_1023;
wire n_1118;
wire n_14268;
wire n_194;
wire n_2949;
wire n_10297;
wire n_12553;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_14127;
wire n_440;
wire n_3806;
wire n_8827;
wire n_2931;
wire n_3866;
wire n_17937;
wire n_9549;
wire n_14894;
wire n_12866;
wire n_17801;
wire n_4157;
wire n_6845;
wire n_9482;
wire n_3629;
wire n_969;
wire n_8877;
wire n_9412;
wire n_15561;
wire n_6321;
wire n_6819;
wire n_10136;
wire n_15148;
wire n_16457;
wire n_19560;
wire n_11356;
wire n_1379;
wire n_15955;
wire n_214;
wire n_8688;
wire n_4910;
wire n_3083;
wire n_10692;
wire n_14826;
wire n_16421;
wire n_15776;
wire n_11280;
wire n_14987;
wire n_8686;
wire n_12239;
wire n_17641;
wire n_3830;
wire n_8403;
wire n_11493;
wire n_17742;
wire n_3117;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_5623;
wire n_15269;
wire n_10471;
wire n_2385;
wire n_4112;
wire n_3739;
wire n_14946;
wire n_18727;
wire n_15674;
wire n_4352;
wire n_17933;
wire n_8780;
wire n_17384;
wire n_7958;
wire n_18037;
wire n_4980;
wire n_11885;
wire n_1924;
wire n_15855;
wire n_3363;
wire n_10777;
wire n_3721;
wire n_16490;
wire n_7760;
wire n_13306;
wire n_9753;
wire n_8722;
wire n_16489;
wire n_19580;
wire n_8589;
wire n_3969;
wire n_7573;
wire n_6281;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_4256;
wire n_4938;
wire n_8608;
wire n_12874;
wire n_11480;
wire n_11194;
wire n_10469;
wire n_445;
wire n_18650;
wire n_930;
wire n_9342;
wire n_18062;
wire n_2620;
wire n_9329;
wire n_1945;
wire n_5426;
wire n_19257;
wire n_17119;
wire n_9868;
wire n_1414;
wire n_7048;
wire n_944;
wire n_16491;
wire n_2744;
wire n_1011;
wire n_1566;
wire n_8145;
wire n_8928;
wire n_17638;
wire n_7682;
wire n_990;
wire n_18584;
wire n_6231;
wire n_12509;
wire n_14902;
wire n_6932;
wire n_13527;
wire n_7901;
wire n_870;
wire n_366;
wire n_5709;
wire n_7658;
wire n_10979;
wire n_10055;
wire n_19753;
wire n_19765;
wire n_3802;
wire n_6996;
wire n_15935;
wire n_17674;
wire n_376;
wire n_2111;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_17182;
wire n_6337;
wire n_18212;
wire n_3643;
wire n_2425;
wire n_12936;
wire n_8227;
wire n_18424;
wire n_3060;
wire n_10482;
wire n_4105;
wire n_7405;
wire n_14151;
wire n_4926;
wire n_1518;
wire n_8314;
wire n_9386;
wire n_15120;
wire n_11121;
wire n_3038;
wire n_11270;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_10321;
wire n_5310;
wire n_9661;
wire n_14284;
wire n_3863;
wire n_5722;
wire n_4640;
wire n_13232;
wire n_13001;
wire n_17377;
wire n_9901;
wire n_17334;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_4628;
wire n_8407;
wire n_8567;
wire n_15455;
wire n_11288;
wire n_12772;
wire n_5237;
wire n_409;
wire n_11042;
wire n_10726;
wire n_16534;
wire n_19304;
wire n_4460;
wire n_4108;
wire n_14681;
wire n_11272;
wire n_14230;
wire n_5853;
wire n_8283;
wire n_5011;
wire n_14546;
wire n_9882;
wire n_16484;
wire n_10637;
wire n_9205;
wire n_17464;
wire n_7972;
wire n_1675;
wire n_13512;
wire n_7916;
wire n_9368;
wire n_13069;
wire n_12362;
wire n_19038;
wire n_6167;
wire n_13233;
wire n_18495;
wire n_8008;
wire n_18833;
wire n_13297;
wire n_2553;
wire n_6307;
wire n_149;
wire n_632;
wire n_2038;
wire n_7483;
wire n_14873;
wire n_9504;
wire n_14840;
wire n_16556;
wire n_6267;
wire n_5998;
wire n_17861;
wire n_6568;
wire n_19083;
wire n_7507;
wire n_7159;
wire n_18038;
wire n_6028;
wire n_1417;
wire n_16072;
wire n_14083;
wire n_681;
wire n_10189;
wire n_8697;
wire n_6813;
wire n_6669;
wire n_422;
wire n_8420;
wire n_8297;
wire n_3079;
wire n_10881;
wire n_13519;
wire n_16583;
wire n_15641;
wire n_16007;
wire n_17129;
wire n_4853;
wire n_8639;
wire n_16796;
wire n_16510;
wire n_531;
wire n_15892;
wire n_4272;
wire n_14049;
wire n_1025;
wire n_7562;
wire n_3111;
wire n_336;
wire n_12019;
wire n_8176;
wire n_14529;
wire n_17624;
wire n_16106;
wire n_10891;
wire n_9026;
wire n_10803;
wire n_13190;
wire n_6188;
wire n_5262;
wire n_4670;
wire n_4882;
wire n_11695;
wire n_17595;
wire n_4738;
wire n_8113;
wire n_18922;
wire n_15877;
wire n_1307;
wire n_11453;
wire n_19233;
wire n_17896;
wire n_19088;
wire n_5713;
wire n_16445;
wire n_168;
wire n_6318;
wire n_2353;
wire n_16997;
wire n_4099;
wire n_14690;
wire n_19252;
wire n_17356;
wire n_1738;
wire n_10290;
wire n_19705;
wire n_11862;
wire n_14839;
wire n_15409;
wire n_16207;
wire n_9433;
wire n_18568;
wire n_11660;
wire n_14249;
wire n_14241;
wire n_6604;
wire n_2386;
wire n_5373;
wire n_1724;
wire n_16101;
wire n_3708;
wire n_6391;
wire n_10284;
wire n_14446;
wire n_14719;
wire n_15575;
wire n_12971;
wire n_8522;
wire n_7942;
wire n_16599;
wire n_6473;
wire n_18620;
wire n_15696;
wire n_14558;
wire n_19695;
wire n_11318;
wire n_17198;
wire n_7725;
wire n_16950;
wire n_8626;
wire n_1393;
wire n_1867;
wire n_1603;
wire n_19277;
wire n_5466;
wire n_19475;
wire n_15095;
wire n_5955;
wire n_658;
wire n_1874;
wire n_11487;
wire n_2825;
wire n_8441;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_7778;
wire n_758;
wire n_2256;
wire n_4060;
wire n_8397;
wire n_5796;
wire n_17916;
wire n_8726;
wire n_17250;
wire n_770;
wire n_6958;
wire n_15417;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_14713;
wire n_4687;
wire n_7531;
wire n_18686;
wire n_1404;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_14202;
wire n_15859;
wire n_11933;
wire n_14554;
wire n_9887;
wire n_4600;
wire n_13211;
wire n_8316;
wire n_5829;
wire n_19654;
wire n_8057;
wire n_5191;
wire n_1231;
wire n_14874;
wire n_18198;
wire n_2370;
wire n_18550;
wire n_4253;
wire n_407;
wire n_913;
wire n_16824;
wire n_15098;
wire n_867;
wire n_16832;
wire n_13336;
wire n_1333;
wire n_2496;
wire n_16074;
wire n_3189;
wire n_19487;
wire n_18664;
wire n_13102;
wire n_4691;
wire n_12894;
wire n_10492;
wire n_15769;
wire n_4297;
wire n_9247;
wire n_17340;
wire n_8378;
wire n_2907;
wire n_577;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_9570;
wire n_5675;
wire n_12356;
wire n_2778;
wire n_19454;
wire n_11077;
wire n_1909;
wire n_5020;
wire n_9846;
wire n_13262;
wire n_1123;
wire n_10764;
wire n_18005;
wire n_18429;
wire n_9677;
wire n_3934;
wire n_4033;
wire n_6804;
wire n_6603;
wire n_17812;
wire n_3193;
wire n_7534;
wire n_8201;
wire n_4354;
wire n_16485;
wire n_9348;
wire n_14262;
wire n_1530;
wire n_8696;
wire n_938;
wire n_6396;
wire n_12630;
wire n_6890;
wire n_549;
wire n_4377;
wire n_12022;
wire n_905;
wire n_10741;
wire n_6109;
wire n_14727;
wire n_12425;
wire n_14762;
wire n_322;
wire n_689;
wire n_13507;
wire n_10915;
wire n_18290;
wire n_558;
wire n_3036;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_17133;
wire n_17729;
wire n_15410;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_16002;
wire n_16258;
wire n_13594;
wire n_10680;
wire n_3599;
wire n_5543;
wire n_5885;
wire n_14228;
wire n_5356;
wire n_3772;
wire n_5458;
wire n_16131;
wire n_11473;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_11726;
wire n_15944;
wire n_12574;
wire n_8833;
wire n_10142;
wire n_7828;
wire n_9918;
wire n_18643;
wire n_15932;
wire n_16345;
wire n_4427;
wire n_9390;
wire n_10069;
wire n_17325;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_18233;
wire n_5510;
wire n_5555;
wire n_13678;
wire n_12458;
wire n_19291;
wire n_6066;
wire n_14582;
wire n_6897;
wire n_13523;
wire n_9619;
wire n_15117;
wire n_11171;
wire n_4886;
wire n_9187;
wire n_2733;
wire n_16621;
wire n_13819;
wire n_15777;
wire n_14424;
wire n_18398;
wire n_14523;
wire n_11063;
wire n_18846;
wire n_9989;
wire n_8319;
wire n_4200;
wire n_3460;
wire n_12853;
wire n_12942;
wire n_9259;
wire n_3519;
wire n_12397;
wire n_16555;
wire n_15336;
wire n_14161;
wire n_6573;
wire n_16760;
wire n_7634;
wire n_5078;
wire n_13290;
wire n_13500;
wire n_11440;
wire n_16844;
wire n_10483;
wire n_17758;
wire n_4737;
wire n_4116;
wire n_7285;
wire n_11337;
wire n_12005;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_18610;
wire n_9824;
wire n_342;
wire n_15089;
wire n_2658;
wire n_2665;
wire n_8233;
wire n_6130;
wire n_7273;
wire n_14750;
wire n_17939;
wire n_5976;
wire n_14074;
wire n_840;
wire n_2913;
wire n_12800;
wire n_2230;
wire n_1969;
wire n_1565;
wire n_16574;
wire n_15145;
wire n_17516;
wire n_8187;
wire n_9399;
wire n_15838;
wire n_15297;
wire n_13979;
wire n_9740;
wire n_615;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_17178;
wire n_9764;
wire n_4854;
wire n_15160;
wire n_3789;
wire n_605;
wire n_12354;
wire n_7597;
wire n_12666;
wire n_14297;
wire n_17388;
wire n_16368;
wire n_12631;
wire n_1646;
wire n_19154;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_18426;
wire n_18073;
wire n_6921;
wire n_14675;
wire n_18905;
wire n_9826;
wire n_3171;
wire n_3608;
wire n_11942;
wire n_15998;
wire n_3459;
wire n_19138;
wire n_6624;
wire n_6956;
wire n_12966;
wire n_15851;
wire n_15884;
wire n_5656;
wire n_5125;
wire n_7329;
wire n_14502;
wire n_14533;
wire n_5652;
wire n_17935;
wire n_10752;
wire n_18630;
wire n_10067;
wire n_18021;
wire n_10399;
wire n_12498;
wire n_656;
wire n_11010;
wire n_9590;
wire n_16017;
wire n_2717;
wire n_11588;
wire n_16346;
wire n_738;
wire n_13956;
wire n_3497;
wire n_7418;
wire n_6880;
wire n_19305;
wire n_3580;
wire n_12387;
wire n_19783;
wire n_9497;
wire n_13255;
wire n_15911;
wire n_2307;
wire n_3704;
wire n_684;
wire n_9219;
wire n_17376;
wire n_8028;
wire n_4280;
wire n_8914;
wire n_1181;
wire n_15276;
wire n_8391;
wire n_16343;
wire n_13749;
wire n_15552;
wire n_17722;
wire n_19370;
wire n_16228;
wire n_803;
wire n_1817;
wire n_12862;
wire n_13621;
wire n_8216;
wire n_2868;
wire n_16953;
wire n_2231;
wire n_3609;
wire n_9982;
wire n_7804;
wire n_18948;
wire n_12656;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_19150;
wire n_8263;
wire n_6438;
wire n_11936;
wire n_19132;
wire n_10374;
wire n_7332;
wire n_10382;
wire n_18247;
wire n_4455;
wire n_8374;
wire n_13223;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_18909;
wire n_13728;
wire n_4806;
wire n_7386;
wire n_17824;
wire n_11018;
wire n_10981;
wire n_16014;
wire n_2682;
wire n_13379;
wire n_13781;
wire n_19311;
wire n_5098;
wire n_17513;
wire n_10344;
wire n_5707;
wire n_14613;
wire n_19451;
wire n_11515;
wire n_17466;
wire n_3505;
wire n_15881;
wire n_7637;
wire n_16577;
wire n_10318;
wire n_4796;
wire n_4442;
wire n_18422;
wire n_2581;
wire n_18091;
wire n_12890;
wire n_3590;
wire n_5344;
wire n_954;
wire n_13994;
wire n_4419;
wire n_17060;
wire n_11972;
wire n_13484;
wire n_17298;
wire n_8460;
wire n_3327;
wire n_17468;
wire n_14593;
wire n_2701;
wire n_16013;
wire n_1080;
wire n_7409;
wire n_19266;
wire n_10735;
wire n_17153;
wire n_13807;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_16942;
wire n_2421;
wire n_17569;
wire n_4387;
wire n_2618;
wire n_2464;
wire n_5128;
wire n_18661;
wire n_14033;
wire n_2224;
wire n_10393;
wire n_1092;
wire n_15221;
wire n_5467;
wire n_16090;
wire n_18467;
wire n_4890;
wire n_1784;
wire n_9045;
wire n_12281;
wire n_9373;
wire n_14337;
wire n_2929;
wire n_11809;
wire n_17994;
wire n_9967;
wire n_13553;
wire n_4236;
wire n_7187;
wire n_19039;
wire n_17063;
wire n_19692;
wire n_1831;
wire n_9182;
wire n_5079;
wire n_9365;
wire n_18960;
wire n_10909;
wire n_10083;
wire n_6336;
wire n_18891;
wire n_9224;
wire n_10347;
wire n_6541;
wire n_12410;
wire n_4706;
wire n_16327;
wire n_19238;
wire n_14707;
wire n_16043;
wire n_19677;
wire n_4622;
wire n_14612;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_2732;
wire n_17688;
wire n_4206;
wire n_2249;
wire n_18794;
wire n_5835;
wire n_7979;
wire n_13382;
wire n_11675;
wire n_15543;
wire n_15906;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_2955;
wire n_11083;
wire n_17418;
wire n_2158;
wire n_7866;
wire n_3367;
wire n_7205;
wire n_18283;
wire n_2202;
wire n_736;
wire n_11728;
wire n_2993;
wire n_4754;
wire n_11698;
wire n_4647;
wire n_9556;
wire n_8590;
wire n_16682;
wire n_4030;
wire n_1995;
wire n_17038;
wire n_15798;
wire n_4760;
wire n_11326;
wire n_6421;
wire n_19743;
wire n_11870;
wire n_7407;
wire n_6328;
wire n_11283;
wire n_6236;
wire n_11834;
wire n_13361;
wire n_17286;
wire n_4509;
wire n_15061;
wire n_2875;
wire n_1103;
wire n_6144;
wire n_11506;
wire n_13161;
wire n_10135;
wire n_144;
wire n_2219;
wire n_14010;
wire n_16413;
wire n_999;
wire n_4897;
wire n_19796;
wire n_15030;
wire n_18205;
wire n_9152;
wire n_3539;
wire n_16451;
wire n_19590;
wire n_8364;
wire n_3276;
wire n_15228;
wire n_15832;
wire n_10720;
wire n_10535;
wire n_19349;
wire n_17629;
wire n_17536;
wire n_3886;
wire n_6708;
wire n_11236;
wire n_18793;
wire n_4420;
wire n_892;
wire n_18529;
wire n_6242;
wire n_12379;
wire n_1468;
wire n_2855;
wire n_2156;
wire n_18222;
wire n_12932;
wire n_14078;
wire n_3548;
wire n_18985;
wire n_8548;
wire n_19793;
wire n_10672;
wire n_7645;
wire n_14222;
wire n_16990;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_12114;
wire n_10308;
wire n_11608;
wire n_14430;
wire n_1015;
wire n_10623;
wire n_4797;
wire n_6285;
wire n_4270;
wire n_16545;
wire n_19339;
wire n_13709;
wire n_4945;
wire n_17713;
wire n_5677;
wire n_9454;
wire n_10586;
wire n_8742;
wire n_12626;
wire n_11967;
wire n_9253;
wire n_15084;
wire n_13559;
wire n_8874;
wire n_5927;
wire n_15071;
wire n_11996;
wire n_9566;
wire n_11338;
wire n_13426;
wire n_1356;
wire n_4333;
wire n_18826;
wire n_7666;
wire n_11250;
wire n_15328;
wire n_1452;
wire n_2854;
wire n_7963;
wire n_6398;
wire n_8329;
wire n_302;
wire n_9503;
wire n_8270;
wire n_16051;
wire n_11738;
wire n_18196;
wire n_3217;
wire n_1983;
wire n_11522;
wire n_7737;
wire n_16569;
wire n_8614;
wire n_18459;
wire n_9568;
wire n_15621;
wire n_18411;
wire n_8816;
wire n_9119;
wire n_19337;
wire n_13529;
wire n_6224;
wire n_3279;
wire n_18293;
wire n_2402;
wire n_1081;
wire n_19616;
wire n_1084;
wire n_6614;
wire n_5912;
wire n_18395;
wire n_3501;
wire n_374;
wire n_12554;
wire n_8035;
wire n_12722;
wire n_6735;
wire n_17445;
wire n_10491;
wire n_921;
wire n_12037;
wire n_15371;
wire n_17572;
wire n_13453;
wire n_15080;
wire n_5265;
wire n_2257;
wire n_9943;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_7152;
wire n_2200;
wire n_9575;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_10521;
wire n_9610;
wire n_16483;
wire n_14016;
wire n_12323;
wire n_15566;
wire n_10527;
wire n_3115;
wire n_7570;
wire n_2084;
wire n_4875;
wire n_7817;
wire n_5682;
wire n_5387;
wire n_654;
wire n_11394;
wire n_2458;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_13897;
wire n_2527;
wire n_14792;
wire n_16290;
wire n_14248;
wire n_8370;
wire n_164;
wire n_13300;
wire n_16296;
wire n_5681;
wire n_7566;
wire n_11940;
wire n_1271;
wire n_4901;
wire n_9217;
wire n_12901;
wire n_4040;
wire n_10518;
wire n_2406;
wire n_7617;
wire n_15170;
wire n_16936;
wire n_19262;
wire n_9771;
wire n_15774;
wire n_5316;
wire n_7718;
wire n_244;
wire n_13844;
wire n_19246;
wire n_7396;
wire n_282;
wire n_18543;
wire n_5703;
wire n_18930;
wire n_833;
wire n_523;
wire n_7998;
wire n_12432;
wire n_7561;
wire n_18349;
wire n_6810;
wire n_2196;
wire n_17010;
wire n_17040;
wire n_16130;
wire n_12879;
wire n_5564;
wire n_13746;
wire n_12559;
wire n_13508;
wire n_14660;
wire n_4530;
wire n_9899;
wire n_13004;
wire n_5406;
wire n_13479;
wire n_8277;
wire n_652;
wire n_18014;
wire n_1906;
wire n_14437;
wire n_4841;
wire n_1758;
wire n_13759;
wire n_5806;
wire n_4338;
wire n_10486;
wire n_306;
wire n_16613;
wire n_8724;
wire n_5738;
wire n_15938;
wire n_17216;
wire n_3151;
wire n_15146;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_9995;
wire n_5710;
wire n_9076;
wire n_12351;
wire n_16360;
wire n_19146;
wire n_13359;
wire n_10372;
wire n_3558;
wire n_14867;
wire n_1984;
wire n_2236;
wire n_6044;
wire n_9491;
wire n_8867;
wire n_4326;
wire n_12702;
wire n_17811;
wire n_15188;
wire n_2834;
wire n_12439;
wire n_19478;
wire n_11008;
wire n_6125;
wire n_7314;
wire n_786;
wire n_14186;
wire n_7526;
wire n_17816;
wire n_5040;
wire n_14023;
wire n_19758;
wire n_17890;
wire n_10736;
wire n_19550;
wire n_11575;
wire n_7004;
wire n_14418;
wire n_8308;
wire n_18897;
wire n_151;
wire n_8165;
wire n_14283;
wire n_4788;
wire n_8400;
wire n_18177;
wire n_5977;
wire n_10446;
wire n_7879;
wire n_16372;
wire n_1908;
wire n_15958;
wire n_18853;
wire n_7696;
wire n_11570;
wire n_16567;
wire n_12952;
wire n_19096;
wire n_2045;
wire n_14795;
wire n_3687;
wire n_2216;
wire n_19318;
wire n_3621;
wire n_16425;
wire n_16769;
wire n_10603;
wire n_12004;
wire n_6962;
wire n_8217;
wire n_12830;
wire n_8858;
wire n_7246;
wire n_10255;
wire n_2719;
wire n_11490;
wire n_8689;
wire n_10113;
wire n_15086;
wire n_680;
wire n_3339;
wire n_10188;
wire n_6853;
wire n_10686;
wire n_9841;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_16838;
wire n_10974;
wire n_11067;
wire n_8627;
wire n_13659;
wire n_12034;
wire n_16586;
wire n_1399;
wire n_16056;
wire n_13303;
wire n_6894;
wire n_13346;
wire n_13702;
wire n_9179;
wire n_2358;
wire n_15894;
wire n_8752;
wire n_2186;
wire n_18237;
wire n_3034;
wire n_4408;
wire n_18367;
wire n_10937;
wire n_643;
wire n_12134;
wire n_400;
wire n_12449;
wire n_2814;
wire n_16399;
wire n_789;
wire n_327;
wire n_6284;
wire n_10167;
wire n_12524;
wire n_18113;
wire n_6883;
wire n_12963;
wire n_10428;
wire n_16860;
wire n_17869;
wire n_19199;
wire n_18682;
wire n_12366;
wire n_747;
wire n_14951;
wire n_11068;
wire n_11035;
wire n_5495;
wire n_535;
wire n_19148;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_9420;
wire n_3851;
wire n_16995;
wire n_14336;
wire n_7825;
wire n_10079;
wire n_7212;
wire n_19436;
wire n_6966;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_6035;
wire n_1652;
wire n_15435;
wire n_8634;
wire n_9531;
wire n_12605;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_2914;
wire n_12828;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_8532;
wire n_19109;
wire n_12661;
wire n_10588;
wire n_8991;
wire n_8065;
wire n_3100;
wire n_11140;
wire n_3573;
wire n_17882;
wire n_17677;
wire n_8518;
wire n_197;
wire n_18226;
wire n_13017;
wire n_1083;
wire n_16884;
wire n_15199;
wire n_18153;
wire n_1721;
wire n_9812;
wire n_1737;
wire n_15419;
wire n_752;
wire n_7361;
wire n_9949;
wire n_1028;
wire n_14889;
wire n_7228;
wire n_9576;
wire n_5872;
wire n_1973;
wire n_3181;
wire n_6338;
wire n_15267;
wire n_19366;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_6266;
wire n_14796;
wire n_2242;
wire n_19125;
wire n_11364;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_19069;
wire n_17397;
wire n_7018;
wire n_5873;
wire n_7975;
wire n_10009;
wire n_9279;
wire n_11902;
wire n_924;
wire n_16782;
wire n_11993;
wire n_2318;
wire n_10443;
wire n_3170;
wire n_17317;
wire n_12813;
wire n_13534;
wire n_3304;
wire n_4968;
wire n_10384;
wire n_5085;
wire n_5736;
wire n_2433;
wire n_829;
wire n_7978;
wire n_10293;
wire n_17422;
wire n_12312;
wire n_10074;
wire n_13097;
wire n_17850;
wire n_15786;
wire n_4208;
wire n_9632;
wire n_12256;
wire n_11812;
wire n_9711;
wire n_9431;
wire n_4779;
wire n_14650;
wire n_18068;
wire n_481;
wire n_14610;
wire n_997;
wire n_11505;
wire n_4437;
wire n_7316;
wire n_17938;
wire n_1306;
wire n_3264;
wire n_18955;
wire n_7103;
wire n_14601;
wire n_436;
wire n_11363;
wire n_15794;
wire n_17066;
wire n_2426;
wire n_2478;
wire n_14645;
wire n_1133;
wire n_4642;
wire n_11151;
wire n_15825;
wire n_10716;
wire n_10664;
wire n_2578;
wire n_3709;
wire n_11434;
wire n_3738;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_5812;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_19536;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_8788;
wire n_10992;
wire n_19380;
wire n_1629;
wire n_10160;
wire n_10560;
wire n_7404;
wire n_12857;
wire n_13171;
wire n_18615;
wire n_1260;
wire n_309;
wire n_9854;
wire n_14854;
wire n_812;
wire n_15266;
wire n_1006;
wire n_7271;
wire n_9713;
wire n_16501;
wire n_257;
wire n_19264;
wire n_1311;
wire n_10300;
wire n_9588;
wire n_14218;
wire n_15107;
wire n_6842;
wire n_13876;
wire n_4803;
wire n_18935;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_14487;
wire n_9127;
wire n_5996;
wire n_16767;
wire n_9869;
wire n_315;
wire n_14449;
wire n_17094;
wire n_12885;
wire n_2579;
wire n_15539;
wire n_2105;
wire n_135;
wire n_9715;
wire n_17112;
wire n_8618;
wire n_18916;
wire n_3387;
wire n_12108;
wire n_7535;
wire n_11531;
wire n_19450;
wire n_9407;
wire n_2912;
wire n_14476;
wire n_3409;
wire n_15244;
wire n_2320;
wire n_19574;
wire n_11824;
wire n_1259;
wire n_6957;
wire n_9361;
wire n_13976;
wire n_16578;
wire n_18949;
wire n_13579;
wire n_11566;
wire n_17452;
wire n_16650;
wire n_14639;
wire n_8990;
wire n_17067;
wire n_6444;
wire n_19170;
wire n_226;
wire n_7944;
wire n_19235;
wire n_11374;
wire n_8647;
wire n_15857;
wire n_2003;
wire n_7016;
wire n_10782;
wire n_13557;
wire n_3301;
wire n_16709;
wire n_6379;
wire n_15589;
wire n_17491;
wire n_2324;
wire n_17757;
wire n_12754;
wire n_245;
wire n_13583;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_17333;
wire n_19043;
wire n_2847;
wire n_17749;
wire n_16658;
wire n_4050;
wire n_13455;
wire n_883;
wire n_19136;
wire n_6232;
wire n_9132;
wire n_1032;
wire n_10861;
wire n_17035;
wire n_8879;
wire n_1099;
wire n_19639;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_2211;
wire n_6362;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_9332;
wire n_17097;
wire n_369;
wire n_16765;
wire n_11030;
wire n_4179;
wire n_1285;
wire n_6326;
wire n_10073;
wire n_14619;
wire n_1590;
wire n_5072;
wire n_7241;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_15427;
wire n_17364;
wire n_10333;
wire n_12430;
wire n_18330;
wire n_7235;
wire n_6239;
wire n_2340;
wire n_13407;
wire n_5896;
wire n_13676;
wire n_18391;
wire n_16694;
wire n_12557;
wire n_13788;
wire n_6974;
wire n_16537;
wire n_18227;
wire n_18666;
wire n_8939;
wire n_13584;
wire n_428;
wire n_15471;
wire n_12139;
wire n_9030;
wire n_7657;
wire n_822;
wire n_2791;
wire n_19433;
wire n_9665;
wire n_5044;
wire n_5134;
wire n_7096;
wire n_3063;
wire n_13327;
wire n_1550;
wire n_19098;
wire n_11197;
wire n_491;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_10093;
wire n_15428;
wire n_15014;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_7999;
wire n_10675;
wire n_6087;
wire n_16311;
wire n_538;
wire n_4164;
wire n_10107;
wire n_3225;
wire n_15536;
wire n_13224;
wire n_11469;
wire n_5022;
wire n_14046;
wire n_7041;
wire n_10742;
wire n_10829;
wire n_19115;
wire n_12389;
wire n_9309;
wire n_19632;
wire n_10620;
wire n_13971;
wire n_16750;
wire n_7672;
wire n_2551;
wire n_5047;
wire n_7318;
wire n_19325;
wire n_12995;
wire n_18261;
wire n_14406;
wire n_13209;
wire n_11883;
wire n_14959;
wire n_3269;
wire n_15387;
wire n_11901;
wire n_6352;
wire n_15973;
wire n_8542;
wire n_19747;
wire n_10859;
wire n_18446;
wire n_8576;
wire n_14807;
wire n_8038;
wire n_11572;
wire n_5141;
wire n_3603;
wire n_14493;
wire n_18306;
wire n_13113;
wire n_13387;
wire n_8716;
wire n_3822;
wire n_5535;
wire n_19411;
wire n_3812;
wire n_16807;
wire n_18538;
wire n_2696;
wire n_17576;
wire n_4080;
wire n_6002;
wire n_541;
wire n_18665;
wire n_15538;
wire n_2073;
wire n_2273;
wire n_4941;
wire n_5506;
wire n_11399;
wire n_17578;
wire n_8768;
wire n_10884;
wire n_1162;
wire n_15870;
wire n_12035;
wire n_13006;
wire n_12791;
wire n_7600;
wire n_14742;
wire n_2831;
wire n_4158;
wire n_6644;
wire n_17878;
wire n_4795;
wire n_19528;
wire n_12810;
wire n_16930;
wire n_3824;
wire n_13947;
wire n_11322;
wire n_17562;
wire n_4544;
wire n_5841;
wire n_12241;
wire n_9343;
wire n_15895;
wire n_16554;
wire n_17779;
wire n_5108;
wire n_7347;
wire n_11057;
wire n_2355;
wire n_10969;
wire n_14474;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_8863;
wire n_18501;
wire n_7759;
wire n_11551;
wire n_18049;
wire n_7479;
wire n_2866;
wire n_10598;
wire n_8947;
wire n_15494;
wire n_10717;
wire n_11118;
wire n_18579;
wire n_3649;
wire n_2821;
wire n_6067;
wire n_12674;
wire n_17727;
wire n_17839;
wire n_8510;
wire n_12230;
wire n_11410;
wire n_19282;
wire n_1563;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_17122;
wire n_1359;
wire n_5367;
wire n_16778;
wire n_3794;
wire n_12220;
wire n_6868;
wire n_1335;
wire n_5970;
wire n_16133;
wire n_12283;
wire n_7174;
wire n_9421;
wire n_5202;
wire n_19055;
wire n_13383;
wire n_18787;
wire n_17079;
wire n_8021;
wire n_3346;
wire n_7803;
wire n_15124;
wire n_12595;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_13983;
wire n_9416;
wire n_6225;
wire n_5502;
wire n_3428;
wire n_4552;
wire n_6218;
wire n_17489;
wire n_12920;
wire n_13317;
wire n_9929;
wire n_2519;
wire n_9953;
wire n_1063;
wire n_6648;
wire n_15578;
wire n_10955;
wire n_7927;
wire n_11011;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_12141;
wire n_9346;
wire n_7920;
wire n_437;
wire n_12774;
wire n_4169;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_697;
wire n_17399;
wire n_388;
wire n_7025;
wire n_15886;
wire n_17022;
wire n_15856;
wire n_1757;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_14357;
wire n_13044;
wire n_13228;
wire n_13518;
wire n_4070;
wire n_19763;
wire n_3885;
wire n_1369;
wire n_14008;
wire n_17069;
wire n_12746;
wire n_4031;
wire n_16162;
wire n_10970;
wire n_16285;
wire n_14927;
wire n_13881;
wire n_3209;
wire n_17205;
wire n_5547;
wire n_13747;
wire n_1391;
wire n_12532;
wire n_10238;
wire n_8931;
wire n_5596;
wire n_4653;
wire n_4435;
wire n_8334;
wire n_4019;
wire n_1071;
wire n_11681;
wire n_10890;
wire n_11202;
wire n_19513;
wire n_10552;
wire n_5815;
wire n_15254;
wire n_6595;
wire n_8539;
wire n_10205;
wire n_16947;
wire n_15747;
wire n_3727;
wire n_13899;
wire n_6306;
wire n_19386;
wire n_1714;
wire n_16235;
wire n_11663;
wire n_542;
wire n_11331;
wire n_305;
wire n_19472;
wire n_9528;
wire n_14348;
wire n_7583;
wire n_12201;
wire n_19334;
wire n_14086;
wire n_12499;
wire n_19173;
wire n_12448;
wire n_10610;
wire n_12761;
wire n_11187;
wire n_16455;
wire n_15004;
wire n_16625;
wire n_16025;
wire n_5520;
wire n_2638;
wire n_14552;
wire n_7353;
wire n_9490;
wire n_19767;
wire n_5669;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_145;
wire n_4775;
wire n_16249;
wire n_16435;
wire n_4674;
wire n_16723;
wire n_11446;
wire n_10910;
wire n_294;
wire n_8242;
wire n_11540;
wire n_13248;
wire n_17296;
wire n_19237;
wire n_9819;
wire n_15338;
wire n_8184;
wire n_425;
wire n_6525;
wire n_4286;
wire n_13119;
wire n_2958;
wire n_12642;
wire n_3731;
wire n_1822;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_2489;
wire n_17361;
wire n_16080;
wire n_4525;
wire n_9992;
wire n_15180;
wire n_15692;
wire n_5712;
wire n_12669;
wire n_14296;
wire n_6702;
wire n_19490;
wire n_11179;
wire n_17074;
wire n_2520;
wire n_446;
wire n_7749;
wire n_10078;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_18496;
wire n_8705;
wire n_19107;
wire n_11779;
wire n_7508;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_14211;
wire n_7574;
wire n_4306;
wire n_13516;
wire n_14273;
wire n_12462;
wire n_4453;
wire n_16462;
wire n_18648;
wire n_4005;
wire n_6169;
wire n_18775;
wire n_15230;
wire n_3546;
wire n_3661;
wire n_12735;
wire n_10709;
wire n_12646;
wire n_15875;
wire n_7352;
wire n_10244;
wire n_755;
wire n_18512;
wire n_12999;
wire n_12682;
wire n_14802;
wire n_6848;
wire n_17415;
wire n_3509;
wire n_10043;
wire n_14834;
wire n_5919;
wire n_8159;
wire n_14346;
wire n_16955;
wire n_7439;
wire n_17653;
wire n_2504;
wire n_14506;
wire n_2623;
wire n_18822;
wire n_16018;
wire n_14615;
wire n_15222;
wire n_6850;
wire n_18991;
wire n_15285;
wire n_5005;
wire n_13294;
wire n_6098;
wire n_7112;
wire n_11307;
wire n_19021;
wire n_17860;
wire n_18274;
wire n_9545;
wire n_596;
wire n_9629;
wire n_9603;
wire n_18003;
wire n_12719;
wire n_10342;
wire n_15361;
wire n_3322;
wire n_19037;
wire n_16244;
wire n_17862;
wire n_4654;
wire n_13438;
wire n_3640;
wire n_1159;
wire n_995;
wire n_15850;
wire n_9930;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_14988;
wire n_9659;
wire n_3226;
wire n_2780;
wire n_16293;
wire n_9897;
wire n_9241;
wire n_14590;
wire n_14603;
wire n_8185;
wire n_11466;
wire n_5061;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_9291;
wire n_4063;
wire n_11982;
wire n_2601;
wire n_773;
wire n_11873;
wire n_15821;
wire n_920;
wire n_10185;
wire n_11182;
wire n_3212;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_18807;
wire n_4721;
wire n_14145;
wire n_11991;
wire n_848;
wire n_12875;
wire n_15064;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_13918;
wire n_13775;
wire n_9851;
wire n_11799;
wire n_8009;
wire n_7852;
wire n_1881;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_18307;
wire n_2720;
wire n_18110;
wire n_14973;
wire n_16751;
wire n_7220;
wire n_18015;
wire n_1323;
wire n_2627;
wire n_18242;
wire n_6550;
wire n_3004;
wire n_8841;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_15136;
wire n_1764;
wire n_10354;
wire n_7465;
wire n_13177;
wire n_4546;
wire n_12724;
wire n_14958;
wire n_6672;
wire n_16744;
wire n_17876;
wire n_1551;
wire n_15992;
wire n_7738;
wire n_17406;
wire n_19079;
wire n_8395;
wire n_6634;
wire n_14758;
wire n_18392;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_16802;
wire n_17909;
wire n_18439;
wire n_5735;
wire n_19022;
wire n_13311;
wire n_19700;
wire n_2278;
wire n_16020;
wire n_11513;
wire n_7464;
wire n_8937;
wire n_7115;
wire n_2924;
wire n_12087;
wire n_13675;
wire n_15022;
wire n_18693;
wire n_3595;
wire n_6104;
wire n_10537;
wire n_421;
wire n_6082;
wire n_18305;
wire n_1270;
wire n_10426;
wire n_1852;
wire n_9167;
wire n_12082;
wire n_9655;
wire n_11436;
wire n_11729;
wire n_3230;
wire n_19276;
wire n_1499;
wire n_12989;
wire n_504;
wire n_5877;
wire n_8845;
wire n_15198;
wire n_6018;
wire n_17902;
wire n_13620;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_17144;
wire n_12464;
wire n_9560;
wire n_18362;
wire n_18886;
wire n_1182;
wire n_15007;
wire n_15197;
wire n_167;
wire n_8519;
wire n_5582;
wire n_5886;
wire n_1216;
wire n_6032;
wire n_18982;
wire n_9319;
wire n_5446;
wire n_3010;
wire n_12450;
wire n_5224;
wire n_19776;
wire n_14648;
wire n_11767;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_9401;
wire n_11586;
wire n_12149;
wire n_12002;
wire n_12836;
wire n_19506;
wire n_17084;
wire n_13548;
wire n_15710;
wire n_2232;
wire n_11195;
wire n_4038;
wire n_16240;
wire n_2790;
wire n_9747;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_17190;
wire n_3784;
wire n_17973;
wire n_220;
wire n_8586;
wire n_9058;
wire n_18707;
wire n_1472;
wire n_18547;
wire n_16700;
wire n_5454;
wire n_800;
wire n_10780;
wire n_17940;
wire n_8756;
wire n_1840;
wire n_4434;
wire n_13406;
wire n_16371;
wire n_7923;
wire n_14040;
wire n_14054;
wire n_8602;
wire n_1346;
wire n_13469;
wire n_10411;
wire n_13249;
wire n_12984;
wire n_18840;
wire n_13587;
wire n_5913;
wire n_10090;
wire n_14872;
wire n_1102;
wire n_8112;
wire n_18959;
wire n_258;
wire n_11567;
wire n_2766;
wire n_19428;
wire n_9292;
wire n_18771;
wire n_12197;
wire n_356;
wire n_17753;
wire n_19134;
wire n_4833;
wire n_11580;
wire n_13326;
wire n_13082;
wire n_6474;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_18518;
wire n_10856;
wire n_12403;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_9584;
wire n_13692;
wire n_8194;
wire n_8055;
wire n_8579;
wire n_10914;
wire n_8360;
wire n_4279;
wire n_6425;
wire n_1456;
wire n_6493;
wire n_14382;
wire n_13396;
wire n_10071;
wire n_8755;
wire n_2099;
wire n_11565;
wire n_3388;
wire n_14911;
wire n_15405;
wire n_5810;
wire n_4461;
wire n_3245;
wire n_4007;
wire n_15643;
wire n_15420;
wire n_13052;
wire n_11013;
wire n_5991;
wire n_1676;
wire n_1319;
wire n_16634;
wire n_16762;
wire n_10035;
wire n_5702;
wire n_18094;
wire n_18673;
wire n_18980;
wire n_14962;
wire n_1633;
wire n_17435;
wire n_8108;
wire n_2820;
wire n_17065;
wire n_12068;
wire n_5250;
wire n_3074;
wire n_17285;
wire n_10041;
wire n_15499;
wire n_5590;
wire n_14514;
wire n_17612;
wire n_8498;
wire n_14256;
wire n_17073;
wire n_16773;
wire n_2727;
wire n_2533;
wire n_5349;
wire n_19320;
wire n_2759;
wire n_2361;
wire n_2266;
wire n_14082;
wire n_7280;
wire n_5833;
wire n_7886;
wire n_15728;
wire n_6884;
wire n_7664;
wire n_18292;
wire n_7012;
wire n_299;
wire n_1248;
wire n_17354;
wire n_12486;
wire n_902;
wire n_2189;
wire n_7376;
wire n_5816;
wire n_15347;
wire n_10137;
wire n_12084;
wire n_16517;
wire n_706;
wire n_1794;
wire n_1236;
wire n_11863;
wire n_17868;
wire n_17033;
wire n_17234;
wire n_430;
wire n_16174;
wire n_18059;
wire n_19015;
wire n_10794;
wire n_14703;
wire n_13533;
wire n_6274;
wire n_8838;
wire n_12109;
wire n_16283;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_2975;
wire n_16088;
wire n_2856;
wire n_4498;
wire n_12320;
wire n_19245;
wire n_9759;
wire n_6992;
wire n_15226;
wire n_19742;
wire n_646;
wire n_528;
wire n_10206;
wire n_1329;
wire n_17736;
wire n_6322;
wire n_5167;
wire n_15425;
wire n_5661;
wire n_16878;
wire n_3589;
wire n_262;
wire n_897;
wire n_7616;
wire n_1800;
wire n_18294;
wire n_9733;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_13011;
wire n_9981;
wire n_18514;
wire n_5558;
wire n_5687;
wire n_16513;
wire n_6378;
wire n_14495;
wire n_1759;
wire n_16879;
wire n_12269;
wire n_853;
wire n_13486;
wire n_11463;
wire n_3585;
wire n_17541;
wire n_5954;
wire n_5025;
wire n_933;
wire n_17394;
wire n_7587;
wire n_3135;
wire n_17496;
wire n_6930;
wire n_17472;
wire n_19121;
wire n_12802;
wire n_11569;
wire n_10064;
wire n_7197;
wire n_9676;
wire n_7393;
wire n_11332;
wire n_13629;
wire n_13207;
wire n_310;
wire n_5766;
wire n_18025;
wire n_7358;
wire n_2796;
wire n_9950;
wire n_18088;
wire n_13589;
wire n_15730;
wire n_18089;
wire n_4534;
wire n_17967;
wire n_19731;
wire n_6929;
wire n_16706;
wire n_11309;
wire n_955;
wire n_8045;
wire n_16032;
wire n_19740;
wire n_19741;
wire n_18910;
wire n_2969;
wire n_2395;
wire n_16959;
wire n_8209;
wire n_14477;
wire n_9213;
wire n_7291;
wire n_14522;
wire n_669;
wire n_16971;
wire n_2290;
wire n_2005;
wire n_13561;
wire n_14720;
wire n_7437;
wire n_16873;
wire n_1408;
wire n_7618;
wire n_8575;
wire n_5733;
wire n_6620;
wire n_6597;
wire n_11105;
wire n_13698;
wire n_13894;
wire n_452;
wire n_6586;
wire n_10474;
wire n_12689;
wire n_18939;
wire n_8789;
wire n_7953;
wire n_19775;
wire n_13540;
wire n_6428;
wire n_5328;
wire n_14642;
wire n_12042;
wire n_14827;
wire n_15481;
wire n_5657;
wire n_174;
wire n_1173;
wire n_13465;
wire n_11130;
wire n_16149;
wire n_11664;
wire n_18705;
wire n_17430;
wire n_15388;
wire n_19242;
wire n_10652;
wire n_13733;
wire n_13098;
wire n_3334;
wire n_9388;
wire n_12654;
wire n_4985;
wire n_10869;
wire n_3823;
wire n_18708;
wire n_19112;
wire n_11783;
wire n_2255;
wire n_17837;
wire n_4678;
wire n_2649;
wire n_9911;
wire n_19603;
wire n_5579;
wire n_414;
wire n_16317;
wire n_1922;
wire n_15187;
wire n_17897;
wire n_12419;
wire n_13763;
wire n_10346;
wire n_4363;
wire n_10473;
wire n_15712;
wire n_5107;
wire n_16985;
wire n_5095;
wire n_8493;
wire n_10957;
wire n_13517;
wire n_11188;
wire n_3404;
wire n_10442;
wire n_1509;
wire n_3290;
wire n_13973;
wire n_7150;
wire n_8252;
wire n_11774;
wire n_3671;
wire n_7015;
wire n_2015;
wire n_3982;
wire n_13206;
wire n_7249;
wire n_1161;
wire n_15939;
wire n_3840;
wire n_3461;
wire n_7985;
wire n_13637;
wire n_3513;
wire n_16705;
wire n_18163;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_15904;
wire n_592;
wire n_12768;
wire n_1156;
wire n_18369;
wire n_16047;
wire n_3508;
wire n_10165;
wire n_8156;
wire n_868;
wire n_19674;
wire n_14923;
wire n_13031;
wire n_19029;
wire n_19316;
wire n_17912;
wire n_13155;
wire n_469;
wire n_1218;
wire n_13410;
wire n_19581;
wire n_7814;
wire n_8660;
wire n_985;
wire n_2440;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_19546;
wire n_561;
wire n_8606;
wire n_9663;
wire n_16584;
wire n_18340;
wire n_1244;
wire n_9743;
wire n_19048;
wire n_11584;
wire n_2285;
wire n_5280;
wire n_14169;
wire n_7700;
wire n_4451;
wire n_10158;
wire n_10582;
wire n_16151;
wire n_10427;
wire n_11816;
wire n_18808;
wire n_3563;
wire n_16420;
wire n_201;
wire n_11693;
wire n_3495;
wire n_15429;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_10835;
wire n_975;
wire n_11411;
wire n_5576;
wire n_19681;
wire n_13823;
wire n_11386;
wire n_11604;
wire n_13323;
wire n_3359;
wire n_12164;
wire n_16919;
wire n_12824;
wire n_13434;
wire n_16680;
wire n_16938;
wire n_3187;
wire n_10844;
wire n_17793;
wire n_14153;
wire n_6802;
wire n_10654;
wire n_6909;
wire n_13445;
wire n_17177;
wire n_19074;
wire n_18182;
wire n_4336;
wire n_15760;
wire n_16712;
wire n_14746;
wire n_11097;
wire n_4981;
wire n_14606;
wire n_12052;
wire n_9746;
wire n_8073;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_8821;
wire n_9440;
wire n_3955;
wire n_17253;
wire n_2280;
wire n_203;
wire n_1868;
wire n_17264;
wire n_2079;
wire n_15475;
wire n_8663;
wire n_2185;
wire n_5861;
wire n_1836;
wire n_10553;
wire n_19770;
wire n_8309;
wire n_1486;
wire n_5258;
wire n_8945;
wire n_15121;
wire n_10988;
wire n_19209;
wire n_784;
wire n_6112;
wire n_16192;
wire n_18030;
wire n_9041;
wire n_862;
wire n_8166;
wire n_2098;
wire n_5606;
wire n_1935;
wire n_10108;
wire n_13865;
wire n_5920;
wire n_10307;
wire n_1449;
wire n_361;
wire n_8215;
wire n_19538;
wire n_17497;
wire n_6180;
wire n_8809;
wire n_12382;
wire n_5527;
wire n_6476;
wire n_14428;
wire n_6566;
wire n_5172;
wire n_11173;
wire n_16218;
wire n_6872;
wire n_13998;
wire n_5254;
wire n_17825;
wire n_10587;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_7967;
wire n_13522;
wire n_15609;
wire n_16423;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_19016;
wire n_7180;
wire n_13530;
wire n_8604;
wire n_16362;
wire n_7263;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_677;
wire n_14318;
wire n_4686;
wire n_17673;
wire n_17004;
wire n_11802;
wire n_3706;
wire n_8005;
wire n_2179;
wire n_13942;
wire n_18230;
wire n_1547;
wire n_12570;
wire n_11905;
wire n_19326;
wire n_893;
wire n_3801;
wire n_5267;
wire n_10202;
wire n_3564;
wire n_9104;
wire n_15295;
wire n_17050;
wire n_17408;
wire n_15445;
wire n_8272;
wire n_13997;
wire n_14402;
wire n_14882;
wire n_11051;
wire n_11214;
wire n_2628;
wire n_7000;
wire n_7398;
wire n_18335;
wire n_1078;
wire n_14232;
wire n_12882;
wire n_19300;
wire n_18057;
wire n_12617;
wire n_8236;
wire n_13137;
wire n_3345;
wire n_19612;
wire n_15933;
wire n_17188;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_12495;
wire n_10348;
wire n_9581;
wire n_8070;
wire n_4696;
wire n_18468;
wire n_16786;
wire n_7802;
wire n_17118;
wire n_3877;
wire n_15353;
wire n_19623;
wire n_1455;
wire n_6629;
wire n_15993;
wire n_5279;
wire n_5894;
wire n_17699;
wire n_19605;
wire n_8175;
wire n_567;
wire n_8953;
wire n_17546;
wire n_17279;
wire n_19111;
wire n_4814;
wire n_10373;
wire n_3979;
wire n_3077;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_19511;
wire n_6914;
wire n_14121;
wire n_10381;
wire n_713;
wire n_1400;
wire n_10947;
wire n_16984;
wire n_6015;
wire n_11261;
wire n_16012;
wire n_1560;
wire n_734;
wire n_13929;
wire n_17739;
wire n_10767;
wire n_19684;
wire n_14646;
wire n_14095;
wire n_15069;
wire n_14520;
wire n_14780;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_12652;
wire n_15507;
wire n_8142;
wire n_11627;
wire n_6404;
wire n_12209;
wire n_6674;
wire n_5680;
wire n_17883;
wire n_13606;
wire n_11659;
wire n_13501;
wire n_4102;
wire n_9106;
wire n_4662;
wire n_8869;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_17149;
wire n_9520;
wire n_2080;
wire n_14931;
wire n_18774;
wire n_7770;
wire n_6968;
wire n_16268;
wire n_12371;
wire n_4507;
wire n_11497;
wire n_14900;
wire n_792;
wire n_15846;
wire n_13454;
wire n_5306;
wire n_16662;
wire n_9042;
wire n_17329;
wire n_3488;
wire n_8987;
wire n_11805;
wire n_1910;
wire n_14935;
wire n_2998;
wire n_237;
wire n_6282;
wire n_12770;
wire n_4294;
wire n_19551;
wire n_11635;
wire n_15434;
wire n_16530;
wire n_12951;
wire n_9453;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_10281;
wire n_3927;
wire n_3888;
wire n_764;
wire n_12831;
wire n_2895;
wire n_6431;
wire n_733;
wire n_19620;
wire n_15767;
wire n_1290;
wire n_12427;
wire n_1354;
wire n_7533;
wire n_16026;
wire n_7221;
wire n_15159;
wire n_1701;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8246;
wire n_8952;
wire n_3875;
wire n_5609;
wire n_4717;
wire n_871;
wire n_15154;
wire n_9680;
wire n_12172;
wire n_5658;
wire n_4731;
wire n_12923;
wire n_12147;
wire n_3052;
wire n_19624;
wire n_13227;
wire n_19683;
wire n_12825;
wire n_8848;
wire n_5667;
wire n_8259;
wire n_2624;
wire n_5865;
wire n_15182;
wire n_8349;
wire n_6836;
wire n_11998;
wire n_8776;
wire n_19391;
wire n_7753;
wire n_6771;
wire n_14732;
wire n_9947;
wire n_16659;
wire n_1750;
wire n_1462;
wire n_10138;
wire n_12117;
wire n_10375;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_12960;
wire n_18972;
wire n_14094;
wire n_13033;
wire n_15703;
wire n_19353;
wire n_7648;
wire n_515;
wire n_4418;
wire n_12131;
wire n_12851;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_514;
wire n_15518;
wire n_14217;
wire n_10903;
wire n_17596;
wire n_15574;
wire n_14062;
wire n_8453;
wire n_12740;
wire n_2393;
wire n_2921;
wire n_3237;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_17580;
wire n_10517;
wire n_16889;
wire n_10323;
wire n_10842;
wire n_17620;
wire n_3542;
wire n_16465;
wire n_2763;
wire n_2762;
wire n_11146;
wire n_10883;
wire n_17785;
wire n_1296;
wire n_19249;
wire n_3073;
wire n_5343;
wire n_1294;
wire n_3696;
wire n_12278;
wire n_18918;
wire n_19018;
wire n_1779;
wire n_524;
wire n_17672;
wire n_4329;
wire n_18036;
wire n_5135;
wire n_17414;
wire n_10123;
wire n_10651;
wire n_4697;
wire n_3763;
wire n_17483;
wire n_17689;
wire n_18975;
wire n_14785;
wire n_8500;
wire n_17857;
wire n_2145;
wire n_4964;
wire n_12804;
wire n_12116;
wire n_17438;
wire n_1932;
wire n_13755;
wire n_1101;
wire n_10468;
wire n_4636;
wire n_14126;
wire n_14105;
wire n_8285;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_4287;
wire n_19145;
wire n_17696;
wire n_1451;
wire n_639;
wire n_11370;
wire n_16731;
wire n_4576;
wire n_9020;
wire n_4615;
wire n_1018;
wire n_9895;
wire n_16452;
wire n_11585;
wire n_13140;
wire n_13962;
wire n_4389;
wire n_13753;
wire n_1376;
wire n_15365;
wire n_17141;
wire n_948;
wire n_12560;
wire n_19295;
wire n_18171;
wire n_977;
wire n_13610;
wire n_536;
wire n_8851;
wire n_13332;
wire n_15293;
wire n_19405;
wire n_6097;
wire n_19214;
wire n_19779;
wire n_7093;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_432;
wire n_3700;
wire n_3104;
wire n_2239;
wire n_7840;
wire n_18797;
wire n_10024;
wire n_16386;
wire n_17101;
wire n_15695;
wire n_7080;
wire n_17984;
wire n_2191;
wire n_14156;
wire n_10711;
wire n_7624;
wire n_1426;
wire n_16185;
wire n_9186;
wire n_10818;
wire n_1529;
wire n_4634;
wire n_2069;
wire n_18851;
wire n_2362;
wire n_4096;
wire n_15178;
wire n_2698;
wire n_12222;
wire n_11951;
wire n_7003;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_17163;
wire n_10563;
wire n_8810;
wire n_3631;
wire n_2772;
wire n_14518;
wire n_16310;
wire n_16477;
wire n_13397;
wire n_10178;
wire n_5052;
wire n_4541;
wire n_17731;
wire n_15360;
wire n_929;
wire n_4551;
wire n_2857;
wire n_13132;
wire n_6609;
wire n_10115;
wire n_17157;
wire n_5326;
wire n_16927;
wire n_12793;
wire n_11778;
wire n_1183;
wire n_2494;
wire n_12406;
wire n_998;
wire n_717;
wire n_1383;
wire n_7484;
wire n_16639;
wire n_6414;
wire n_1000;
wire n_9470;
wire n_3810;
wire n_552;
wire n_15516;
wire n_3006;
wire n_216;
wire n_13792;
wire n_5010;
wire n_1201;
wire n_4592;
wire n_18229;
wire n_9405;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_17426;
wire n_13480;
wire n_1955;
wire n_19583;
wire n_312;
wire n_13571;
wire n_10984;
wire n_5104;
wire n_19723;
wire n_18742;
wire n_12001;
wire n_7883;
wire n_589;
wire n_1310;
wire n_13715;
wire n_3591;
wire n_16675;
wire n_2797;
wire n_7458;
wire n_4746;
wire n_15186;
wire n_16935;
wire n_18576;
wire n_13810;
wire n_14403;
wire n_7435;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_19292;
wire n_13473;
wire n_18267;
wire n_5985;
wire n_556;
wire n_15963;
wire n_14353;
wire n_16589;
wire n_1602;
wire n_19213;
wire n_11742;
wire n_6891;
wire n_10031;
wire n_276;
wire n_19163;
wire n_12235;
wire n_5232;
wire n_7663;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_14386;
wire n_18784;
wire n_16472;
wire n_17830;
wire n_12098;
wire n_4428;
wire n_1533;
wire n_7917;
wire n_12579;
wire n_2274;
wire n_9203;
wire n_15073;
wire n_7532;
wire n_9613;
wire n_5761;
wire n_13982;
wire n_18703;
wire n_12611;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_7968;
wire n_6382;
wire n_317;
wire n_18542;
wire n_1679;
wire n_9141;
wire n_15867;
wire n_5760;
wire n_2146;
wire n_11027;
wire n_11852;
wire n_5472;
wire n_8377;
wire n_9913;
wire n_2575;
wire n_9286;
wire n_19646;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_10819;
wire n_1179;
wire n_324;
wire n_14521;
wire n_9704;
wire n_19468;
wire n_19025;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_8814;
wire n_8530;
wire n_9193;
wire n_16882;
wire n_7711;
wire n_16181;
wire n_15948;
wire n_8984;
wire n_17123;
wire n_3663;
wire n_3299;
wire n_9290;
wire n_351;
wire n_259;
wire n_14580;
wire n_5745;
wire n_1645;
wire n_14028;
wire n_19131;
wire n_14772;
wire n_956;
wire n_13827;
wire n_14542;
wire n_18632;
wire n_3845;
wire n_664;
wire n_1869;
wire n_7230;
wire n_17552;
wire n_7989;
wire n_9778;
wire n_18986;
wire n_2016;
wire n_5171;
wire n_18280;
wire n_15003;
wire n_13200;
wire n_1937;
wire n_16783;
wire n_12848;
wire n_18963;
wire n_341;
wire n_1744;
wire n_828;
wire n_10315;
wire n_18321;
wire n_607;
wire n_19104;
wire n_17187;
wire n_4028;
wire n_17031;
wire n_11455;
wire n_12368;
wire n_5255;
wire n_3756;
wire n_17240;
wire n_19795;
wire n_3406;
wire n_13193;
wire n_951;
wire n_19798;
wire n_952;
wire n_8462;
wire n_18953;
wire n_9380;
wire n_10062;
wire n_18235;
wire n_19476;
wire n_2375;
wire n_1934;
wire n_8429;
wire n_10514;
wire n_1434;
wire n_12785;
wire n_3981;
wire n_15312;
wire n_14155;
wire n_1275;
wire n_1510;
wire n_7620;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_15818;
wire n_6079;
wire n_16481;
wire n_16430;
wire n_19313;
wire n_3864;
wire n_16715;
wire n_8492;
wire n_16565;
wire n_248;
wire n_2302;
wire n_8135;
wire n_16620;
wire n_8445;
wire n_1037;
wire n_6427;
wire n_3592;
wire n_468;
wire n_4230;
wire n_14978;
wire n_2637;
wire n_18353;
wire n_12639;
wire n_991;
wire n_8895;
wire n_3817;
wire n_7811;
wire n_340;
wire n_14649;
wire n_15940;
wire n_12175;
wire n_5003;
wire n_13536;
wire n_10512;
wire n_14714;
wire n_11384;
wire n_4827;
wire n_8273;
wire n_12353;
wire n_14129;
wire n_6065;
wire n_9761;
wire n_16962;
wire n_4610;
wire n_9087;
wire n_4472;
wire n_17832;
wire n_3081;
wire n_17316;
wire n_15333;
wire n_10434;
wire n_12869;
wire n_8312;
wire n_6781;
wire n_18585;
wire n_13830;
wire n_6133;
wire n_14184;
wire n_11889;
wire n_14183;
wire n_4990;
wire n_6127;
wire n_19172;
wire n_17751;
wire n_2498;
wire n_11362;
wire n_19256;
wire n_8078;
wire n_4515;
wire n_14200;
wire n_6006;
wire n_16558;
wire n_7926;
wire n_19118;
wire n_6598;
wire n_172;
wire n_15568;
wire n_12502;
wire n_2392;
wire n_4131;
wire n_16859;
wire n_1043;
wire n_18800;
wire n_16703;
wire n_2305;
wire n_19666;
wire n_13191;
wire n_10131;
wire n_15464;
wire n_17741;
wire n_6867;
wire n_12600;
wire n_14536;
wire n_16338;
wire n_6139;
wire n_12133;
wire n_7965;
wire n_12919;
wire n_3356;
wire n_10273;
wire n_11416;
wire n_3210;
wire n_937;
wire n_17485;
wire n_14321;
wire n_1682;
wire n_7474;
wire n_11169;
wire n_8650;
wire n_17843;
wire n_14654;
wire n_10503;
wire n_4905;
wire n_14664;
wire n_13215;
wire n_4601;
wire n_16834;
wire n_962;
wire n_10465;
wire n_16073;
wire n_10590;
wire n_3647;
wire n_13782;
wire n_15476;
wire n_8526;
wire n_1186;
wire n_13751;
wire n_17150;
wire n_14019;
wire n_19140;
wire n_19418;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_19806;
wire n_7028;
wire n_9890;
wire n_11492;
wire n_19653;
wire n_394;
wire n_18904;
wire n_6535;
wire n_18801;
wire n_16644;
wire n_9817;
wire n_1524;
wire n_11160;
wire n_18899;
wire n_9782;
wire n_1920;
wire n_3292;
wire n_1225;
wire n_12319;
wire n_10805;
wire n_17214;
wire n_6643;
wire n_17982;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_2506;
wire n_17012;
wire n_14896;
wire n_17440;
wire n_12930;
wire n_17181;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_9069;
wire n_17371;
wire n_3562;
wire n_14030;
wire n_8603;
wire n_17274;
wire n_16660;
wire n_11343;
wire n_3007;
wire n_19143;
wire n_12575;
wire n_11451;
wire n_4571;
wire n_16853;
wire n_3698;
wire n_13384;
wire n_3355;
wire n_2114;
wire n_16048;
wire n_16262;
wire n_17127;
wire n_15422;
wire n_9003;
wire n_2154;
wire n_18874;
wire n_12418;
wire n_5290;
wire n_4185;
wire n_14837;
wire n_7312;
wire n_4219;
wire n_11269;
wire n_16849;
wire n_3985;
wire n_1447;
wire n_14103;
wire n_4774;
wire n_6689;
wire n_7632;
wire n_9172;
wire n_14653;
wire n_4232;
wire n_3000;
wire n_19464;
wire n_17275;
wire n_8980;
wire n_5571;
wire n_17573;
wire n_11311;
wire n_6698;
wire n_18553;
wire n_17345;
wire n_17770;
wire n_13242;
wire n_7707;
wire n_13282;
wire n_14436;
wire n_12113;
wire n_14599;
wire n_16087;
wire n_4736;
wire n_1725;
wire n_3743;
wire n_13352;
wire n_17648;
wire n_18116;
wire n_17853;
wire n_14812;
wire n_17871;
wire n_11293;
wire n_14728;
wire n_19184;
wire n_545;
wire n_2671;
wire n_6363;
wire n_2715;
wire n_8619;
wire n_3511;
wire n_19224;
wire n_18217;
wire n_18812;
wire n_15122;
wire n_10134;
wire n_11603;
wire n_1477;
wire n_7277;
wire n_11271;
wire n_14778;
wire n_15714;
wire n_17270;
wire n_12015;
wire n_8146;
wire n_13690;
wire n_2833;
wire n_11562;
wire n_10194;
wire n_17085;
wire n_8910;
wire n_1001;
wire n_6408;
wire n_6150;
wire n_10077;
wire n_4708;
wire n_13619;
wire n_4657;
wire n_18508;
wire n_12031;
wire n_1191;
wire n_9278;
wire n_855;
wire n_10889;
wire n_10010;
wire n_14996;
wire n_12126;
wire n_14543;
wire n_8550;
wire n_11094;
wire n_14747;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_9739;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_17886;
wire n_1976;
wire n_12195;
wire n_19369;
wire n_6679;
wire n_19294;
wire n_1824;
wire n_13289;
wire n_13182;
wire n_16265;
wire n_16466;
wire n_13324;
wire n_9541;
wire n_11286;
wire n_15215;
wire n_18947;
wire n_17748;
wire n_16379;
wire n_16728;
wire n_823;
wire n_1074;
wire n_7097;
wire n_8140;
wire n_15111;
wire n_1097;
wire n_781;
wire n_18563;
wire n_1810;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_18917;
wire n_1583;
wire n_17621;
wire n_2295;
wire n_1643;
wire n_19570;
wire n_7909;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_15759;
wire n_10734;
wire n_16441;
wire n_15383;
wire n_11560;
wire n_10395;
wire n_3617;
wire n_14966;
wire n_11435;
wire n_1598;
wire n_15255;
wire n_6214;
wire n_9370;
wire n_918;
wire n_13136;
wire n_763;
wire n_6692;
wire n_2485;
wire n_14322;
wire n_12331;
wire n_8093;
wire n_6036;
wire n_13349;
wire n_9956;
wire n_17007;
wire n_6552;
wire n_17096;
wire n_8327;
wire n_13096;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_17005;
wire n_1702;
wire n_4947;
wire n_9487;
wire n_16791;
wire n_14608;
wire n_7306;
wire n_16153;
wire n_10118;
wire n_795;
wire n_18791;
wire n_7470;
wire n_13800;
wire n_19593;
wire n_1245;
wire n_7693;
wire n_3215;
wire n_4740;
wire n_15662;
wire n_1112;
wire n_10002;
wire n_2081;
wire n_911;
wire n_11242;
wire n_17974;
wire n_2862;
wire n_472;
wire n_15923;
wire n_2474;
wire n_3703;
wire n_13694;
wire n_4863;
wire n_17494;
wire n_2267;
wire n_668;
wire n_1821;
wire n_9660;
wire n_16233;
wire n_17344;
wire n_13093;
wire n_9328;
wire n_16511;
wire n_15274;
wire n_16410;
wire n_7653;
wire n_8354;
wire n_14276;
wire n_6959;
wire n_8353;
wire n_6388;
wire n_5045;
wire n_13185;
wire n_11053;
wire n_18635;
wire n_12159;
wire n_9434;
wire n_18450;
wire n_13855;
wire n_10902;
wire n_19596;
wire n_8348;
wire n_7032;
wire n_19086;
wire n_18806;
wire n_8211;
wire n_1816;
wire n_11304;
wire n_9681;
wire n_5848;
wire n_7475;
wire n_10485;
wire n_18448;
wire n_4612;
wire n_6435;
wire n_10536;
wire n_2531;
wire n_9079;
wire n_15544;
wire n_18738;
wire n_19564;
wire n_16145;
wire n_19424;
wire n_17512;
wire n_18931;
wire n_18988;
wire n_714;
wire n_8653;
wire n_8920;
wire n_17521;
wire n_10950;
wire n_5485;
wire n_17477;
wire n_6682;
wire n_6823;
wire n_14550;
wire n_9089;
wire n_4390;
wire n_15346;
wire n_13477;
wire n_18200;
wire n_2095;
wire n_8942;
wire n_10978;
wire n_8222;
wire n_13808;
wire n_6822;
wire n_3295;
wire n_8553;
wire n_1998;
wire n_240;
wire n_19608;
wire n_17068;
wire n_10187;
wire n_11014;
wire n_17508;
wire n_15033;
wire n_2640;
wire n_3288;
wire n_583;
wire n_17789;
wire n_3876;
wire n_9564;
wire n_7391;
wire n_9230;
wire n_19301;
wire n_941;
wire n_19297;
wire n_10768;
wire n_14067;
wire n_6389;
wire n_15903;
wire n_2471;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_13970;
wire n_15247;
wire n_16656;
wire n_4580;
wire n_1055;
wire n_2197;
wire n_10065;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_13408;
wire n_17585;
wire n_15248;
wire n_13727;
wire n_17500;
wire n_13025;
wire n_10268;
wire n_18728;
wire n_14801;
wire n_12601;
wire n_15399;
wire n_17549;
wire n_13641;
wire n_2634;
wire n_1761;
wire n_19588;
wire n_19493;
wire n_8750;
wire n_17473;
wire n_17746;
wire n_5868;
wire n_10305;
wire n_2308;
wire n_16862;
wire n_3001;
wire n_12807;
wire n_15669;
wire n_18018;
wire n_3795;
wire n_7321;
wire n_5289;
wire n_8200;
wire n_4138;
wire n_16055;
wire n_19053;
wire n_18179;
wire n_18564;
wire n_3815;
wire n_12981;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_339;
wire n_434;
wire n_13542;
wire n_288;
wire n_8212;
wire n_5612;
wire n_14426;
wire n_9016;
wire n_15456;
wire n_11545;
wire n_8846;
wire n_4834;
wire n_12665;
wire n_19469;
wire n_16526;
wire n_16397;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_12592;
wire n_17467;
wire n_9029;
wire n_6837;
wire n_3813;
wire n_18860;
wire n_1613;
wire n_11043;
wire n_9414;
wire n_18539;
wire n_7023;
wire n_9615;
wire n_14205;
wire n_1189;
wire n_18532;
wire n_5034;
wire n_726;
wire n_10779;
wire n_11061;
wire n_16495;
wire n_17922;
wire n_5375;
wire n_15742;
wire n_16686;
wire n_16347;
wire n_5370;
wire n_9811;
wire n_5784;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_16385;
wire n_19141;
wire n_1708;
wire n_805;
wire n_14723;
wire n_2051;
wire n_5112;
wire n_19205;
wire n_1402;
wire n_1691;
wire n_10520;
wire n_17437;
wire n_13531;
wire n_7797;
wire n_3668;
wire n_18641;
wire n_13880;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_18251;
wire n_4087;
wire n_7582;
wire n_10541;
wire n_14587;
wire n_8959;
wire n_17326;
wire n_10614;
wire n_18834;
wire n_7809;
wire n_461;
wire n_16877;
wire n_18169;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_9910;
wire n_16790;
wire n_10217;
wire n_17255;
wire n_2513;
wire n_10743;
wire n_2247;
wire n_13424;
wire n_14658;
wire n_15066;
wire n_1579;
wire n_9651;
wire n_3275;
wire n_836;
wire n_15474;
wire n_15316;
wire n_10270;
wire n_11115;
wire n_8001;
wire n_2094;
wire n_1511;
wire n_17417;
wire n_7529;
wire n_14233;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_6881;
wire n_3371;
wire n_19269;
wire n_9544;
wire n_3261;
wire n_17324;
wire n_666;
wire n_7520;
wire n_9831;
wire n_4187;
wire n_940;
wire n_18245;
wire n_9697;
wire n_18878;
wire n_5317;
wire n_18414;
wire n_494;
wire n_8362;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_8256;
wire n_5716;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_12091;
wire n_8704;
wire n_17589;
wire n_6132;
wire n_5211;
wire n_17493;
wire n_9294;
wire n_11747;
wire n_6395;
wire n_976;
wire n_7054;
wire n_2686;
wire n_5327;
wire n_4392;
wire n_11858;
wire n_14027;
wire n_7433;
wire n_16316;
wire n_10075;
wire n_10423;
wire n_17762;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_17291;
wire n_17895;
wire n_5519;
wire n_11895;
wire n_13458;
wire n_4047;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_10886;
wire n_18720;
wire n_13003;
wire n_3791;
wire n_13091;
wire n_6387;
wire n_10192;
wire n_9465;
wire n_13811;
wire n_5139;
wire n_757;
wire n_19459;
wire n_14011;
wire n_166;
wire n_10436;
wire n_19026;
wire n_12794;
wire n_15496;
wire n_6342;
wire n_17744;
wire n_15260;
wire n_15104;
wire n_12483;
wire n_16374;
wire n_18173;
wire n_17251;
wire n_3883;
wire n_18945;
wire n_261;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_5822;
wire n_17381;
wire n_9959;
wire n_15055;
wire n_3949;
wire n_11015;
wire n_18712;
wire n_5364;
wire n_3315;
wire n_9631;
wire n_14751;
wire n_6194;
wire n_4893;
wire n_18313;
wire n_12815;
wire n_15913;
wire n_10431;
wire n_9945;
wire n_1413;
wire n_2228;
wire n_17694;
wire n_5039;
wire n_16314;
wire n_2455;
wire n_4772;
wire n_15115;
wire n_8746;
wire n_11183;
wire n_10019;
wire n_8531;
wire n_12093;
wire n_19296;
wire n_11581;
wire n_4468;
wire n_4161;
wire n_6459;
wire n_8379;
wire n_13100;
wire n_4961;
wire n_4454;
wire n_16154;
wire n_12334;
wire n_18397;
wire n_9209;
wire n_7311;
wire n_3686;
wire n_18234;
wire n_7669;
wire n_8793;
wire n_12355;
wire n_19340;
wire n_15052;
wire n_9767;
wire n_9838;
wire n_1713;
wire n_4277;
wire n_9300;
wire n_11500;
wire n_12943;
wire n_17598;
wire n_530;
wire n_17956;
wire n_618;
wire n_11021;
wire n_8543;
wire n_16502;
wire n_3069;
wire n_7189;
wire n_13067;
wire n_6258;
wire n_16688;
wire n_10243;
wire n_9700;
wire n_18114;
wire n_18802;
wire n_3725;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_5554;
wire n_1175;
wire n_10596;
wire n_19671;
wire n_903;
wire n_12140;
wire n_1802;
wire n_286;
wire n_254;
wire n_8063;
wire n_3961;
wire n_12599;
wire n_2347;
wire n_19419;
wire n_816;
wire n_8032;
wire n_7427;
wire n_2967;
wire n_13250;
wire n_11190;
wire n_11794;
wire n_10519;
wire n_2467;
wire n_17630;
wire n_10163;
wire n_17409;
wire n_3983;
wire n_3538;
wire n_16544;
wire n_2824;
wire n_17529;
wire n_18979;
wire n_12330;
wire n_950;
wire n_8129;
wire n_14819;
wire n_14890;
wire n_15871;
wire n_13906;
wire n_3009;
wire n_5824;
wire n_6760;
wire n_14265;
wire n_13664;
wire n_13566;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_3526;
wire n_4367;
wire n_10874;
wire n_6825;
wire n_19558;
wire n_11831;
wire n_16213;
wire n_14399;
wire n_9628;
wire n_18940;
wire n_19348;
wire n_2583;
wire n_18279;
wire n_19655;
wire n_10250;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_18658;
wire n_14063;
wire n_16657;
wire n_2078;
wire n_2932;
wire n_3431;
wire n_3450;
wire n_17584;
wire n_12041;
wire n_449;
wire n_16734;
wire n_17783;
wire n_2728;
wire n_15157;
wire n_13074;
wire n_3183;
wire n_1067;
wire n_14716;
wire n_255;
wire n_1952;
wire n_12876;
wire n_15286;
wire n_14698;
wire n_19152;
wire n_18633;
wire n_6468;
wire n_3937;
wire n_3159;
wire n_14323;
wire n_18565;
wire n_13071;
wire n_6857;
wire n_3576;
wire n_1863;
wire n_12536;
wire n_10795;
wire n_16333;
wire n_872;
wire n_15116;
wire n_8049;
wire n_7762;
wire n_9467;
wire n_7186;
wire n_13739;
wire n_11157;
wire n_19809;
wire n_9097;
wire n_1513;
wire n_14364;
wire n_15472;
wire n_837;
wire n_5087;
wire n_13234;
wire n_9314;
wire n_7017;
wire n_16718;
wire n_2060;
wire n_7830;
wire n_5131;
wire n_19217;
wire n_17380;
wire n_8084;
wire n_14113;
wire n_8289;
wire n_11178;
wire n_5887;
wire n_16428;
wire n_19010;
wire n_14938;
wire n_14784;
wire n_2816;
wire n_11432;
wire n_14179;
wire n_17755;
wire n_7191;
wire n_14979;
wire n_10412;
wire n_12650;
wire n_4443;
wire n_14324;
wire n_614;
wire n_5460;
wire n_1615;
wire n_4114;
wire n_12859;
wire n_2119;
wire n_17763;
wire n_7961;
wire n_5899;
wire n_17176;
wire n_10617;
wire n_3185;
wire n_2605;
wire n_16524;
wire n_10544;
wire n_13030;
wire n_2848;
wire n_919;
wire n_17819;
wire n_18475;
wire n_15094;
wire n_16880;
wire n_11952;
wire n_6422;
wire n_1299;
wire n_13896;
wire n_5339;
wire n_3837;
wire n_16473;
wire n_1436;
wire n_9873;
wire n_13299;
wire n_13042;
wire n_4818;
wire n_15658;
wire n_10095;
wire n_15873;
wire n_8268;
wire n_6160;
wire n_19749;
wire n_7066;
wire n_18128;
wire n_796;
wire n_7789;
wire n_184;
wire n_6192;
wire n_10056;
wire n_16597;
wire n_17627;
wire n_18815;
wire n_6039;
wire n_2144;
wire n_11919;
wire n_1142;
wire n_11414;
wire n_17705;
wire n_5719;
wire n_17728;
wire n_19457;
wire n_17618;
wire n_7344;
wire n_9888;
wire n_10037;
wire n_2259;
wire n_18029;
wire n_6707;
wire n_12744;
wire n_19601;
wire n_11136;
wire n_19790;
wire n_3142;
wire n_19527;
wire n_19672;
wire n_6787;
wire n_11620;
wire n_15480;
wire n_10179;
wire n_4709;
wire n_2132;
wire n_14038;
wire n_18726;
wire n_11215;
wire n_2860;
wire n_2330;
wire n_11890;
wire n_9366;
wire n_14253;
wire n_7915;
wire n_5893;
wire n_9077;
wire n_2281;
wire n_8406;
wire n_15919;
wire n_16652;
wire n_12443;
wire n_6463;
wire n_11683;
wire n_8554;
wire n_386;
wire n_6051;
wire n_2301;
wire n_7538;
wire n_12934;
wire n_3270;
wire n_19547;
wire n_18981;
wire n_970;
wire n_6799;
wire n_19368;
wire n_444;
wire n_3913;
wire n_3311;
wire n_6487;
wire n_8818;
wire n_16648;
wire n_4348;
wire n_16724;
wire n_10466;
wire n_11953;
wire n_4404;
wire n_439;
wire n_6563;
wire n_2828;
wire n_7554;
wire n_2384;
wire n_4204;
wire n_19005;
wire n_759;
wire n_18881;
wire n_2724;
wire n_15926;
wire n_4513;
wire n_16943;
wire n_11089;
wire n_6341;
wire n_13422;
wire n_7421;
wire n_10166;
wire n_7489;
wire n_1647;
wire n_14702;
wire n_13179;
wire n_15844;
wire n_2306;
wire n_11839;
wire n_18039;
wire n_3683;
wire n_4801;
wire n_13834;
wire n_401;
wire n_18277;
wire n_2550;
wire n_8341;
wire n_11193;
wire n_17800;
wire n_17613;
wire n_7188;
wire n_3736;
wire n_11217;
wire n_15651;
wire n_17759;
wire n_6923;
wire n_9287;
wire n_7991;
wire n_10877;
wire n_16737;
wire n_14686;
wire n_3284;
wire n_12214;
wire n_427;
wire n_16259;
wire n_8926;
wire n_2995;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_13924;
wire n_4149;
wire n_9608;
wire n_501;
wire n_19539;
wire n_8817;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_11488;
wire n_13671;
wire n_14876;
wire n_18571;
wire n_1129;
wire n_6987;
wire n_18265;
wire n_11037;
wire n_16925;
wire n_18740;
wire n_14319;
wire n_2911;
wire n_1429;
wire n_5706;
wire n_16763;
wire n_3429;
wire n_17462;
wire n_1593;
wire n_15287;
wire n_1202;
wire n_7671;
wire n_13150;
wire n_5431;
wire n_15103;
wire n_12541;
wire n_8649;
wire n_19757;
wire n_14818;
wire n_19508;
wire n_8303;
wire n_6153;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_18364;
wire n_11665;
wire n_6579;
wire n_13590;
wire n_16747;
wire n_11138;
wire n_5798;
wire n_575;
wire n_11731;
wire n_5875;
wire n_16257;
wire n_5621;
wire n_16200;
wire n_16041;
wire n_16023;
wire n_732;
wire n_2983;
wire n_6789;
wire n_12100;
wire n_1042;
wire n_15327;
wire n_17718;
wire n_1728;
wire n_13471;
wire n_17615;
wire n_845;
wire n_19063;
wire n_140;
wire n_8862;
wire n_16161;
wire n_10580;
wire n_17287;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_768;
wire n_9675;
wire n_7786;
wire n_16923;
wire n_11454;
wire n_7609;
wire n_3449;
wire n_2598;
wire n_8900;
wire n_597;
wire n_12523;
wire n_6934;
wire n_1403;
wire n_6737;
wire n_18388;
wire n_4488;
wire n_3767;
wire n_8478;
wire n_16988;
wire n_6695;
wire n_12395;
wire n_4211;
wire n_5867;
wire n_17475;
wire n_17363;
wire n_4656;
wire n_3839;
wire n_8497;
wire n_10770;
wire n_6410;
wire n_17873;
wire n_4915;
wire n_15592;
wire n_16064;
wire n_18524;
wire n_15319;
wire n_235;
wire n_5662;
wire n_3730;
wire n_14452;
wire n_17894;
wire n_13464;
wire n_12670;
wire n_16817;
wire n_18336;
wire n_7667;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_17835;
wire n_2737;
wire n_17459;
wire n_10082;
wire n_7182;
wire n_7365;
wire n_10467;
wire n_9849;
wire n_1622;
wire n_17476;
wire n_9856;
wire n_18449;
wire n_17591;
wire n_18672;
wire n_18848;
wire n_11668;
wire n_7885;
wire n_15684;
wire n_2171;
wire n_16720;
wire n_9349;
wire n_17423;
wire n_3136;
wire n_11091;
wire n_4192;
wire n_10940;
wire n_16463;
wire n_15976;
wire n_2808;
wire n_18100;
wire n_17723;
wire n_8839;
wire n_4174;
wire n_12891;
wire n_11615;
wire n_1171;
wire n_11059;
wire n_16403;
wire n_1827;
wire n_14616;
wire n_16799;
wire n_2187;
wire n_6058;
wire n_17965;
wire n_7745;
wire n_12941;
wire n_2872;
wire n_14258;
wire n_12200;
wire n_14024;
wire n_2046;
wire n_17212;
wire n_8684;
wire n_13682;
wire n_6249;
wire n_11060;
wire n_5480;
wire n_18943;
wire n_4831;
wire n_11461;
wire n_10714;
wire n_6969;
wire n_7459;
wire n_6161;
wire n_2970;
wire n_8206;
wire n_18070;
wire n_2882;
wire n_4260;
wire n_18338;
wire n_6607;
wire n_9335;
wire n_1974;
wire n_4122;
wire n_9452;
wire n_11427;
wire n_19293;
wire n_934;
wire n_5284;
wire n_12673;
wire n_14694;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_19208;
wire n_9427;
wire n_17817;
wire n_6294;
wire n_543;
wire n_9611;
wire n_18371;
wire n_9021;
wire n_16269;
wire n_9250;
wire n_11212;
wire n_13145;
wire n_804;
wire n_9550;
wire n_16591;
wire n_11263;
wire n_10641;
wire n_959;
wire n_4312;
wire n_18805;
wire n_16566;
wire n_13195;
wire n_8694;
wire n_13965;
wire n_5048;
wire n_11994;
wire n_13358;
wire n_2195;
wire n_3208;
wire n_18759;
wire n_16693;
wire n_14519;
wire n_6123;
wire n_11000;
wire n_16125;
wire n_4935;
wire n_19403;
wire n_8191;
wire n_10325;
wire n_16354;
wire n_10298;
wire n_6922;
wire n_16701;
wire n_7698;
wire n_12854;
wire n_16427;
wire n_16336;
wire n_8431;
wire n_19631;
wire n_2945;
wire n_3061;
wire n_16248;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_10400;
wire n_19081;
wire n_9177;
wire n_9060;
wire n_11947;
wire n_14496;
wire n_9096;
wire n_13952;
wire n_11697;
wire n_16963;
wire n_18074;
wire n_7891;
wire n_14413;
wire n_8517;
wire n_3008;
wire n_4776;
wire n_4153;
wire n_10901;
wire n_11034;
wire n_10549;
wire n_12115;
wire n_1962;
wire n_11499;
wire n_10825;
wire n_4723;
wire n_17292;
wire n_4269;
wire n_18023;
wire n_14777;
wire n_14057;
wire n_5459;
wire n_17788;
wire n_4143;
wire n_876;
wire n_16406;
wire n_12558;
wire n_11984;
wire n_11948;
wire n_4719;
wire n_7477;
wire n_17028;
wire n_15654;
wire n_1904;
wire n_17289;
wire n_2588;
wire n_11402;
wire n_1353;
wire n_11401;
wire n_17828;
wire n_19679;
wire n_17820;
wire n_2366;
wire n_10581;
wire n_14949;
wire n_17487;
wire n_4423;
wire n_2210;
wire n_3602;
wire n_18372;
wire n_12086;
wire n_1411;
wire n_16952;
wire n_566;
wire n_16449;
wire n_2951;
wire n_11589;
wire n_11246;
wire n_1807;
wire n_18266;
wire n_16606;
wire n_14460;
wire n_13216;
wire n_209;
wire n_12849;
wire n_11312;
wire n_13786;
wire n_5909;
wire n_9344;
wire n_671;
wire n_19719;
wire n_10865;
wire n_740;
wire n_10738;
wire n_7378;
wire n_9798;
wire n_15491;
wire n_14925;
wire n_11612;
wire n_4229;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_13414;
wire n_3865;
wire n_4073;
wire n_5400;
wire n_7498;
wire n_3846;
wire n_11916;
wire n_180;
wire n_3512;
wire n_7501;
wire n_5201;
wire n_10421;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_12764;
wire n_15325;
wire n_1326;
wire n_4783;
wire n_18987;
wire n_19091;
wire n_14238;
wire n_16918;
wire n_12409;
wire n_11625;
wire n_1130;
wire n_17054;
wire n_6592;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_14042;
wire n_9220;
wire n_17312;
wire n_12763;
wire n_378;
wire n_18460;
wire n_17272;
wire n_16394;
wire n_18869;
wire n_15310;
wire n_17989;
wire n_1283;
wire n_4917;
wire n_8698;
wire n_12584;
wire n_14435;
wire n_4432;
wire n_10376;
wire n_15510;
wire n_7515;
wire n_17567;
wire n_344;
wire n_9994;
wire n_14226;
wire n_7309;
wire n_15811;
wire n_5114;
wire n_1392;
wire n_8559;
wire n_5693;
wire n_17670;
wire n_15618;
wire n_2463;
wire n_10224;
wire n_15849;
wire n_611;
wire n_18758;
wire n_3062;
wire n_2679;
wire n_9391;
wire n_16105;
wire n_8514;
wire n_9134;
wire n_14159;
wire n_14515;
wire n_12268;
wire n_18990;
wire n_12077;
wire n_15321;
wire n_14757;
wire n_1017;
wire n_5396;
wire n_12534;
wire n_6846;
wire n_13271;
wire n_11481;
wire n_10175;
wire n_15812;
wire n_16292;
wire n_18458;
wire n_6886;
wire n_17019;
wire n_5365;
wire n_8405;
wire n_15223;
wire n_11350;
wire n_626;
wire n_11925;
wire n_16033;
wire n_8672;
wire n_1104;
wire n_4920;
wire n_1253;
wire n_6446;
wire n_3256;
wire n_9430;
wire n_19279;
wire n_7218;
wire n_11407;
wire n_2118;
wire n_19548;
wire n_12710;
wire n_19331;
wire n_2188;
wire n_8440;
wire n_7005;
wire n_9776;
wire n_16736;
wire n_6777;
wire n_18156;
wire n_11987;
wire n_18208;
wire n_19206;
wire n_8475;
wire n_8029;
wire n_18845;
wire n_18527;
wire n_4861;
wire n_4064;
wire n_1829;
wire n_13089;
wire n_15459;
wire n_15192;
wire n_5266;
wire n_4828;
wire n_1638;
wire n_18360;
wire n_16836;
wire n_13167;
wire n_12329;
wire n_519;
wire n_15013;
wire n_6953;
wire n_3669;
wire n_16710;
wire n_14945;
wire n_4316;
wire n_5122;
wire n_5390;
wire n_18660;
wire n_18348;
wire n_19658;
wire n_18487;
wire n_9834;
wire n_16353;
wire n_2047;
wire n_12318;
wire n_5385;
wire n_13278;
wire n_13597;
wire n_5322;
wire n_3989;
wire n_7089;
wire n_2490;
wire n_18232;
wire n_3841;
wire n_1996;
wire n_6332;
wire n_1442;
wire n_7403;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_4909;
wire n_13938;
wire n_13251;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_18913;
wire n_8317;
wire n_12229;
wire n_269;
wire n_6116;
wire n_7492;
wire n_13319;
wire n_9071;
wire n_10415;
wire n_7694;
wire n_11711;
wire n_18637;
wire n_15666;
wire n_11931;
wire n_8109;
wire n_2055;
wire n_18971;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_7987;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_7434;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_15359;
wire n_9063;
wire n_7787;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_15035;
wire n_18500;
wire n_19085;
wire n_18536;
wire n_6261;
wire n_4281;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_10025;
wire n_412;
wire n_18779;
wire n_6299;
wire n_11753;
wire n_7425;
wire n_19061;
wire n_1059;
wire n_11150;
wire n_18199;
wire n_4360;
wire n_16111;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_9726;
wire n_1748;
wire n_13884;
wire n_17125;
wire n_7719;
wire n_5615;
wire n_6220;
wire n_12783;
wire n_1885;
wire n_1240;
wire n_17671;
wire n_1234;
wire n_14195;
wire n_18363;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_3152;
wire n_7935;
wire n_8458;
wire n_6772;
wire n_16902;
wire n_16646;
wire n_14300;
wire n_6077;
wire n_1003;
wire n_11512;
wire n_17090;
wire n_14678;
wire n_13599;
wire n_17282;
wire n_15008;
wire n_5188;
wire n_13647;
wire n_4490;
wire n_13683;
wire n_1575;
wire n_19094;
wire n_10147;
wire n_17921;
wire n_17197;
wire n_18503;
wire n_9298;
wire n_18058;
wire n_16939;
wire n_14497;
wire n_1991;
wire n_5161;
wire n_14280;
wire n_4078;
wire n_13724;
wire n_9301;
wire n_3046;
wire n_5382;
wire n_12054;
wire n_15827;
wire n_5659;
wire n_8099;
wire n_17256;
wire n_11595;
wire n_17806;
wire n_13768;
wire n_1415;
wire n_16707;
wire n_8578;
wire n_1370;
wire n_7222;
wire n_13838;
wire n_10046;
wire n_2291;
wire n_2184;
wire n_10397;
wire n_2982;
wire n_19379;
wire n_10936;
wire n_12442;
wire n_8611;
wire n_1517;
wire n_8819;
wire n_17927;
wire n_2630;
wire n_15123;
wire n_9835;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_7875;
wire n_13153;
wire n_7643;
wire n_13441;
wire n_16082;
wire n_10207;
wire n_13857;
wire n_18872;
wire n_1143;
wire n_10401;
wire n_19352;
wire n_7242;
wire n_17737;
wire n_19240;
wire n_13816;
wire n_18355;
wire n_2013;
wire n_17215;
wire n_19737;
wire n_14736;
wire n_10139;
wire n_13246;
wire n_14061;
wire n_12986;
wire n_11381;
wire n_16378;
wire n_16109;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_16611;
wire n_16172;
wire n_7746;
wire n_3662;
wire n_2981;
wire n_18108;
wire n_16598;
wire n_16277;
wire n_17588;
wire n_12516;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_6653;
wire n_16806;
wire n_15512;
wire n_18836;
wire n_12377;
wire n_638;
wire n_18486;
wire n_5492;
wire n_9965;
wire n_13650;
wire n_16789;
wire n_887;
wire n_15636;
wire n_15946;
wire n_6501;
wire n_18063;
wire n_9990;
wire n_10005;
wire n_12905;
wire n_11426;
wire n_2599;
wire n_15311;
wire n_8505;
wire n_3368;
wire n_17667;
wire n_7884;
wire n_11258;
wire n_15498;
wire n_7417;
wire n_18097;
wire n_4881;
wire n_12513;
wire n_5734;
wire n_13395;
wire n_4255;
wire n_4071;
wire n_7388;
wire n_3568;
wire n_11657;
wire n_8717;
wire n_5770;
wire n_5705;
wire n_3313;
wire n_9064;
wire n_17420;
wire n_2725;
wire n_14135;
wire n_16482;
wire n_8571;
wire n_4305;
wire n_12514;
wire n_10048;
wire n_16809;
wire n_14194;
wire n_619;
wire n_13825;
wire n_18942;
wire n_8243;
wire n_6347;
wire n_9593;
wire n_606;
wire n_13398;
wire n_8449;
wire n_17605;
wire n_630;
wire n_13204;
wire n_4094;
wire n_14331;
wire n_18994;
wire n_4765;
wire n_2522;
wire n_4364;
wire n_9406;
wire n_8967;
wire n_9322;
wire n_15017;
wire n_5959;
wire n_3720;
wire n_8031;
wire n_15591;
wire n_264;
wire n_12188;
wire n_16609;
wire n_4745;
wire n_5642;
wire n_9232;
wire n_15167;
wire n_12299;
wire n_16739;
wire n_15706;
wire n_1680;
wire n_3842;
wire n_993;
wire n_1605;
wire n_11327;
wire n_4979;
wire n_1988;
wire n_15900;
wire n_12000;
wire n_17281;
wire n_19004;
wire n_1233;
wire n_14182;
wire n_241;
wire n_10279;
wire n_15853;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_14352;
wire n_13889;
wire n_17864;
wire n_7081;
wire n_13015;
wire n_7319;
wire n_15831;
wire n_7644;
wire n_11176;
wire n_9883;
wire n_11135;
wire n_5668;
wire n_11275;
wire n_268;
wire n_18850;
wire n_5463;
wire n_12700;
wire n_12904;
wire n_5489;
wire n_1165;
wire n_14623;
wire n_4773;
wire n_7910;
wire n_6009;
wire n_3281;
wire n_9034;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_8074;
wire n_13639;
wire n_15989;
wire n_8860;
wire n_2676;
wire n_3940;
wire n_1214;
wire n_15514;
wire n_9266;
wire n_3453;
wire n_3410;
wire n_16210;
wire n_10027;
wire n_12784;
wire n_1813;
wire n_18639;
wire n_825;
wire n_12877;
wire n_14261;
wire n_14677;
wire n_18020;
wire n_10616;
wire n_8587;
wire n_5366;
wire n_16016;
wire n_15550;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_9078;
wire n_16297;
wire n_16896;
wire n_13198;
wire n_15914;
wire n_3289;
wire n_13741;
wire n_12610;
wire n_14416;
wire n_11251;
wire n_12293;
wire n_2036;
wire n_6470;
wire n_11598;
wire n_8368;
wire n_15691;
wire n_17560;
wire n_8322;
wire n_16127;
wire n_6187;
wire n_8300;
wire n_9378;
wire n_678;
wire n_12206;
wire n_18112;
wire n_17488;
wire n_17427;
wire n_11400;
wire n_19532;
wire n_6693;
wire n_15848;
wire n_11563;
wire n_362;
wire n_12444;
wire n_18586;
wire n_16409;
wire n_5419;
wire n_14513;
wire n_2943;
wire n_12778;
wire n_12485;
wire n_3253;
wire n_15995;
wire n_14602;
wire n_11468;
wire n_16150;
wire n_4603;
wire n_9683;
wire n_17403;
wire n_15132;
wire n_1527;
wire n_495;
wire n_5732;
wire n_11878;
wire n_15843;
wire n_16666;
wire n_4471;
wire n_15749;
wire n_7449;
wire n_15638;
wire n_16547;
wire n_14289;
wire n_1493;
wire n_16479;
wire n_10751;
wire n_16967;
wire n_10240;
wire n_10691;
wire n_2535;
wire n_9561;
wire n_19351;
wire n_16104;
wire n_9773;
wire n_2436;
wire n_3838;
wire n_9745;
wire n_3941;
wire n_15413;
wire n_10216;
wire n_15628;
wire n_17733;
wire n_1514;
wire n_10150;
wire n_12581;
wire n_17395;
wire n_4994;
wire n_6652;
wire n_10971;
wire n_5168;
wire n_4661;
wire n_18506;
wire n_7674;
wire n_14516;
wire n_18484;
wire n_12305;
wire n_12170;
wire n_2853;
wire n_9630;
wire n_13927;
wire n_13313;
wire n_15308;
wire n_17025;
wire n_9255;
wire n_10231;
wire n_8310;
wire n_16500;
wire n_9758;
wire n_15175;
wire n_8936;
wire n_7126;
wire n_18413;
wire n_15206;
wire n_9691;
wire n_12997;
wire n_14005;
wire n_14293;
wire n_14334;
wire n_7690;
wire n_15245;
wire n_15225;
wire n_3229;
wire n_11223;
wire n_13562;
wire n_14537;
wire n_6950;
wire n_10038;
wire n_17794;
wire n_15614;
wire n_2012;
wire n_5066;
wire n_18101;
wire n_2842;
wire n_19087;
wire n_11221;
wire n_15772;
wire n_14245;
wire n_17659;
wire n_11448;
wire n_17321;
wire n_18272;
wire n_1809;
wire n_8328;
wire n_15502;
wire n_15076;
wire n_12576;
wire n_7258;
wire n_10579;
wire n_13345;
wire n_3677;
wire n_8336;
wire n_3996;
wire n_17492;
wire n_19324;
wire n_4218;
wire n_11445;
wire n_13151;
wire n_3685;
wire n_11552;
wire n_15102;
wire n_14733;
wire n_417;
wire n_14317;
wire n_19807;
wire n_4459;
wire n_16220;
wire n_9852;
wire n_11623;
wire n_3019;
wire n_3471;
wire n_5295;
wire n_2368;
wire n_18599;
wire n_14131;
wire n_10676;
wire n_8041;
wire n_4175;
wire n_10299;
wire n_10540;
wire n_17931;
wire n_16993;
wire n_12845;
wire n_11645;
wire n_10200;
wire n_3259;
wire n_2524;
wire n_13164;
wire n_2460;
wire n_13662;
wire n_3867;
wire n_3593;
wire n_1073;
wire n_16275;
wire n_17062;
wire n_13340;
wire n_17887;
wire n_17192;
wire n_4140;
wire n_2481;
wire n_9939;
wire n_7766;
wire n_19397;
wire n_12797;
wire n_6758;
wire n_5160;
wire n_19709;
wire n_9481;
wire n_7955;
wire n_17081;
wire n_1207;
wire n_12012;
wire n_7287;
wire n_10076;
wire n_880;
wire n_6464;
wire n_18675;
wire n_3540;
wire n_11554;
wire n_150;
wire n_1478;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_4533;
wire n_9635;
wire n_19619;
wire n_1410;
wire n_14308;
wire n_5408;
wire n_1736;
wire n_3848;
wire n_319;
wire n_8181;
wire n_2511;
wire n_8254;
wire n_13452;
wire n_8071;
wire n_5271;
wire n_17480;
wire n_562;
wire n_5964;
wire n_6004;
wire n_11628;
wire n_1136;
wire n_11549;
wire n_17162;
wire n_12286;
wire n_9001;
wire n_19517;
wire n_2329;
wire n_16107;
wire n_14545;
wire n_18031;
wire n_8013;
wire n_146;
wire n_19670;
wire n_193;
wire n_16683;
wire n_17804;
wire n_12347;
wire n_19346;
wire n_17424;
wire n_296;
wire n_651;
wire n_3407;
wire n_5992;
wire n_217;
wire n_1185;
wire n_19394;
wire n_215;
wire n_17818;
wire n_12698;
wire n_2621;
wire n_6540;
wire n_16086;
wire n_5513;
wire n_5614;
wire n_497;
wire n_17383;
wire n_11871;
wire n_16857;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_15326;
wire n_17555;
wire n_18957;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_4056;
wire n_9240;
wire n_8293;
wire n_14726;
wire n_14180;
wire n_18697;
wire n_10548;
wire n_12957;
wire n_11616;
wire n_8791;
wire n_8288;
wire n_1091;
wire n_1425;
wire n_12786;
wire n_983;
wire n_10678;
wire n_6757;
wire n_17752;
wire n_18045;
wire n_1390;
wire n_2289;
wire n_8323;
wire n_10391;
wire n_13176;
wire n_9784;
wire n_19647;
wire n_7990;
wire n_18368;
wire n_10036;
wire n_17631;
wire n_5278;
wire n_14905;
wire n_15128;
wire n_3688;
wire n_8720;
wire n_12205;
wire n_11989;
wire n_16912;
wire n_16215;
wire n_1905;
wire n_14009;
wire n_3466;
wire n_5704;
wire n_15787;
wire n_7148;
wire n_5956;
wire n_9417;
wire n_2139;
wire n_12020;
wire n_18875;
wire n_6835;
wire n_1203;
wire n_11624;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_19290;
wire n_5516;
wire n_2841;
wire n_6247;
wire n_11234;
wire n_10919;
wire n_12099;
wire n_12858;
wire n_4399;
wire n_15351;
wire n_2487;
wire n_18170;
wire n_19159;
wire n_7544;
wire n_9336;
wire n_19750;
wire n_3572;
wire n_8854;
wire n_6645;
wire n_16177;
wire n_10727;
wire n_10885;
wire n_443;
wire n_13201;
wire n_14759;
wire n_13274;
wire n_18621;
wire n_9312;
wire n_5174;
wire n_7469;
wire n_5538;
wire n_5017;
wire n_10895;
wire n_198;
wire n_11977;
wire n_15576;
wire n_11696;
wire n_11734;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11507;
wire n_17290;
wire n_15337;
wire n_17276;
wire n_7082;
wire n_14749;
wire n_18731;
wire n_3108;
wire n_19306;
wire n_11320;
wire n_11837;
wire n_19458;
wire n_8260;
wire n_3417;
wire n_13898;
wire n_16507;
wire n_4124;
wire n_16543;
wire n_11938;
wire n_6418;
wire n_17003;
wire n_5153;
wire n_18814;
wire n_609;
wire n_10571;
wire n_19202;
wire n_19664;
wire n_9807;
wire n_9057;
wire n_8706;
wire n_2607;
wire n_7945;
wire n_8894;
wire n_19244;
wire n_2890;
wire n_12053;
wire n_15947;
wire n_17738;
wire n_12619;
wire n_1320;
wire n_11289;
wire n_13555;
wire n_2499;
wire n_12582;
wire n_5487;
wire n_18919;
wire n_12423;
wire n_15426;
wire n_14137;
wire n_16905;
wire n_17765;
wire n_14163;
wire n_15523;
wire n_2472;
wire n_7328;
wire n_19298;
wire n_10958;
wire n_15682;
wire n_9479;
wire n_15556;
wire n_3957;
wire n_14041;
wire n_18622;
wire n_9181;
wire n_19338;
wire n_19385;
wire n_6578;
wire n_3040;
wire n_14763;
wire n_19319;
wire n_17686;
wire n_18381;
wire n_10879;
wire n_19481;
wire n_5951;
wire n_6589;
wire n_1864;
wire n_10639;
wire n_16359;
wire n_3475;
wire n_17448;
wire n_18657;
wire n_16037;
wire n_9276;
wire n_13351;
wire n_579;
wire n_5152;
wire n_16805;
wire n_15937;
wire n_16141;
wire n_4927;
wire n_5574;
wire n_9821;
wire n_11723;
wire n_4258;
wire n_2699;
wire n_11112;
wire n_650;
wire n_16647;
wire n_1940;
wire n_1405;
wire n_5469;
wire n_14393;
wire n_456;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_6567;
wire n_313;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_3134;
wire n_16231;
wire n_896;
wire n_4553;
wire n_3278;
wire n_17805;
wire n_17318;
wire n_11906;
wire n_2673;
wire n_2456;
wire n_14298;
wire n_9741;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_2871;
wire n_420;
wire n_10180;
wire n_4183;
wire n_14112;
wire n_10650;
wire n_12120;
wire n_12021;
wire n_10157;
wire n_7423;
wire n_10402;
wire n_12515;
wire n_17283;
wire n_9166;
wire n_1640;
wire n_12895;
wire n_12045;
wire n_2141;
wire n_6940;
wire n_12726;
wire n_12668;
wire n_7835;
wire n_15437;
wire n_6320;
wire n_799;
wire n_3044;
wire n_9969;
wire n_11437;
wire n_14068;
wire n_14853;
wire n_11869;
wire n_16735;
wire n_5620;
wire n_10836;
wire n_159;
wire n_16375;
wire n_2125;
wire n_8072;
wire n_13117;
wire n_7130;
wire n_2992;
wire n_1241;
wire n_3221;
wire n_11282;
wire n_17720;
wire n_14700;
wire n_16382;
wire n_7491;
wire n_1706;
wire n_18944;
wire n_18474;
wire n_4052;
wire n_9636;
wire n_7559;
wire n_13175;
wire n_2441;
wire n_9833;
wire n_9095;
wire n_15757;
wire n_18465;
wire n_5907;
wire n_15979;
wire n_19076;
wire n_1559;
wire n_6731;
wire n_4315;
wire n_2888;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_3744;
wire n_12038;
wire n_8210;
wire n_12644;
wire n_1360;
wire n_11826;
wire n_18241;
wire n_3781;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_16764;
wire n_14808;
wire n_2126;
wire n_18135;
wire n_3843;
wire n_11764;
wire n_6600;
wire n_817;
wire n_14140;
wire n_5402;
wire n_10696;
wire n_7355;
wire n_18688;
wire n_9331;
wire n_10170;
wire n_6031;
wire n_14479;
wire n_8331;
wire n_3216;
wire n_332;
wire n_1882;
wire n_18109;
wire n_14172;
wire n_7270;
wire n_591;
wire n_18721;
wire n_5417;
wire n_6967;
wire n_19241;
wire n_6742;
wire n_18117;
wire n_13525;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_14997;
wire n_15931;
wire n_6691;
wire n_14799;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_19062;
wire n_12634;
wire n_14774;
wire n_12680;
wire n_11613;
wire n_10233;
wire n_751;
wire n_19721;
wire n_15492;
wire n_18443;
wire n_17343;
wire n_4652;
wire n_10810;
wire n_12176;
wire n_10311;
wire n_9140;
wire n_2163;
wire n_18533;
wire n_2815;
wire n_19427;
wire n_4577;
wire n_4748;
wire n_337;
wire n_5814;
wire n_12094;
wire n_3231;
wire n_9736;
wire n_2979;
wire n_5531;
wire n_12517;
wire n_6517;
wire n_18431;
wire n_15441;
wire n_9225;
wire n_17353;
wire n_2946;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_3430;
wire n_2269;
wire n_8105;
wire n_9031;
wire n_4225;
wire n_19406;
wire n_13087;
wire n_13972;
wire n_15436;
wire n_17920;
wire n_15633;
wire n_2565;
wire n_12339;
wire n_10602;
wire n_16630;
wire n_14632;
wire n_5655;
wire n_15969;
wire n_6393;
wire n_8154;
wire n_2175;
wire n_2182;
wire n_13849;
wire n_11131;
wire n_10778;
wire n_17961;
wire n_13258;
wire n_1506;
wire n_3473;
wire n_957;
wire n_1994;
wire n_9014;
wire n_13166;
wire n_8509;
wire n_6364;
wire n_16754;
wire n_15482;
wire n_16217;
wire n_19467;
wire n_11003;
wire n_6061;
wire n_18132;
wire n_12723;
wire n_19762;
wire n_14097;
wire n_18741;
wire n_2685;
wire n_8372;
wire n_17042;
wire n_10088;
wire n_14887;
wire n_7225;
wire n_8077;
wire n_18530;
wire n_16948;
wire n_6755;
wire n_18934;
wire n_2265;
wire n_13762;
wire n_13037;
wire n_11573;
wire n_4409;
wire n_7509;
wire n_10145;
wire n_14225;
wire n_11005;
wire n_4629;
wire n_6255;
wire n_18611;
wire n_4638;
wire n_6840;
wire n_17675;
wire n_8423;
wire n_9577;
wire n_19149;
wire n_12589;
wire n_14143;
wire n_6488;
wire n_904;
wire n_8337;
wire n_709;
wire n_7164;
wire n_14044;
wire n_17431;
wire n_3868;
wire n_18249;
wire n_18561;
wire n_18134;
wire n_17000;
wire n_12699;
wire n_1085;
wire n_12927;
wire n_2042;
wire n_16588;
wire n_771;
wire n_8199;
wire n_17456;
wire n_1149;
wire n_8656;
wire n_265;
wire n_14909;
wire n_10918;
wire n_13122;
wire n_2592;
wire n_15553;
wire n_2666;
wire n_1585;
wire n_12663;
wire n_1799;
wire n_2564;
wire n_16349;
wire n_17165;
wire n_15841;
wire n_17623;
wire n_4259;
wire n_2035;
wire n_11127;
wire n_18083;
wire n_7134;
wire n_4572;
wire n_9547;
wire n_4104;
wire n_16350;
wire n_8346;
wire n_8761;
wire n_15458;
wire n_9085;
wire n_13734;
wire n_8226;
wire n_17532;
wire n_7079;
wire n_9084;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_3219;
wire n_14051;
wire n_17680;
wire n_9889;
wire n_12375;
wire n_12556;
wire n_2010;
wire n_1198;
wire n_13723;
wire n_10168;
wire n_2174;
wire n_12156;
wire n_13128;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_17663;
wire n_14913;
wire n_10621;
wire n_9731;
wire n_6572;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_15382;
wire n_4051;
wire n_7755;
wire n_16031;
wire n_6080;
wire n_4865;
wire n_8387;
wire n_12076;
wire n_10613;
wire n_6717;
wire n_7473;
wire n_11359;
wire n_19404;
wire n_19064;
wire n_15997;
wire n_19562;
wire n_10561;
wire n_19335;
wire n_14695;
wire n_16251;
wire n_13212;
wire n_16978;
wire n_15166;
wire n_18304;
wire n_15138;
wire n_16516;
wire n_18517;
wire n_2879;
wire n_17533;
wire n_14405;
wire n_967;
wire n_7038;
wire n_14081;
wire n_4341;
wire n_1819;
wire n_8177;
wire n_17616;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_16137;
wire n_6145;
wire n_6539;
wire n_6926;
wire n_13421;
wire n_1632;
wire n_13495;
wire n_13474;
wire n_14903;
wire n_13949;
wire n_12383;
wire n_11912;
wire n_4973;
wire n_14967;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3950;
wire n_9423;
wire n_16619;
wire n_2927;
wire n_4750;
wire n_12962;
wire n_18823;
wire n_16263;
wire n_11666;
wire n_12459;
wire n_2166;
wire n_2899;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_16369;
wire n_5903;
wire n_17213;
wire n_5986;
wire n_3065;
wire n_6710;
wire n_1423;
wire n_19745;
wire n_18326;
wire n_19402;
wire n_17664;
wire n_4959;
wire n_9056;
wire n_4426;
wire n_12496;
wire n_12814;
wire n_3002;
wire n_649;
wire n_15943;
wire n_18714;
wire n_11921;
wire n_8495;
wire n_14532;
wire n_8783;
wire n_14557;
wire n_19805;
wire n_1199;
wire n_12603;
wire n_15392;
wire n_14340;
wire n_18444;
wire n_14032;
wire n_16944;
wire n_15702;
wire n_7262;
wire n_212;
wire n_3773;
wire n_12967;
wire n_14899;
wire n_12232;
wire n_18115;
wire n_18847;
wire n_11859;
wire n_15773;
wire n_798;
wire n_19771;
wire n_15307;
wire n_14111;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9553;
wire n_11633;
wire n_7506;
wire n_8551;
wire n_14361;
wire n_12760;
wire n_18291;
wire n_2647;
wire n_19633;
wire n_14943;
wire n_4578;
wire n_4777;
wire n_2672;
wire n_12590;
wire n_2299;
wire n_15605;
wire n_5871;
wire n_18951;
wire n_17711;
wire n_12577;
wire n_7142;
wire n_10182;
wire n_16813;
wire n_13928;
wire n_19342;
wire n_7125;
wire n_1172;
wire n_11655;
wire n_3626;
wire n_2313;
wire n_12069;
wire n_16899;
wire n_15656;
wire n_18455;
wire n_16957;
wire n_10317;
wire n_4029;
wire n_375;
wire n_12270;
wire n_4617;
wire n_16021;
wire n_9196;
wire n_4010;
wire n_1649;
wire n_5882;
wire n_5650;
wire n_6057;
wire n_14555;
wire n_10893;
wire n_1572;
wire n_5021;
wire n_9251;
wire n_9973;
wire n_11117;
wire n_8064;
wire n_8468;
wire n_4325;
wire n_3251;
wire n_10201;
wire n_2212;
wire n_12210;
wire n_8778;
wire n_17106;
wire n_14168;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_15342;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_5625;
wire n_11777;
wire n_17402;
wire n_4919;
wire n_3737;
wire n_13975;
wire n_5969;
wire n_10121;
wire n_8198;
wire n_19054;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_12189;
wire n_1211;
wire n_9270;
wire n_14142;
wire n_6041;
wire n_9099;
wire n_7350;
wire n_10814;
wire n_5276;
wire n_16034;
wire n_9627;
wire n_17008;
wire n_16563;
wire n_6664;
wire n_196;
wire n_17575;
wire n_2985;
wire n_13131;
wire n_14941;
wire n_1446;
wire n_3938;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_5855;
wire n_3531;
wire n_16128;
wire n_10975;
wire n_1054;
wire n_9460;
wire n_17698;
wire n_11652;
wire n_14320;
wire n_11056;
wire n_19229;
wire n_6238;
wire n_13932;
wire n_2397;
wire n_16804;
wire n_3931;
wire n_15606;
wire n_10459;
wire n_2113;
wire n_1918;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_15866;
wire n_9766;
wire n_4163;
wire n_10463;
wire n_14764;
wire n_645;
wire n_7074;
wire n_8734;
wire n_2633;
wire n_12564;
wire n_19443;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_7037;
wire n_13697;
wire n_11784;
wire n_5298;
wire n_9025;
wire n_3396;
wire n_14244;
wire n_7928;
wire n_12886;
wire n_6532;
wire n_821;
wire n_4372;
wire n_7293;
wire n_18638;
wire n_13000;
wire n_14362;
wire n_5640;
wire n_15996;
wire n_408;
wire n_4318;
wire n_6721;
wire n_18825;
wire n_2123;
wire n_3716;
wire n_6108;
wire n_10370;
wire n_8258;
wire n_18537;
wire n_9597;
wire n_11892;
wire n_5744;
wire n_5384;
wire n_3248;
wire n_15731;
wire n_134;
wire n_8299;
wire n_12473;
wire n_4032;
wire n_1064;
wire n_11421;
wire n_1396;
wire n_18704;
wire n_11966;
wire n_19530;
wire n_17450;
wire n_18011;
wire n_12748;
wire n_4337;
wire n_16829;
wire n_3092;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_3734;
wire n_17305;
wire n_18047;
wire n_7078;
wire n_13831;
wire n_2580;
wire n_8188;
wire n_16792;
wire n_18572;
wire n_11423;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_18378;
wire n_9567;
wire n_9061;
wire n_3419;
wire n_1297;
wire n_17154;
wire n_16922;
wire n_8664;
wire n_922;
wire n_16552;
wire n_16867;
wire n_16638;
wire n_14783;
wire n_13268;
wire n_10740;
wire n_10457;
wire n_19042;
wire n_17968;
wire n_1896;
wire n_3058;
wire n_14158;
wire n_9701;
wire n_675;
wire n_19247;
wire n_14236;
wire n_1540;
wire n_18849;
wire n_13510;
wire n_14640;
wire n_6659;
wire n_9709;
wire n_242;
wire n_9295;
wire n_4371;
wire n_2994;
wire n_3689;
wire n_16678;
wire n_10264;
wire n_5850;
wire n_15029;
wire n_14286;
wire n_12528;
wire n_17640;
wire n_6182;
wire n_12717;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_1965;
wire n_2476;
wire n_17651;
wire n_17662;
wire n_598;
wire n_11547;
wire n_19680;
wire n_13520;
wire n_19668;
wire n_8501;
wire n_10301;
wire n_3271;
wire n_295;
wire n_4248;
wire n_13018;
wire n_18240;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_15139;
wire n_8076;
wire n_6826;
wire n_1792;
wire n_11395;
wire n_9107;
wire n_19630;
wire n_3809;
wire n_11279;
wire n_18370;
wire n_11724;
wire n_11789;
wire n_14152;
wire n_3139;
wire n_14869;
wire n_19354;
wire n_881;
wire n_8014;
wire n_19030;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_4018;
wire n_14651;
wire n_694;
wire n_7982;
wire n_8804;
wire n_297;
wire n_3337;
wire n_11383;
wire n_1044;
wire n_2165;
wire n_15882;
wire n_17740;
wire n_6879;
wire n_17059;
wire n_7567;
wire n_8433;
wire n_6074;
wire n_4588;
wire n_585;
wire n_10932;
wire n_10619;
wire n_1756;
wire n_5411;
wire n_17263;
wire n_9156;
wire n_16113;
wire n_16848;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_18749;
wire n_10248;
wire n_9748;
wire n_3616;
wire n_13365;
wire n_7771;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_16289;
wire n_2151;
wire n_7701;
wire n_16342;
wire n_1839;
wire n_17278;
wire n_5235;
wire n_6720;
wire n_11930;
wire n_6888;
wire n_826;
wire n_3747;
wire n_12628;
wire n_8122;
wire n_17095;
wire n_13444;
wire n_16504;
wire n_8432;
wire n_4330;
wire n_7592;
wire n_14209;
wire n_19462;
wire n_18651;
wire n_5311;
wire n_6590;
wire n_3522;
wire n_2747;
wire n_18243;
wire n_791;
wire n_11876;
wire n_5572;
wire n_19110;
wire n_7151;
wire n_8950;
wire n_18683;
wire n_10758;
wire n_2861;
wire n_13431;
wire n_3975;
wire n_1838;
wire n_4683;
wire n_12538;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_2316;
wire n_15954;
wire n_9355;
wire n_5060;
wire n_15386;
wire n_4986;
wire n_14620;
wire n_5888;
wire n_15349;
wire n_9582;
wire n_2208;
wire n_5884;
wire n_11009;
wire n_9288;
wire n_6308;
wire n_7897;
wire n_17701;
wire n_7118;
wire n_2134;
wire n_8284;
wire n_9702;
wire n_18767;
wire n_15378;
wire n_7422;
wire n_1431;
wire n_17881;
wire n_3835;
wire n_6738;
wire n_12307;
wire n_8703;
wire n_15839;
wire n_16135;
wire n_17661;
wire n_14999;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_19377;
wire n_3557;
wire n_2610;
wire n_3620;
wire n_13720;
wire n_478;
wire n_7339;
wire n_3832;
wire n_13706;
wire n_13903;
wire n_3693;
wire n_9051;
wire n_8545;
wire n_10385;
wire n_10105;
wire n_2372;
wire n_1490;
wire n_15785;
wire n_19056;
wire n_3674;
wire n_2959;
wire n_17114;
wire n_10251;
wire n_15234;
wire n_293;
wire n_18796;
wire n_1070;
wire n_2403;
wire n_4700;
wire n_17524;
wire n_9980;
wire n_14394;
wire n_4224;
wire n_18679;
wire n_6005;
wire n_17261;
wire n_9555;
wire n_14845;
wire n_1358;
wire n_7713;
wire n_4564;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_16182;
wire n_2424;
wire n_3201;
wire n_19239;
wire n_1475;
wire n_10304;
wire n_3103;
wire n_5860;
wire n_6936;
wire n_15934;
wire n_16827;
wire n_16121;
wire n_7487;
wire n_9986;
wire n_527;
wire n_13794;
wire n_3627;
wire n_13537;
wire n_9397;
wire n_18616;
wire n_1137;
wire n_3612;
wire n_17574;
wire n_4695;
wire n_9855;
wire n_10568;
wire n_2966;
wire n_2294;
wire n_13463;
wire n_600;
wire n_9496;
wire n_16241;
wire n_10796;
wire n_10016;
wire n_10030;
wire n_12864;
wire n_9653;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_1339;
wire n_13936;
wire n_13933;
wire n_7815;
wire n_403;
wire n_7934;
wire n_3244;
wire n_11578;
wire n_6865;
wire n_1141;
wire n_7276;
wire n_18595;
wire n_1755;
wire n_5043;
wire n_8739;
wire n_17078;
wire n_6747;
wire n_13714;
wire n_2025;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_2250;
wire n_3033;
wire n_16079;
wire n_11908;
wire n_18166;
wire n_6462;
wire n_17372;
wire n_6034;
wire n_13159;
wire n_9781;
wire n_418;
wire n_14788;
wire n_13287;
wire n_11913;
wire n_7034;
wire n_1618;
wire n_4867;
wire n_13389;
wire n_17726;
wire n_1653;
wire n_9906;
wire n_4237;
wire n_5029;
wire n_12317;
wire n_13302;
wire n_10092;
wire n_6833;
wire n_6793;
wire n_16766;
wire n_17834;
wire n_11815;
wire n_6295;
wire n_3386;
wire n_11231;
wire n_463;
wire n_13740;
wire n_17966;
wire n_19278;
wire n_8137;
wire n_12027;
wire n_3205;
wire n_15218;
wire n_17366;
wire n_19114;
wire n_17514;
wire n_17975;
wire n_7014;
wire n_10430;
wire n_16697;
wire n_8305;
wire n_18147;
wire n_1636;
wire n_4001;
wire n_18751;
wire n_6709;
wire n_17525;
wire n_960;
wire n_6712;
wire n_7416;
wire n_778;
wire n_14553;
wire n_5177;
wire n_9657;
wire n_16594;
wire n_16370;
wire n_6743;
wire n_16223;
wire n_1610;
wire n_12412;
wire n_11880;
wire n_5785;
wire n_14528;
wire n_4583;
wire n_9485;
wire n_13940;
wire n_2515;
wire n_11249;
wire n_15449;
wire n_4054;
wire n_10119;
wire n_11986;
wire n_14798;
wire n_5966;
wire n_3349;
wire n_17579;
wire n_368;
wire n_12118;
wire n_14409;
wire n_14724;
wire n_18451;
wire n_14291;
wire n_1020;
wire n_8625;
wire n_4214;
wire n_6919;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_9192;
wire n_1138;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_8179;
wire n_19360;
wire n_11861;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_4413;
wire n_7453;
wire n_10684;
wire n_2381;
wire n_18095;
wire n_2052;
wire n_5081;
wire n_15039;
wire n_17929;
wire n_17027;
wire n_8806;
wire n_17400;
wire n_6619;
wire n_19234;
wire n_16434;
wire n_5189;
wire n_13930;
wire n_8149;
wire n_3041;
wire n_603;
wire n_10390;
wire n_1657;
wire n_7210;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_6718;
wire n_4238;
wire n_3011;
wire n_15400;
wire n_2061;
wire n_17411;
wire n_16866;
wire n_15485;
wire n_18499;
wire n_18789;
wire n_14841;
wire n_16726;
wire n_13624;
wire n_5632;
wire n_5425;
wire n_18603;
wire n_19480;
wire n_8269;
wire n_13805;
wire n_18786;
wire n_3650;
wire n_16243;
wire n_8968;
wire n_7855;
wire n_14029;
wire n_4590;
wire n_3137;
wire n_14056;
wire n_5678;
wire n_13695;
wire n_6981;
wire n_13288;
wire n_19465;
wire n_16917;
wire n_3238;
wire n_218;
wire n_11519;
wire n_13065;
wire n_11229;
wire n_18655;
wire n_16159;
wire n_17570;
wire n_11397;
wire n_12840;
wire n_5437;
wire n_12846;
wire n_14705;
wire n_17660;
wire n_8401;
wire n_7854;
wire n_10577;
wire n_11324;
wire n_12945;
wire n_5307;
wire n_17385;
wire n_10151;
wire n_6439;
wire n_2446;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_16193;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_9305;
wire n_9999;
wire n_17495;
wire n_1121;
wire n_11361;
wire n_1963;
wire n_6945;
wire n_18617;
wire n_3790;
wire n_7029;
wire n_19009;
wire n_10186;
wire n_17236;
wire n_11841;
wire n_6618;
wire n_14453;
wire n_17545;
wire n_13094;
wire n_7317;
wire n_17558;
wire n_3977;
wire n_227;
wire n_9461;
wire n_6816;
wire n_10928;
wire n_5008;
wire n_6502;
wire n_6250;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_4133;
wire n_9618;
wire n_6118;
wire n_18961;
wire n_4561;
wire n_464;
wire n_19772;
wire n_11808;
wire n_17970;
wire n_13257;
wire n_17160;
wire n_18778;
wire n_4239;
wire n_18509;
wire n_4184;
wire n_17636;
wire n_1830;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_13922;
wire n_13423;
wire n_18149;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2293;
wire n_10252;
wire n_16641;
wire n_11555;
wire n_6869;
wire n_3102;
wire n_14625;
wire n_10345;
wire n_2026;
wire n_10059;
wire n_8325;
wire n_7621;
wire n_7359;
wire n_550;
wire n_3321;
wire n_2322;
wire n_12394;
wire n_4782;
wire n_13578;
wire n_19540;
wire n_14204;
wire n_9005;
wire n_4378;
wire n_8274;
wire n_12954;
wire n_4876;
wire n_19703;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_14688;
wire n_10644;
wire n_12801;
wire n_18594;
wire n_13708;
wire n_10365;
wire n_11781;
wire n_9648;
wire n_2653;
wire n_12965;
wire n_12788;
wire n_9498;
wire n_15707;
wire n_16328;
wire n_3156;
wire n_15396;
wire n_19804;
wire n_15909;
wire n_672;
wire n_3483;
wire n_11884;
wire n_19516;
wire n_19734;
wire n_13371;
wire n_4493;
wire n_7971;
wire n_743;
wire n_12264;
wire n_8232;
wire n_9649;
wire n_8904;
wire n_16977;
wire n_19287;
wire n_10629;
wire n_660;
wire n_7070;
wire n_8382;
wire n_4421;
wire n_18950;
wire n_2839;
wire n_4793;
wire n_13856;
wire n_15607;
wire n_15879;
wire n_7259;
wire n_12274;
wire n_14588;
wire n_2944;
wire n_8128;
wire n_15746;
wire n_3831;
wire n_15921;
wire n_19545;
wire n_5932;
wire n_5830;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12586;
wire n_3391;
wire n_8794;
wire n_11760;
wire n_19203;
wire n_1463;
wire n_4505;
wire n_17222;
wire n_1826;
wire n_5126;
wire n_8205;
wire n_9907;
wire n_13088;
wire n_6976;
wire n_13538;
wire n_11024;
wire n_18437;
wire n_6304;
wire n_5236;
wire n_7640;
wire n_13701;
wire n_10498;
wire n_11424;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_1256;
wire n_10635;
wire n_13626;
wire n_19218;
wire n_12832;
wire n_8067;
wire n_12301;
wire n_9643;
wire n_4630;
wire n_18973;
wire n_18402;
wire n_15822;
wire n_11881;
wire n_14980;
wire n_2109;
wire n_7727;
wire n_18968;
wire n_11935;
wire n_17561;
wire n_18766;
wire n_1204;
wire n_18901;
wire n_233;
wire n_8719;
wire n_16140;
wire n_19223;
wire n_18046;
wire n_2787;
wire n_15493;
wire n_12615;
wire n_13357;
wire n_10802;
wire n_17148;
wire n_769;
wire n_4786;
wire n_7565;
wire n_16624;
wire n_7631;
wire n_13869;
wire n_16903;
wire n_7387;
wire n_9212;
wire n_12167;
wire n_9473;
wire n_13026;
wire n_10490;
wire n_15019;
wire n_13499;
wire n_17107;
wire n_14843;
wire n_2736;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_16781;
wire n_19738;
wire n_12298;
wire n_10081;
wire n_3774;
wire n_12569;
wire n_2910;
wire n_14929;
wire n_18497;
wire n_5148;
wire n_2584;
wire n_866;
wire n_12456;
wire n_8655;
wire n_17039;
wire n_10808;
wire n_6333;
wire n_8745;
wire n_5791;
wire n_18504;
wire n_8086;
wire n_15466;
wire n_13943;
wire n_17124;
wire n_7379;
wire n_17530;
wire n_11078;
wire n_8901;
wire n_8695;
wire n_4911;
wire n_8173;
wire n_12072;
wire n_4436;
wire n_10545;
wire n_1174;
wire n_17945;
wire n_16557;
wire n_14141;
wire n_5602;
wire n_647;
wire n_9379;
wire n_11992;
wire n_15790;
wire n_844;
wire n_17061;
wire n_14880;
wire n_13142;
wire n_13180;
wire n_3584;
wire n_10453;
wire n_16975;
wire n_3556;
wire n_16716;
wire n_13785;
wire n_5831;
wire n_7742;
wire n_9274;
wire n_3456;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_17230;
wire n_12863;
wire n_10352;
wire n_19449;
wire n_1122;
wire n_4059;
wire n_16830;
wire n_1109;
wire n_17851;
wire n_3309;
wire n_8507;
wire n_8415;
wire n_2609;
wire n_10713;
wire n_6680;
wire n_10954;
wire n_7432;
wire n_16036;
wire n_13978;
wire n_13941;
wire n_15339;
wire n_13439;
wire n_228;
wire n_16152;
wire n_14133;
wire n_14433;
wire n_13187;
wire n_13162;
wire n_2600;
wire n_7505;
wire n_18521;
wire n_15059;
wire n_8244;
wire n_7494;
wire n_18380;
wire n_4353;
wire n_735;
wire n_17071;
wire n_13661;
wire n_9546;
wire n_7589;
wire n_17764;
wire n_4346;
wire n_4351;
wire n_11296;
wire n_13770;
wire n_18636;
wire n_8723;
wire n_13511;
wire n_18016;
wire n_11019;
wire n_980;
wire n_7843;
wire n_1651;
wire n_19544;
wire n_4784;
wire n_19258;
wire n_14569;
wire n_7902;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_15744;
wire n_7756;
wire n_2844;
wire n_15557;
wire n_18244;
wire n_8940;
wire n_8342;
wire n_14154;
wire n_8472;
wire n_4332;
wire n_810;
wire n_10000;
wire n_12812;
wire n_7988;
wire n_14174;
wire n_7500;
wire n_10246;
wire n_3198;
wire n_18236;
wire n_14269;
wire n_9822;
wire n_13991;
wire n_17523;
wire n_14821;
wire n_17330;
wire n_15096;
wire n_5272;
wire n_14992;
wire n_10125;
wire n_9065;
wire n_16637;
wire n_3218;
wire n_18627;
wire n_9153;
wire n_9086;
wire n_10505;
wire n_582;
wire n_861;
wire n_11064;
wire n_6908;
wire n_8237;
wire n_9093;
wire n_19046;
wire n_2968;
wire n_4201;
wire n_7266;
wire n_17928;
wire n_8046;
wire n_5646;
wire n_13284;
wire n_4852;
wire n_4210;
wire n_16521;
wire n_2709;
wire n_9198;
wire n_8335;
wire n_9142;
wire n_17697;
wire n_15820;
wire n_18239;
wire n_5214;
wire n_15486;
wire n_9493;
wire n_19371;
wire n_11330;
wire n_12720;
wire n_7794;
wire n_19139;
wire n_13318;
wire n_15917;
wire n_1274;
wire n_3333;
wire n_6605;
wire n_12687;
wire n_18278;
wire n_19748;
wire n_17510;
wire n_19106;
wire n_13208;
wire n_13867;
wire n_15594;
wire n_17807;
wire n_17841;
wire n_5380;
wire n_5776;
wire n_11796;
wire n_18339;
wire n_16881;
wire n_12789;
wire n_2677;
wire n_12127;
wire n_17232;
wire n_3283;
wire n_16976;
wire n_8037;
wire n_13673;
wire n_14119;
wire n_1742;
wire n_16775;
wire n_12573;
wire n_2542;
wire n_1671;
wire n_19400;
wire n_15214;
wire n_13045;
wire n_741;
wire n_1351;
wire n_17347;
wire n_18684;
wire n_6806;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_5019;
wire n_2332;
wire n_5138;
wire n_4388;
wire n_6960;
wire n_3089;
wire n_8169;
wire n_12265;
wire n_783;
wire n_5409;
wire n_5301;
wire n_17777;
wire n_188;
wire n_1854;
wire n_3222;
wire n_7504;
wire n_15971;
wire n_442;
wire n_11678;
wire n_8023;
wire n_12251;
wire n_1975;
wire n_16307;
wire n_8130;
wire n_16911;
wire n_15294;
wire n_5055;
wire n_18676;
wire n_16288;
wire n_7116;
wire n_4249;
wire n_17992;
wire n_6999;
wire n_14741;
wire n_11046;
wire n_11079;
wire n_5548;
wire n_15581;
wire n_11065;
wire n_8339;
wire n_19058;
wire n_14215;
wire n_17368;
wire n_852;
wire n_544;
wire n_5900;
wire n_4273;
wire n_18104;
wire n_8499;
wire n_15356;
wire n_18525;
wire n_6882;
wire n_10775;
wire n_2129;
wire n_9526;
wire n_17511;
wire n_18762;
wire n_15571;
wire n_7983;
wire n_10863;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_17138;
wire n_17700;
wire n_13993;
wire n_10986;
wire n_8366;
wire n_8102;
wire n_19126;
wire n_18087;
wire n_8022;
wire n_17226;
wire n_19212;
wire n_10262;
wire n_5239;
wire n_1781;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_2004;
wire n_1106;
wire n_18183;
wire n_8913;
wire n_155;
wire n_4956;
wire n_16772;
wire n_14699;
wire n_454;
wire n_10335;
wire n_15362;
wire n_5129;
wire n_11301;
wire n_15101;
wire n_5070;
wire n_18154;
wire n_11703;
wire n_6374;
wire n_17013;
wire n_6628;
wire n_13483;
wire n_18923;
wire n_4262;
wire n_16551;
wire n_17803;
wire n_1894;
wire n_6570;
wire n_8556;
wire n_8040;
wire n_11821;
wire n_13121;
wire n_13989;
wire n_10755;
wire n_16998;
wire n_15200;
wire n_17349;
wire n_10682;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_2613;
wire n_3535;
wire n_8595;
wire n_2708;
wire n_1648;
wire n_2011;
wire n_5684;
wire n_15887;
wire n_10022;
wire n_5729;
wire n_13803;
wire n_14066;
wire n_7856;
wire n_564;
wire n_6148;
wire n_7625;
wire n_686;
wire n_1641;
wire n_3871;
wire n_12775;
wire n_7863;
wire n_6989;
wire n_8958;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_13687;
wire n_7623;
wire n_7217;
wire n_1699;
wire n_14540;
wire n_16784;
wire n_8115;
wire n_608;
wire n_2101;
wire n_9398;
wire n_15320;
wire n_3484;
wire n_4677;
wire n_12915;
wire n_6196;
wire n_13149;
wire n_18748;
wire n_2616;
wire n_5275;
wire n_14091;
wire n_15755;
wire n_8412;
wire n_2811;
wire n_6485;
wire n_14478;
wire n_17848;
wire n_10177;
wire n_6107;
wire n_16689;
wire n_11944;
wire n_1075;
wire n_7796;
wire n_6994;
wire n_15986;
wire n_14570;
wire n_16068;
wire n_13797;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_175;
wire n_9446;
wire n_11129;
wire n_7234;
wire n_3914;
wire n_8119;
wire n_10296;
wire n_8641;
wire n_12988;
wire n_17136;
wire n_13344;
wire n_11139;
wire n_17766;
wire n_12685;
wire n_8436;
wire n_14239;
wire n_8659;
wire n_14045;
wire n_19575;
wire n_4369;
wire n_7849;
wire n_12667;
wire n_18747;
wire n_15635;
wire n_4331;
wire n_7297;
wire n_15183;
wire n_10018;
wire n_4972;
wire n_4993;
wire n_15118;
wire n_7298;
wire n_5536;
wire n_10141;
wire n_9129;
wire n_14162;
wire n_8224;
wire n_2678;
wire n_15679;
wire n_4613;
wire n_13014;
wire n_19744;
wire n_1167;
wire n_2428;
wire n_10897;
wire n_210;
wire n_10449;
wire n_7861;
wire n_14303;
wire n_7039;
wire n_11349;
wire n_5046;
wire n_2749;
wire n_3273;
wire n_7077;
wire n_12540;
wire n_19160;
wire n_5305;
wire n_4681;
wire n_13239;
wire n_15942;
wire n_17583;
wire n_4752;
wire n_18552;
wire n_9143;
wire n_8287;
wire n_2092;
wire n_7950;
wire n_8607;
wire n_2514;
wire n_604;
wire n_17032;
wire n_6248;
wire n_16768;
wire n_16134;
wire n_10452;
wire n_7806;
wire n_3942;
wire n_15928;
wire n_16092;
wire n_7595;
wire n_8066;
wire n_5795;
wire n_12349;
wire n_14282;
wire n_5552;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_890;
wire n_16266;
wire n_8416;
wire n_4518;
wire n_14167;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_10363;
wire n_2252;
wire n_13623;
wire n_11511;
wire n_15833;
wire n_16046;
wire n_760;
wire n_9393;
wire n_15974;
wire n_13845;
wire n_12709;
wire n_13432;
wire n_12771;
wire n_17760;
wire n_1858;
wire n_14787;
wire n_19502;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_17100;
wire n_10781;
wire n_7315;
wire n_9886;
wire n_1164;
wire n_13244;
wire n_4288;
wire n_18969;
wire n_6185;
wire n_5529;
wire n_3733;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_17191;
wire n_13404;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_18689;
wire n_7268;
wire n_4228;
wire n_3423;
wire n_10094;
wire n_16295;
wire n_10084;
wire n_19259;
wire n_13870;
wire n_13791;
wire n_3644;
wire n_6955;
wire n_2706;
wire n_1127;
wire n_1512;
wire n_9932;
wire n_16745;
wire n_320;
wire n_13900;
wire n_16224;
wire n_14652;
wire n_1139;
wire n_3179;
wire n_8741;
wire n_4000;
wire n_2897;
wire n_3970;
wire n_7232;
wire n_7377;
wire n_19461;
wire n_996;
wire n_16132;
wire n_19425;
wire n_6646;
wire n_19789;
wire n_15149;
wire n_14844;
wire n_16907;
wire n_14391;
wire n_6033;
wire n_11541;
wire n_15495;
wire n_4873;
wire n_9801;
wire n_19312;
wire n_3782;
wire n_8773;
wire n_6369;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_581;
wire n_7542;
wire n_5636;
wire n_13213;
wire n_12231;
wire n_989;
wire n_17643;
wire n_8410;
wire n_14756;
wire n_18144;
wire n_7739;
wire n_4939;
wire n_19474;
wire n_14384;
wire n_15905;
wire n_5530;
wire n_2473;
wire n_12552;
wire n_11069;
wire n_2539;
wire n_4123;
wire n_5595;
wire n_9941;
wire n_16795;
wire n_17131;
wire n_3119;
wire n_3735;
wire n_11369;
wire n_4379;
wire n_14210;
wire n_486;
wire n_5388;
wire n_4718;
wire n_15788;
wire n_13362;
wire n_5962;
wire n_7010;
wire n_648;
wire n_9728;
wire n_16690;
wire n_2057;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_15694;
wire n_8774;
wire n_18690;
wire n_19494;
wire n_7299;
wire n_4872;
wire n_9936;
wire n_6195;
wire n_9530;
wire n_14692;
wire n_7471;
wire n_10455;
wire n_15488;
wire n_5300;
wire n_11393;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_16525;
wire n_7790;
wire n_16315;
wire n_19283;
wire n_6149;
wire n_17918;
wire n_7002;
wire n_12428;
wire n_3025;
wire n_1626;
wire n_15814;
wire n_1388;
wire n_10265;
wire n_16676;
wire n_18736;
wire n_15756;
wire n_19495;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_14378;
wire n_18299;
wire n_11371;
wire n_5394;
wire n_14191;
wire n_19267;
wire n_16546;
wire n_18252;
wire n_17454;
wire n_16144;
wire n_16669;
wire n_474;
wire n_6902;
wire n_3331;
wire n_10100;
wire n_18607;
wire n_5741;
wire n_15743;
wire n_2773;
wire n_7478;
wire n_19587;
wire n_19130;
wire n_5405;
wire n_7456;
wire n_13600;
wire n_964;
wire n_8503;
wire n_4756;
wire n_8196;
wire n_16062;
wire n_17712;
wire n_10846;
wire n_9787;
wire n_13363;
wire n_19648;
wire n_4970;
wire n_211;
wire n_9786;
wire n_18681;
wire n_14908;
wire n_2292;
wire n_12908;
wire n_18692;
wire n_3441;
wire n_17168;
wire n_2416;
wire n_311;
wire n_14201;
wire n_8923;
wire n_13315;
wire n_18900;
wire n_6736;
wire n_19231;
wire n_1769;
wire n_14597;
wire n_15663;
wire n_3605;
wire n_4633;
wire n_3306;
wire n_9115;
wire n_4584;
wire n_3090;
wire n_11833;
wire n_3724;
wire n_4276;
wire n_11897;
wire n_2990;
wire n_19675;
wire n_1773;
wire n_5001;
wire n_5176;
wire n_7443;
wire n_11285;
wire n_3323;
wire n_9977;
wire n_8051;
wire n_16719;
wire n_518;
wire n_9242;
wire n_4618;
wire n_4679;
wire n_914;
wire n_11262;
wire n_4496;
wire n_12880;
wire n_4805;
wire n_8651;
wire n_13959;
wire n_3454;
wire n_10732;
wire n_6885;
wire n_10851;
wire n_10221;
wire n_3547;
wire n_9299;
wire n_11162;
wire n_13685;
wire n_3816;
wire n_14693;
wire n_8842;
wire n_3214;
wire n_19780;
wire n_16915;
wire n_1917;
wire n_14486;
wire n_1580;
wire n_7730;
wire n_11592;
wire n_15090;
wire n_8467;
wire n_17043;
wire n_15385;
wire n_3109;
wire n_16094;
wire n_2863;
wire n_6417;
wire n_13281;
wire n_1731;
wire n_5648;
wire n_15627;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_10996;
wire n_858;
wire n_8676;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_17170;
wire n_19045;
wire n_410;
wire n_17351;
wire n_18060;
wire n_1594;
wire n_15048;
wire n_16393;
wire n_17135;
wire n_6199;
wire n_9823;
wire n_15739;
wire n_12937;
wire n_10698;
wire n_16891;
wire n_18118;
wire n_14665;
wire n_6726;
wire n_580;
wire n_7011;
wire n_5261;
wire n_10870;
wire n_11066;
wire n_17327;
wire n_4252;
wire n_13886;
wire n_16887;
wire n_6576;
wire n_2448;
wire n_8906;
wire n_17117;
wire n_8482;
wire n_7952;
wire n_16242;
wire n_14489;
wire n_13774;
wire n_13847;
wire n_6915;
wire n_19645;
wire n_12529;
wire n_12103;
wire n_7834;
wire n_17072;
wire n_5185;
wire n_8409;
wire n_17889;
wire n_974;
wire n_14053;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_19321;
wire n_5906;
wire n_8930;
wire n_16564;
wire n_14581;
wire n_628;
wire n_18811;
wire n_1573;
wire n_7890;
wire n_3973;
wire n_11950;
wire n_6024;
wire n_12461;
wire n_485;
wire n_11415;
wire n_7265;
wire n_7986;
wire n_17809;
wire n_2024;
wire n_17900;
wire n_202;
wire n_9879;
wire n_1749;
wire n_18744;
wire n_3474;
wire n_11390;
wire n_17238;
wire n_11669;
wire n_1669;
wire n_1024;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_8250;
wire n_10601;
wire n_9158;
wire n_18591;
wire n_1667;
wire n_16945;
wire n_9518;
wire n_7717;
wire n_18187;
wire n_18462;
wire n_18260;
wire n_5143;
wire n_11739;
wire n_10497;
wire n_14561;
wire n_18405;
wire n_1639;
wire n_13301;
wire n_8298;
wire n_466;
wire n_5215;
wire n_7860;
wire n_14212;
wire n_2548;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_13158;
wire n_1108;
wire n_11044;
wire n_15967;
wire n_15530;
wire n_1601;
wire n_11679;
wire n_8450;
wire n_17665;
wire n_3648;
wire n_17799;
wire n_7499;
wire n_3042;
wire n_19718;
wire n_7292;
wire n_12398;
wire n_17089;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_7397;
wire n_10789;
wire n_17020;
wire n_12705;
wire n_1430;
wire n_1316;
wire n_7977;
wire n_12847;
wire n_13047;
wire n_6861;
wire n_14470;
wire n_15497;
wire n_7847;
wire n_15952;
wire n_13178;
wire n_19777;
wire n_3723;
wire n_18609;
wire n_1190;
wire n_12404;
wire n_397;
wire n_11606;
wire n_5978;
wire n_11452;
wire n_15734;
wire n_6217;
wire n_5031;
wire n_10797;
wire n_7289;
wire n_17656;
wire n_14110;
wire n_14806;
wire n_1673;
wire n_7354;
wire n_18312;
wire n_13824;
wire n_3424;
wire n_239;
wire n_7960;
wire n_15620;
wire n_2326;
wire n_18053;
wire n_12912;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_2120;
wire n_16493;
wire n_6048;
wire n_6416;
wire n_2964;
wire n_352;
wire n_6838;
wire n_10068;
wire n_11988;
wire n_3485;
wire n_4077;
wire n_1361;
wire n_19034;
wire n_6256;
wire n_15645;
wire n_6613;
wire n_11438;
wire n_15965;
wire n_5221;
wire n_5641;
wire n_18877;
wire n_6361;
wire n_14981;
wire n_11348;
wire n_9685;
wire n_11685;
wire n_5731;
wire n_6678;
wire n_8662;
wire n_15058;
wire n_16539;
wire n_14971;
wire n_19801;
wire n_12429;
wire n_14734;
wire n_14494;
wire n_14956;
wire n_4623;
wire n_7325;
wire n_14866;
wire n_19123;
wire n_5007;
wire n_3320;
wire n_6370;
wire n_13743;
wire n_9923;
wire n_7166;
wire n_7356;
wire n_13378;
wire n_11319;
wire n_3476;
wire n_16981;
wire n_5629;
wire n_3439;
wire n_7873;
wire n_2688;
wire n_1489;
wire n_16418;
wire n_19363;
wire n_17795;
wire n_12640;
wire n_10063;
wire n_13092;
wire n_2852;
wire n_14292;
wire n_8419;
wire n_1496;
wire n_19497;
wire n_9862;
wire n_11385;
wire n_1485;
wire n_11355;
wire n_18659;
wire n_11674;
wire n_1846;
wire n_12535;
wire n_19031;
wire n_12327;
wire n_879;
wire n_2310;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_8430;
wire n_15719;
wire n_12058;
wire n_14879;
wire n_16143;
wire n_18387;
wire n_5852;
wire n_15164;
wire n_7052;
wire n_16755;
wire n_10496;
wire n_5960;
wire n_14149;
wire n_2454;
wire n_18225;
wire n_5321;
wire n_9960;
wire n_157;
wire n_4215;
wire n_10998;
wire n_19180;
wire n_7502;
wire n_1484;
wire n_14216;
wire n_16380;
wire n_3752;
wire n_7919;
wire n_10800;
wire n_17962;
wire n_7085;
wire n_1373;
wire n_12065;
wire n_3958;
wire n_13950;
wire n_18952;
wire n_5210;
wire n_13732;
wire n_16422;
wire n_14968;
wire n_10993;
wire n_15542;
wire n_14985;
wire n_15910;
wire n_17734;
wire n_14443;
wire n_1047;
wire n_3899;
wire n_16136;
wire n_14285;
wire n_1385;
wire n_9734;
wire n_7288;
wire n_16325;
wire n_16842;
wire n_17355;
wire n_4987;
wire n_10495;
wire n_9004;
wire n_834;
wire n_3818;
wire n_6610;
wire n_3124;
wire n_10612;
wire n_1741;
wire n_10260;
wire n_12285;
wire n_6750;
wire n_9150;
wire n_14508;
wire n_15092;
wire n_12683;
wire n_18535;
wire n_2614;
wire n_19691;
wire n_18457;
wire n_3694;
wire n_14566;
wire n_2937;
wire n_7165;
wire n_7869;
wire n_13386;
wire n_13846;
wire n_4376;
wire n_7683;
wire n_16437;
wire n_9587;
wire n_1076;
wire n_10671;
wire n_10193;
wire n_1377;
wire n_11718;
wire n_19333;
wire n_695;
wire n_14383;
wire n_16695;
wire n_4081;
wire n_11680;
wire n_14683;
wire n_18685;
wire n_17052;
wire n_7322;
wire n_17378;
wire n_11658;
wire n_12226;
wire n_13492;
wire n_14001;
wire n_5562;
wire n_15397;
wire n_978;
wire n_15840;
wire n_7880;
wire n_4382;
wire n_749;
wire n_16855;
wire n_19120;
wire n_16937;
wire n_2140;
wire n_9919;
wire n_12135;
wire n_19485;
wire n_5577;
wire n_568;
wire n_17092;
wire n_8829;
wire n_19308;
wire n_13381;
wire n_739;
wire n_5413;
wire n_8971;
wire n_18076;
wire n_16667;
wire n_1338;
wire n_16897;
wire n_10558;
wire n_9579;
wire n_9475;
wire n_17603;
wire n_15273;
wire n_573;
wire n_9049;
wire n_13718;
wire n_18701;
wire n_4480;
wire n_14775;
wire n_18809;
wire n_11045;
wire n_16756;
wire n_222;
wire n_11340;
wire n_16965;
wire n_7675;
wire n_11903;
wire n_13279;
wire n_19704;
wire n_13644;
wire n_13291;
wire n_742;
wire n_691;
wire n_10174;
wire n_377;
wire n_7524;
wire n_2935;
wire n_15897;
wire n_4046;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_12946;
wire n_16729;
wire n_18406;
wire n_13513;
wire n_4027;
wire n_12916;
wire n_1227;
wire n_3520;
wire n_8471;
wire n_12521;
wire n_18925;
wire n_9800;
wire n_11382;
wire n_19578;
wire n_10098;
wire n_11745;
wire n_1570;
wire n_15240;
wire n_1780;
wire n_15564;
wire n_1347;
wire n_17002;
wire n_14350;
wire n_7733;
wire n_17405;
wire n_18711;
wire n_4631;
wire n_19090;
wire n_1561;
wire n_13773;
wire n_14109;
wire n_6982;
wire n_2168;
wire n_5847;
wire n_7345;
wire n_17526;
wire n_14136;
wire n_7385;
wire n_10923;
wire n_5159;
wire n_2615;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_12635;
wire n_3962;
wire n_8488;
wire n_9543;
wire n_11443;
wire n_15765;
wire n_6855;
wire n_18176;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_4188;
wire n_13467;
wire n_3667;
wire n_712;
wire n_18374;
wire n_18700;
wire n_7907;
wire n_5568;
wire n_6312;
wire n_11532;
wire n_2505;
wire n_9415;
wire n_4115;
wire n_14343;
wire n_18619;
wire n_9147;
wire n_470;
wire n_11209;
wire n_3680;
wire n_15918;
wire n_5723;
wire n_5918;
wire n_16212;
wire n_11790;
wire n_1972;
wire n_19189;
wire n_4491;
wire n_19444;
wire n_363;
wire n_18148;
wire n_16313;
wire n_10420;
wire n_17058;
wire n_18309;
wire n_16363;
wire n_503;
wire n_6131;
wire n_15232;
wire n_12105;
wire n_14329;
wire n_19392;
wire n_15721;
wire n_5163;
wire n_307;
wire n_10444;
wire n_3361;
wire n_11377;
wire n_3478;
wire n_8018;
wire n_18557;
wire n_7937;
wire n_9176;
wire n_7819;
wire n_10631;
wire n_7305;
wire n_6334;
wire n_16780;
wire n_3096;
wire n_2651;
wire n_8884;
wire n_5537;
wire n_19222;
wire n_1574;
wire n_253;
wire n_2918;
wire n_8751;
wire n_4307;
wire n_11864;
wire n_11006;
wire n_15018;
wire n_6617;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_849;
wire n_4091;
wire n_14108;
wire n_1753;
wire n_3095;
wire n_15439;
wire n_16049;
wire n_2807;
wire n_8178;
wire n_14000;
wire n_14372;
wire n_3618;
wire n_4758;
wire n_17911;
wire n_12046;
wire n_10212;
wire n_18566;
wire n_5335;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_11172;
wire n_10089;
wire n_14947;
wire n_5505;
wire n_8560;
wire n_14748;
wire n_18895;
wire n_19722;
wire n_18466;
wire n_10004;
wire n_12488;
wire n_3852;
wire n_1365;
wire n_11110;
wire n_17338;
wire n_16211;
wire n_15001;
wire n_3896;
wire n_8674;
wire n_5274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_13328;
wire n_4093;
wire n_10892;
wire n_18556;
wire n_10493;
wire n_19195;
wire n_10405;
wire n_15037;
wire n_4794;
wire n_17386;
wire n_7964;
wire n_17091;
wire n_629;
wire n_14349;
wire n_6278;
wire n_7022;
wire n_12691;
wire n_11033;
wire n_19760;
wire n_19072;
wire n_18203;
wire n_14356;
wire n_19028;
wire n_5581;
wire n_16926;
wire n_16006;
wire n_992;
wire n_12651;
wire n_19194;
wire n_16476;
wire n_7486;
wire n_6756;
wire n_16373;
wire n_18792;
wire n_14190;
wire n_8563;
wire n_17223;
wire n_15546;
wire n_11534;
wire n_14157;
wire n_14344;
wire n_9221;
wire n_509;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_6411;
wire n_350;
wire n_10285;
wire n_4370;
wire n_14488;
wire n_11032;
wire n_2359;
wire n_13582;
wire n_142;
wire n_17950;
wire n_18162;
wire n_7302;
wire n_19725;
wire n_11174;
wire n_18574;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_18544;
wire n_10294;
wire n_4359;
wire n_10106;
wire n_17865;
wire n_9934;
wire n_3487;
wire n_287;
wire n_9234;
wire n_10674;
wire n_6534;
wire n_3340;
wire n_230;
wire n_5227;
wire n_16011;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_18185;
wire n_8087;
wire n_7607;
wire n_14458;
wire n_17540;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_13565;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_522;
wire n_18965;
wire n_3440;
wire n_13784;
wire n_13468;
wire n_2356;
wire n_12363;
wire n_18201;
wire n_7553;
wire n_1772;
wire n_1119;
wire n_6824;
wire n_19625;
wire n_5788;
wire n_11788;
wire n_2739;
wire n_12544;
wire n_13036;
wire n_14146;
wire n_13199;
wire n_6903;
wire n_2864;
wire n_13009;
wire n_1180;
wire n_10908;
wire n_10339;
wire n_9908;
wire n_9486;
wire n_13002;
wire n_13868;
wire n_7903;
wire n_18596;
wire n_11877;
wire n_8864;
wire n_7384;
wire n_18674;
wire n_13285;
wire n_8610;
wire n_19075;
wire n_7894;
wire n_11750;
wire n_3532;
wire n_7055;
wire n_18722;
wire n_8520;
wire n_16458;
wire n_13374;
wire n_12055;
wire n_381;
wire n_7639;
wire n_16520;
wire n_4327;
wire n_3765;
wire n_4125;
wire n_12811;
wire n_12186;
wire n_13032;
wire n_3067;
wire n_2155;
wire n_11001;
wire n_9512;
wire n_14199;
wire n_17858;
wire n_13684;
wire n_2364;
wire n_9170;
wire n_15108;
wire n_9616;
wire n_3803;
wire n_2085;
wire n_917;
wire n_16898;
wire n_3639;
wire n_9073;
wire n_12897;
wire n_5192;
wire n_18325;
wire n_12272;
wire n_9302;
wire n_19068;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_3413;
wire n_9171;
wire n_3412;
wire n_8279;
wire n_12191;
wire n_17432;
wire n_9580;
wire n_8019;
wire n_13963;
wire n_17707;
wire n_4575;
wire n_699;
wire n_4320;
wire n_18842;
wire n_7832;
wire n_9540;
wire n_17242;
wire n_11137;
wire n_451;
wire n_8390;
wire n_8898;
wire n_14316;
wire n_5231;
wire n_2190;
wire n_8613;
wire n_3438;
wire n_18300;
wire n_8464;
wire n_15701;
wire n_6423;
wire n_1441;
wire n_15612;
wire n_3373;
wire n_18804;
wire n_7441;
wire n_513;
wire n_12112;
wire n_13060;
wire n_16187;
wire n_9449;
wire n_19787;
wire n_14817;
wire n_9050;
wire n_433;
wire n_6121;
wire n_5726;
wire n_14087;
wire n_2792;
wire n_15980;
wire n_3798;
wire n_788;
wire n_329;
wire n_14438;
wire n_2674;
wire n_4641;
wire n_16253;
wire n_7133;
wire n_12202;
wire n_13836;
wire n_1866;
wire n_8661;
wire n_2130;
wire n_7424;
wire n_3714;
wire n_19774;
wire n_16671;
wire n_12870;
wire n_11156;
wire n_10611;
wire n_10715;
wire n_12333;
wire n_8609;
wire n_17666;
wire n_17219;
wire n_7626;
wire n_13576;
wire n_2714;
wire n_2245;
wire n_7310;
wire n_17451;
wire n_12119;
wire n_12618;
wire n_16093;
wire n_1265;
wire n_17266;
wire n_15129;
wire n_17146;
wire n_16209;
wire n_14306;
wire n_8873;
wire n_11891;
wire n_16276;
wire n_199;
wire n_18427;
wire n_12401;
wire n_13055;
wire n_7323;
wire n_7301;
wire n_3715;
wire n_18600;
wire n_612;
wire n_17633;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_3933;
wire n_17815;
wire n_7244;
wire n_10745;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_7633;
wire n_18760;
wire n_13937;
wire n_4146;
wire n_5711;
wire n_9437;
wire n_18724;
wire n_8640;
wire n_14359;
wire n_4855;
wire n_6186;
wire n_16933;
wire n_6803;
wire n_8437;
wire n_8427;
wire n_1188;
wire n_10605;
wire n_14013;
wire n_14419;
wire n_9933;
wire n_11449;
wire n_2916;
wire n_15251;
wire n_9892;
wire n_18976;
wire n_16727;
wire n_9462;
wire n_5972;
wire n_19447;
wire n_15854;
wire n_3145;
wire n_19438;
wire n_5444;
wire n_12501;
wire n_961;
wire n_4356;
wire n_17518;
wire n_8843;
wire n_9891;
wire n_15810;
wire n_2377;
wire n_701;
wire n_10643;
wire n_16974;
wire n_3719;
wire n_4361;
wire n_10872;
wire n_13987;
wire n_15626;
wire n_1630;
wire n_4136;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_2619;
wire n_5329;
wire n_9925;
wire n_16066;
wire n_9757;
wire n_10008;
wire n_13726;
wire n_507;
wire n_14412;
wire n_17587;
wire n_2271;
wire n_12243;
wire n_8562;
wire n_19714;
wire n_12614;
wire n_11378;
wire n_2606;
wire n_14631;
wire n_5728;
wire n_10032;
wire n_462;
wire n_304;
wire n_13425;
wire n_9806;
wire n_17105;
wire n_17233;
wire n_7021;
wire n_13591;
wire n_18296;
wire n_11713;
wire n_16972;
wire n_15586;
wire n_6355;
wire n_2954;
wire n_17821;
wire n_12931;
wire n_15525;
wire n_7215;
wire n_17790;
wire n_2493;
wire n_4802;
wire n_17566;
wire n_2705;
wire n_5523;
wire n_14332;
wire n_18379;
wire n_3405;
wire n_8016;
wire n_5423;
wire n_10645;
wire n_11096;
wire n_10604;
wire n_5074;
wire n_17398;
wire n_4044;
wire n_6564;
wire n_11161;
wire n_8709;
wire n_2631;
wire n_12491;
wire n_11216;
wire n_14368;
wire n_1293;
wire n_18390;
wire n_4701;
wire n_10966;
wire n_794;
wire n_727;
wire n_19310;
wire n_3385;
wire n_19650;
wire n_4851;
wire n_6442;
wire n_18359;
wire n_3293;
wire n_5204;
wire n_7925;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_15126;
wire n_4991;
wire n_19289;
wire n_5422;
wire n_6871;
wire n_16846;
wire n_9389;
wire n_1913;
wire n_12074;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5292;
wire n_19665;
wire n_12745;
wire n_9752;
wire n_14473;
wire n_12887;
wire n_18997;
wire n_10341;
wire n_19521;
wire n_4011;
wire n_15816;
wire n_18314;
wire n_7138;
wire n_17341;
wire n_4753;
wire n_8712;
wire n_631;
wire n_2262;
wire n_3611;
wire n_19254;
wire n_5059;
wire n_8837;
wire n_843;
wire n_17652;
wire n_2604;
wire n_14641;
wire n_16506;
wire n_17543;
wire n_15433;
wire n_15953;
wire n_5219;
wire n_9721;
wire n_11344;
wire n_3537;
wire n_12658;
wire n_1022;
wire n_9197;
wire n_19167;
wire n_1474;
wire n_14740;
wire n_9210;
wire n_6893;
wire n_5686;
wire n_8905;
wire n_13008;
wire n_18832;
wire n_18691;
wire n_7807;
wire n_18126;
wire n_14198;
wire n_14846;
wire n_3654;
wire n_1849;
wire n_9917;
wire n_12056;
wire n_14539;
wire n_8106;
wire n_4264;
wire n_12238;
wire n_5937;
wire n_19226;
wire n_12976;
wire n_14420;
wire n_18562;
wire n_6040;
wire n_11888;
wire n_13243;
wire n_14314;
wire n_16642;
wire n_14227;
wire n_10309;
wire n_11099;
wire n_5465;
wire n_8974;
wire n_4339;
wire n_14164;
wire n_3324;
wire n_10050;
wire n_9871;
wire n_19652;
wire n_1195;
wire n_10306;
wire n_7606;
wire n_1811;
wire n_7193;
wire n_3987;
wire n_1519;
wire n_18180;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_5721;
wire n_1048;
wire n_18142;
wire n_13632;
wire n_13020;
wire n_6012;
wire n_13148;
wire n_1418;
wire n_10429;
wire n_292;
wire n_11470;
wire n_3072;
wire n_13871;
wire n_4874;
wire n_4401;
wire n_889;
wire n_9903;
wire n_17208;
wire n_11102;
wire n_1110;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_17792;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_9522;
wire n_15617;
wire n_15463;
wire n_4658;
wire n_11076;
wire n_14339;
wire n_505;
wire n_1787;
wire n_16005;
wire n_6769;
wire n_9148;
wire n_11054;
wire n_2776;
wire n_10754;
wire n_5742;
wire n_3909;
wire n_9275;
wire n_10223;
wire n_1220;
wire n_8896;
wire n_19727;
wire n_7206;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_2488;
wire n_17979;
wire n_10228;
wire n_1252;
wire n_511;
wire n_8758;
wire n_6026;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_17953;
wire n_13966;
wire n_12530;
wire n_1597;
wire n_9463;
wire n_4839;
wire n_2596;
wire n_1153;
wire n_13077;
wire n_16309;
wire n_10425;
wire n_8069;
wire n_6481;
wire n_19144;
wire n_4006;
wire n_15201;
wire n_9997;
wire n_6384;
wire n_13828;
wire n_7541;
wire n_6906;
wire n_14562;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_10366;
wire n_15015;
wire n_19122;
wire n_7334;
wire n_5807;
wire n_16376;
wire n_2227;
wire n_5216;
wire n_14991;
wire n_10225;
wire n_4869;
wire n_6257;
wire n_4386;
wire n_8383;
wire n_12621;
wire n_4955;
wire n_11290;
wire n_17080;
wire n_12518;
wire n_19033;
wire n_3234;
wire n_14047;
wire n_9052;
wire n_856;
wire n_17447;
wire n_2830;
wire n_17678;
wire n_6587;
wire n_7781;
wire n_7360;
wire n_14568;
wire n_2181;
wire n_11702;
wire n_19395;
wire n_16970;
wire n_11372;
wire n_2826;
wire n_10817;
wire n_15324;
wire n_326;
wire n_8355;
wire n_19501;
wire n_17098;
wire n_12741;
wire n_18041;
wire n_7101;
wire n_1635;
wire n_7530;
wire n_15006;
wire n_15619;
wire n_18911;
wire n_9860;
wire n_12510;
wire n_11756;
wire n_2851;
wire n_8369;
wire n_9022;
wire n_160;
wire n_9103;
wire n_17142;
wire n_8831;
wire n_1508;
wire n_5608;
wire n_2240;
wire n_392;
wire n_12233;
wire n_8853;
wire n_4582;
wire n_6252;
wire n_18403;
wire n_6211;
wire n_15716;
wire n_5844;
wire n_17499;
wire n_1549;
wire n_17898;
wire n_17172;
wire n_8081;
wire n_16608;
wire n_17310;
wire n_13442;
wire n_1916;
wire n_14444;
wire n_18531;
wire n_10484;
wire n_11744;
wire n_17247;
wire n_10288;
wire n_18838;
wire n_10388;
wire n_6189;
wire n_15299;
wire n_4016;
wire n_11072;
wire n_621;
wire n_750;
wire n_2823;
wire n_5597;
wire n_13944;
wire n_9492;
wire n_6413;
wire n_7419;
wire n_6506;
wire n_18476;
wire n_1997;
wire n_710;
wire n_1818;
wire n_17086;
wire n_6935;
wire n_9727;
wire n_13019;
wire n_12703;
wire n_13079;
wire n_4397;
wire n_18343;
wire n_5050;
wire n_746;
wire n_3416;
wire n_3498;
wire n_15369;
wire n_15134;
wire n_16110;
wire n_2957;
wire n_1740;
wire n_19420;
wire n_9375;
wire n_17715;
wire n_5980;
wire n_8770;
wire n_3672;
wire n_15453;
wire n_5318;
wire n_6105;
wire n_6022;
wire n_10964;
wire n_3382;
wire n_19739;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_5053;
wire n_9458;
wire n_7841;
wire n_8466;
wire n_6527;
wire n_15275;
wire n_19092;
wire n_8094;
wire n_4824;
wire n_2037;
wire n_4567;
wire n_6430;
wire n_782;
wire n_18268;
wire n_809;
wire n_10987;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_1797;
wire n_4595;
wire n_402;
wire n_1870;
wire n_11965;
wire n_4904;
wire n_1152;
wire n_14696;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_711;
wire n_3105;
wire n_14006;
wire n_6666;
wire n_3692;
wire n_8321;
wire n_19116;
wire n_9954;
wire n_8735;
wire n_1695;
wire n_11722;
wire n_2272;
wire n_2760;
wire n_972;
wire n_12310;
wire n_5348;
wire n_6594;
wire n_624;
wire n_19471;
wire n_7095;
wire n_3045;
wire n_16672;
wire n_11701;
wire n_885;
wire n_3666;
wire n_4916;
wire n_18010;
wire n_13917;
wire n_7184;
wire n_9617;
wire n_13546;
wire n_14595;
wire n_17001;
wire n_7908;
wire n_7974;
wire n_7551;
wire n_11980;
wire n_11255;
wire n_13592;
wire n_3858;
wire n_17224;
wire n_11720;
wire n_3502;
wire n_5461;
wire n_13874;
wire n_6482;
wire n_5147;
wire n_15506;
wire n_1355;
wire n_9810;
wire n_14469;
wire n_16201;
wire n_2562;
wire n_17690;
wire n_1522;
wire n_5755;
wire n_8043;
wire n_16377;
wire n_14492;
wire n_1548;
wire n_1155;
wire n_14134;
wire n_4944;
wire n_11990;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_15457;
wire n_14345;
wire n_16847;
wire n_6841;
wire n_10153;
wire n_17622;
wire n_17952;
wire n_5054;
wire n_2962;
wire n_8171;
wire n_9006;
wire n_19641;
wire n_6774;
wire n_16964;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_14816;
wire n_8710;
wire n_12806;
wire n_4045;
wire n_14302;
wire n_8549;
wire n_10172;
wire n_8054;
wire n_13904;
wire n_16614;
wire n_3258;
wire n_18694;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_17045;
wire n_15784;
wire n_18613;
wire n_3149;
wire n_11969;
wire n_7914;
wire n_16388;
wire n_3365;
wire n_6521;
wire n_3379;
wire n_8857;
wire n_14243;
wire n_9040;
wire n_6162;
wire n_8010;
wire n_3939;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_1650;
wire n_13574;
wire n_12762;
wire n_16740;
wire n_9830;
wire n_18870;
wire n_10761;
wire n_2761;
wire n_3776;
wire n_18781;
wire n_11579;
wire n_1019;
wire n_15303;
wire n_8291;
wire n_18017;
wire n_4170;
wire n_11535;
wire n_2845;
wire n_18400;
wire n_5173;
wire n_12975;
wire n_16291;
wire n_13850;
wire n_6740;
wire n_1113;
wire n_11510;
wire n_6315;
wire n_17866;
wire n_12736;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_9163;
wire n_15461;
wire n_6910;
wire n_6262;
wire n_14800;
wire n_2827;
wire n_7703;
wire n_6319;
wire n_17352;
wire n_14888;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_1879;
wire n_6536;
wire n_256;
wire n_6175;
wire n_7040;
wire n_8280;
wire n_12390;
wire n_367;
wire n_18898;
wire n_2569;
wire n_10235;
wire n_6978;
wire n_5351;
wire n_12805;
wire n_6093;
wire n_11649;
wire n_16306;
wire n_703;
wire n_18485;
wire n_9190;
wire n_6947;
wire n_14918;
wire n_5293;
wire n_8203;
wire n_6099;
wire n_1324;
wire n_1435;
wire n_3920;
wire n_4892;
wire n_6140;
wire n_15489;
wire n_12914;
wire n_17159;
wire n_17721;
wire n_9506;
wire n_18440;
wire n_6415;
wire n_4439;
wire n_18883;
wire n_16542;
wire n_15158;
wire n_10828;
wire n_18866;
wire n_12300;
wire n_15389;
wire n_7549;
wire n_17308;
wire n_17425;
wire n_11281;
wire n_13056;
wire n_16019;
wire n_17732;
wire n_12337;
wire n_18520;
wire n_13466;
wire n_15082;
wire n_8871;
wire n_11114;
wire n_19442;
wire n_8418;
wire n_7740;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_10860;
wire n_18259;
wire n_17517;
wire n_4930;
wire n_16208;
wire n_19327;
wire n_15209;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_12712;
wire n_360;
wire n_2149;
wire n_15078;
wire n_4557;
wire n_13012;
wire n_895;
wire n_8924;
wire n_12752;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_15511;
wire n_4593;
wire n_4465;
wire n_3622;
wire n_19600;
wire n_18204;
wire n_4495;
wire n_14278;
wire n_5117;
wire n_8214;
wire n_12777;
wire n_14706;
wire n_5990;
wire n_7043;
wire n_11462;
wire n_11732;
wire n_5024;
wire n_4559;
wire n_18137;
wire n_12819;
wire n_10214;
wire n_8241;
wire n_838;
wire n_3336;
wire n_8442;
wire n_2952;
wire n_9572;
wire n_15282;
wire n_9229;
wire n_19505;
wire n_16812;
wire n_16038;
wire n_12237;
wire n_18350;
wire n_6134;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_13372;
wire n_2430;
wire n_653;
wire n_11375;
wire n_11267;
wire n_9602;
wire n_9311;
wire n_4335;
wire n_19482;
wire n_2034;
wire n_576;
wire n_6593;
wire n_8630;
wire n_2683;
wire n_19432;
wire n_9884;
wire n_9876;
wire n_9260;
wire n_14534;
wire n_13630;
wire n_16535;
wire n_13700;
wire n_10406;
wire n_3204;
wire n_17859;
wire n_6746;
wire n_11985;
wire n_8447;
wire n_6443;
wire n_14290;
wire n_7980;
wire n_348;
wire n_8828;
wire n_18631;
wire n_17687;
wire n_390;
wire n_1148;
wire n_6749;
wire n_10798;
wire n_10965;
wire n_19657;
wire n_7732;
wire n_13325;
wire n_14850;
wire n_15135;
wire n_16196;
wire n_11911;
wire n_4265;
wire n_11442;
wire n_2950;
wire n_5634;
wire n_719;
wire n_18862;
wire n_14064;
wire n_14524;
wire n_1090;
wire n_8859;
wire n_16883;
wire n_11388;
wire n_11651;
wire n_1362;
wire n_17946;
wire n_10154;
wire n_18663;
wire n_7922;
wire n_17469;
wire n_15826;
wire n_5580;
wire n_1450;
wire n_19101;
wire n_10033;
wire n_1789;
wire n_17877;
wire n_8311;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_9877;
wire n_8764;
wire n_19361;
wire n_16167;
wire n_2161;
wire n_19452;
wire n_12990;
wire n_14246;
wire n_5764;
wire n_6920;
wire n_11817;
wire n_8729;
wire n_10359;
wire n_3344;
wire n_2334;
wire n_14957;
wire n_5133;
wire n_1763;
wire n_13447;
wire n_6907;
wire n_7144;
wire n_16579;
wire n_11479;
wire n_11737;
wire n_8048;
wire n_635;
wire n_12028;
wire n_3786;
wire n_7072;
wire n_13095;
wire n_4254;
wire n_8253;
wire n_4303;
wire n_18592;
wire n_15032;
wire n_1158;
wire n_11600;
wire n_2248;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_10722;
wire n_8088;
wire n_17855;
wire n_10666;
wire n_3147;
wire n_15440;
wire n_753;
wire n_3925;
wire n_3180;
wire n_8516;
wire n_8302;
wire n_17717;
wire n_15610;
wire n_359;
wire n_15329;
wire n_8167;
wire n_7859;
wire n_14315;
wire n_7872;
wire n_1479;
wire n_4768;
wire n_13858;
wire n_17913;
wire n_3717;
wire n_7480;
wire n_5410;
wire n_571;
wire n_2215;
wire n_16255;
wire n_8944;
wire n_1884;
wire n_10023;
wire n_10999;
wire n_665;
wire n_5156;
wire n_18716;
wire n_10410;
wire n_19732;
wire n_4447;
wire n_3445;
wire n_373;
wire n_16983;
wire n_8975;
wire n_1833;
wire n_17009;
wire n_11305;
wire n_17668;
wire n_9101;
wire n_15631;
wire n_14755;
wire n_8825;
wire n_12969;
wire n_1856;
wire n_12260;
wire n_12016;
wire n_8266;
wire n_5691;
wire n_8981;
wire n_4957;
wire n_17082;
wire n_165;
wire n_8771;
wire n_15750;
wire n_4039;
wire n_457;
wire n_3800;
wire n_4566;
wire n_12939;
wire n_15038;
wire n_17925;
wire n_10404;
wire n_8138;
wire n_6638;
wire n_12779;
wire n_17505;
wire n_17199;
wire n_2930;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_9211;
wire n_8124;
wire n_9395;
wire n_7366;
wire n_5269;
wire n_17348;
wire n_1538;
wire n_8147;
wire n_5468;
wire n_4730;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_10700;
wire n_17743;
wire n_10968;
wire n_3579;
wire n_14247;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_700;
wire n_3178;
wire n_16155;
wire n_15418;
wire n_5256;
wire n_11970;
wire n_7918;
wire n_4168;
wire n_6651;
wire n_12308;
wire n_1923;
wire n_10783;
wire n_12163;
wire n_3952;
wire n_11523;
wire n_12944;
wire n_3911;
wire n_7472;
wire n_9737;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_10812;
wire n_14709;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_2997;
wire n_10001;
wire n_13280;
wire n_12145;
wire n_11088;
wire n_5939;
wire n_5509;
wire n_8160;
wire n_3619;
wire n_11405;
wire n_19274;
wire n_1786;
wire n_13103;
wire n_18385;
wire n_15630;
wire n_4198;
wire n_1371;
wire n_10977;
wire n_2886;
wire n_11299;
wire n_10615;
wire n_1803;
wire n_11542;
wire n_4065;
wire n_229;
wire n_7647;
wire n_12426;
wire n_16222;
wire n_15068;
wire n_15442;
wire n_9054;
wire n_2470;
wire n_4446;
wire n_10532;
wire n_17776;
wire n_4417;
wire n_13995;
wire n_13073;
wire n_6728;
wire n_2286;
wire n_4743;
wire n_16029;
wire n_2018;
wire n_1903;
wire n_13556;
wire n_13367;
wire n_10771;
wire n_11441;
wire n_14203;
wire n_17269;
wire n_693;
wire n_1056;
wire n_19802;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_5110;
wire n_10104;
wire n_772;
wire n_2806;
wire n_9117;
wire n_19426;
wire n_3028;
wire n_9381;
wire n_3076;
wire n_12049;
wire n_14498;
wire n_886;
wire n_343;
wire n_3624;
wire n_1820;
wire n_6549;
wire n_539;
wire n_19708;
wire n_6096;
wire n_7853;
wire n_12526;
wire n_2836;
wire n_8890;
wire n_16575;
wire n_7721;
wire n_7192;
wire n_19602;
wire n_11206;
wire n_11593;
wire n_15807;
wire n_3906;
wire n_11786;
wire n_12737;
wire n_4954;
wire n_17258;
wire n_15113;
wire n_9273;
wire n_2612;
wire n_8970;
wire n_16910;
wire n_2591;
wire n_1815;
wire n_10640;
wire n_2593;
wire n_10729;
wire n_14656;
wire n_16052;
wire n_14745;
wire n_19243;
wire n_4605;
wire n_7635;
wire n_19712;
wire n_11268;
wire n_17121;
wire n_14760;
wire n_3943;
wire n_11501;
wire n_7227;
wire n_13390;
wire n_8030;
wire n_6052;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_12010;
wire n_1843;
wire n_9738;
wire n_12026;
wire n_4227;
wire n_521;
wire n_17481;
wire n_8633;
wire n_17645;
wire n_7689;
wire n_6511;
wire n_18470;
wire n_1309;
wire n_916;
wire n_4415;
wire n_7099;
wire n_1970;
wire n_14676;
wire n_6358;
wire n_2059;
wire n_2669;
wire n_18880;
wire n_11313;
wire n_10438;
wire n_6986;
wire n_8801;
wire n_3912;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_16438;
wire n_860;
wire n_8219;
wire n_15373;
wire n_18580;
wire n_1302;
wire n_10575;
wire n_11028;
wire n_12171;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_15211;
wire n_10760;
wire n_4792;
wire n_15334;
wire n_7731;
wire n_11527;
wire n_18404;
wire n_3514;
wire n_16486;
wire n_9535;
wire n_2654;
wire n_5302;
wire n_966;
wire n_12490;
wire n_3357;
wire n_692;
wire n_5781;
wire n_3895;
wire n_8486;
wire n_12829;
wire n_4118;
wire n_2176;
wire n_2459;
wire n_18662;
wire n_1111;
wire n_1251;
wire n_11610;
wire n_12739;
wire n_7132;
wire n_2711;
wire n_17021;
wire n_17710;
wire n_6663;
wire n_12609;
wire n_4441;
wire n_18248;
wire n_8155;
wire n_11360;
wire n_11868;
wire n_1664;
wire n_3022;
wire n_8098;
wire n_9191;
wire n_17791;
wire n_5654;
wire n_2345;
wire n_18202;
wire n_6376;
wire n_18141;
wire n_5113;
wire n_12888;
wire n_5479;
wire n_19407;
wire n_8485;
wire n_14852;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_13070;
wire n_850;
wire n_5692;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_14491;
wire n_15011;
wire n_17607;
wire n_3768;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_9664;
wire n_3785;
wire n_14928;
wire n_2602;
wire n_2980;
wire n_13778;
wire n_696;
wire n_9931;
wire n_16470;
wire n_16419;
wire n_1082;
wire n_1317;
wire n_16956;
wire n_3227;
wire n_4055;
wire n_14634;
wire n_2178;
wire n_10753;
wire n_13174;
wire n_7108;
wire n_14455;
wire n_1796;
wire n_17164;
wire n_11879;
wire n_2082;
wire n_7876;
wire n_17175;
wire n_9656;
wire n_3707;
wire n_8148;
wire n_8150;
wire n_3578;
wire n_909;
wire n_12596;
wire n_15398;
wire n_15593;
wire n_18175;
wire n_4925;
wire n_16424;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_19367;
wire n_12697;
wire n_7260;
wire n_6409;
wire n_11939;
wire n_1634;
wire n_3252;
wire n_627;
wire n_14347;
wire n_7552;
wire n_19052;
wire n_17969;
wire n_12166;
wire n_2133;
wire n_1712;
wire n_1523;
wire n_10646;
wire n_15725;
wire n_1627;
wire n_11704;
wire n_17506;
wire n_18050;
wire n_8763;
wire n_5208;
wire n_8679;
wire n_7239;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_7050;
wire n_17137;
wire n_2573;
wire n_2646;
wire n_6623;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_16924;
wire n_1364;
wire n_13316;
wire n_10313;
wire n_13689;
wire n_8139;
wire n_17268;
wire n_18000;
wire n_19384;
wire n_3037;
wire n_19288;
wire n_3729;
wire n_19431;
wire n_10773;
wire n_18210;
wire n_2537;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_14836;
wire n_12867;
wire n_4988;
wire n_15960;
wire n_15343;
wire n_7568;
wire n_6354;
wire n_6344;
wire n_12123;
wire n_9772;
wire n_18885;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_15370;
wire n_7724;
wire n_18001;
wire n_4284;
wire n_6305;
wire n_1947;
wire n_12547;
wire n_16148;
wire n_15577;
wire n_3426;
wire n_16550;
wire n_4971;
wire n_19066;
wire n_5857;
wire n_8646;
wire n_13415;
wire n_10259;
wire n_7107;
wire n_17111;
wire n_6457;
wire n_17951;
wire n_8597;
wire n_17379;
wire n_987;
wire n_7123;
wire n_5499;
wire n_720;
wire n_8117;
wire n_15169;
wire n_1707;
wire n_10213;
wire n_13888;
wire n_16592;
wire n_8208;
wire n_797;
wire n_2933;
wire n_19373;
wire n_1878;
wire n_8536;
wire n_17252;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_16475;
wire n_5190;
wire n_13892;
wire n_16361;
wire n_14559;
wire n_16831;
wire n_4097;
wire n_1666;
wire n_19696;
wire n_5392;
wire n_17110;
wire n_14052;
wire n_14311;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_11874;
wire n_13926;
wire n_10171;
wire n_15184;
wire n_1228;
wire n_5455;
wire n_18131;
wire n_5442;
wire n_6386;
wire n_12803;
wire n_5948;
wire n_19518;
wire n_5511;
wire n_2898;
wire n_6208;
wire n_6739;
wire n_15779;
wire n_8202;
wire n_15366;
wire n_3200;
wire n_12734;
wire n_3167;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_10269;
wire n_19504;
wire n_12262;
wire n_14910;
wire n_14385;
wire n_14499;
wire n_8738;
wire n_9126;
wire n_15368;
wire n_19077;
wire n_11376;
wire n_9438;
wire n_18433;
wire n_7808;
wire n_6544;
wire n_9122;
wire n_14731;
wire n_683;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_16337;
wire n_17691;
wire n_8721;
wire n_12820;
wire n_9912;
wire n_6356;
wire n_13558;
wire n_3577;
wire n_2432;
wire n_10148;
wire n_19491;
wire n_1363;
wire n_3641;
wire n_2218;
wire n_16890;
wire n_13890;
wire n_5481;
wire n_9264;
wire n_14483;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_15724;
wire n_19303;
wire n_4053;
wire n_10234;
wire n_8836;
wire n_7019;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_13521;
wire n_4167;
wire n_19788;
wire n_14926;
wire n_10731;
wire n_9878;
wire n_14591;
wire n_14363;
wire n_14576;
wire n_4431;
wire n_17797;
wire n_1125;
wire n_11498;
wire n_10513;
wire n_441;
wire n_7296;
wire n_4299;
wire n_7575;
wire n_3571;
wire n_7083;
wire n_1775;
wire n_7720;
wire n_11643;
wire n_1093;
wire n_6268;
wire n_5827;
wire n_5199;
wire n_11103;
wire n_6456;
wire n_16823;
wire n_16966;
wire n_14088;
wire n_5313;
wire n_17926;
wire n_13817;
wire n_3856;
wire n_9971;
wire n_19579;
wire n_3425;
wire n_10894;
wire n_14118;
wire n_18082;
wire n_9524;
wire n_6467;
wire n_9243;
wire n_9282;
wire n_1453;
wire n_6796;
wire n_18821;
wire n_12417;
wire n_4830;
wire n_13225;
wire n_17006;
wire n_1224;
wire n_10208;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_10804;
wire n_6486;
wire n_3960;
wire n_17246;
wire n_17167;
wire n_18357;
wire n_8438;
wire n_13355;
wire n_18160;
wire n_4693;
wire n_18614;
wire n_10793;
wire n_2000;
wire n_14672;
wire n_4267;
wire n_15127;
wire n_6732;
wire n_2270;
wire n_12711;
wire n_12219;
wire n_906;
wire n_10440;
wire n_1733;
wire n_9695;
wire n_11306;
wire n_19169;
wire n_4609;
wire n_1687;
wire n_8757;
wire n_2328;
wire n_13035;
wire n_7020;
wire n_13021;
wire n_613;
wire n_12893;
wire n_8596;
wire n_3314;
wire n_3016;
wire n_11292;
wire n_554;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_5474;
wire n_12289;
wire n_10813;
wire n_1889;
wire n_10757;
wire n_13046;
wire n_13935;
wire n_435;
wire n_16670;
wire n_762;
wire n_11431;
wire n_1778;
wire n_5287;
wire n_13646;
wire n_1079;
wire n_5083;
wire n_6007;
wire n_3338;
wire n_18186;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_8834;
wire n_3636;
wire n_2327;
wire n_16429;
wire n_15262;
wire n_10822;
wire n_18773;
wire n_7104;
wire n_7467;
wire n_14609;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_13380;
wire n_5771;
wire n_17369;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_11836;
wire n_349;
wire n_6602;
wire n_10924;
wire n_17421;
wire n_11186;
wire n_9742;
wire n_6484;
wire n_19642;
wire n_3637;
wire n_12527;
wire n_4574;
wire n_19800;
wire n_1859;
wire n_9019;
wire n_13891;
wire n_1718;
wire n_8985;
wire n_7692;
wire n_19463;
wire n_12477;
wire n_4234;
wire n_14325;
wire n_15503;
wire n_10418;
wire n_1768;
wire n_19589;
wire n_3974;
wire n_10875;
wire n_1847;
wire n_3634;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_11846;
wire n_1397;
wire n_12400;
wire n_901;
wire n_2755;
wire n_4660;
wire n_1623;
wire n_16861;
wire n_9145;
wire n_12092;
wire n_3112;
wire n_12295;
wire n_9754;
wire n_19549;
wire n_9315;
wire n_18483;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_6734;
wire n_7476;
wire n_5570;
wire n_18096;
wire n_785;
wire n_7495;
wire n_7392;
wire n_5435;
wire n_9765;
wire n_3213;
wire n_3820;
wire n_5200;
wire n_6941;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_8680;
wire n_2722;
wire n_4152;
wire n_16522;
wire n_10394;
wire n_11391;
wire n_15462;
wire n_5244;
wire n_12714;
wire n_16779;
wire n_5889;
wire n_19024;
wire n_5391;
wire n_1938;
wire n_9763;
wire n_11070;
wire n_13337;
wire n_15112;
wire n_18146;
wire n_3394;
wire n_9162;
wire n_1715;
wire n_14849;
wire n_1443;
wire n_1272;
wire n_16661;
wire n_5849;
wire n_11648;
wire n_4554;
wire n_19044;
wire n_10322;
wire n_7135;
wire n_8555;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_15912;
wire n_16206;
wire n_8508;
wire n_19509;
wire n_18827;
wire n_16529;
wire n_1705;
wire n_3905;
wire n_8207;
wire n_11653;
wire n_4680;
wire n_3013;
wire n_11717;
wire n_15246;
wire n_14940;
wire n_6165;
wire n_19153;
wire n_17553;
wire n_15395;
wire n_12838;
wire n_2670;
wire n_18813;
wire n_13505;
wire n_5910;
wire n_12776;
wire n_1569;
wire n_7033;
wire n_13156;
wire n_15529;
wire n_10710;
wire n_5557;
wire n_411;
wire n_8850;
wire n_14647;
wire n_18384;
wire n_8002;
wire n_19610;
wire n_1795;
wire n_16722;
wire n_9090;
wire n_16412;
wire n_12008;
wire n_6119;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_9261;
wire n_8301;
wire n_17453;
wire n_12223;
wire n_18706;
wire n_16758;
wire n_548;
wire n_10942;
wire n_11430;
wire n_13010;
wire n_19073;
wire n_345;
wire n_11239;
wire n_4943;
wire n_10953;
wire n_7842;
wire n_2629;
wire n_2172;
wire n_6202;
wire n_17831;
wire n_12898;
wire n_4682;
wire n_19523;
wire n_15540;
wire n_10343;
wire n_4942;
wire n_9258;
wire n_1086;
wire n_10286;
wire n_10371;
wire n_14990;
wire n_2561;
wire n_16691;
wire n_7236;
wire n_10257;
wire n_3305;
wire n_11219;
wire n_10047;
wire n_14541;
wire n_3267;
wire n_16186;
wire n_1914;
wire n_1318;
wire n_13766;
wire n_11226;
wire n_3005;
wire n_16989;
wire n_11413;
wire n_4840;
wire n_1029;
wire n_16617;
wire n_5320;
wire n_5353;
wire n_13710;
wire n_11232;
wire n_2417;
wire n_9105;
wire n_12080;
wire n_16261;
wire n_5093;
wire n_1556;
wire n_19512;
wire n_5979;
wire n_9668;
wire n_13335;
wire n_14022;
wire n_2083;
wire n_5517;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_3401;
wire n_10744;
wire n_3242;
wire n_9870;
wire n_3613;
wire n_11334;
wire n_7678;
wire n_1045;
wire n_13075;
wire n_13736;
wire n_13129;
wire n_9178;
wire n_6063;
wire n_16118;
wire n_1325;
wire n_6504;
wire n_2923;
wire n_1727;
wire n_13586;
wire n_15813;
wire n_10597;
wire n_17382;
wire n_16281;
wire n_11827;
wire n_13049;
wire n_13961;
wire n_17413;
wire n_15745;
wire n_3814;
wire n_6003;
wire n_6684;
wire n_19084;
wire n_13063;
wire n_5451;
wire n_9323;
wire n_19728;
wire n_6961;
wire n_3543;
wire n_13252;
wire n_9922;
wire n_12024;
wire n_13084;
wire n_2903;
wire n_16622;
wire n_15374;
wire n_3808;
wire n_4365;
wire n_18123;
wire n_16440;
wire n_7929;
wire n_16821;
wire n_10572;
wire n_16431;
wire n_1007;
wire n_1929;
wire n_19272;
wire n_1592;
wire n_19455;
wire n_13985;
wire n_3758;
wire n_17594;
wire n_14124;
wire n_19119;
wire n_17658;
wire n_13552;
wire n_18086;
wire n_12681;
wire n_3343;
wire n_18419;
wire n_13022;
wire n_18583;
wire n_2752;
wire n_17047;
wire n_9513;
wire n_16447;
wire n_16124;
wire n_4885;
wire n_15446;
wire n_10555;
wire n_19179;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_13656;
wire n_18967;
wire n_3658;
wire n_6834;
wire n_6817;
wire n_6927;
wire n_5209;
wire n_16841;
wire n_15470;
wire n_6215;
wire n_4212;
wire n_5699;
wire n_181;
wire n_5765;
wire n_15754;
wire n_17375;
wire n_7862;
wire n_16708;
wire n_17439;
wire n_10630;
wire n_17955;
wire n_8808;
wire n_10061;
wire n_300;
wire n_15599;
wire n_11865;
wire n_13024;
wire n_10694;
wire n_11041;
wire n_14490;
wire n_9708;
wire n_5064;
wire n_15479;
wire n_7119;
wire n_8889;
wire n_601;
wire n_13986;
wire n_9790;
wire n_11973;
wire n_5759;
wire n_13329;
wire n_7874;
wire n_8490;
wire n_10329;
wire n_9979;
wire n_8767;
wire n_13946;
wire n_9505;
wire n_2566;
wire n_15028;
wire n_2702;
wire n_7420;
wire n_7102;
wire n_13618;
wire n_4568;
wire n_10662;
wire n_5559;
wire n_18653;
wire n_17534;
wire n_14993;
wire n_14327;
wire n_8624;
wire n_11022;
wire n_10247;
wire n_5377;
wire n_1016;
wire n_8796;
wire n_4106;
wire n_1501;
wire n_17829;
wire n_10733;
wire n_10472;
wire n_12597;
wire n_13744;
wire n_12834;
wire n_10066;
wire n_17239;
wire n_14335;
wire n_6419;
wire n_3553;
wire n_18989;
wire n_2275;
wire n_15087;
wire n_2568;
wire n_2022;
wire n_3494;
wire n_6244;
wire n_6900;
wire n_9337;
wire n_15219;
wire n_908;
wire n_9432;
wire n_17295;
wire n_19563;
wire n_7705;
wire n_2106;
wire n_5350;
wire n_5470;
wire n_18331;
wire n_7932;
wire n_7058;
wire n_15009;
wire n_8262;
wire n_5700;
wire n_9874;
wire n_7981;
wire n_12588;
wire n_17203;
wire n_15648;
wire n_17548;
wire n_5874;
wire n_9231;
wire n_3328;
wire n_18612;
wire n_7973;
wire n_6815;
wire n_15634;
wire n_9569;
wire n_14823;
wire n_14691;
wire n_2530;
wire n_16908;
wire n_16508;
wire n_9719;
wire n_8358;
wire n_9552;
wire n_13822;
wire n_14948;
wire n_6317;
wire n_475;
wire n_492;
wire n_4012;
wire n_10756;
wire n_3645;
wire n_17099;
wire n_14387;
wire n_16572;
wire n_11797;
wire n_18933;
wire n_18889;
wire n_14106;
wire n_18788;
wire n_13616;
wire n_18667;
wire n_7820;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_15468;
wire n_9633;
wire n_3422;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_13627;
wire n_878;
wire n_19040;
wire n_5120;
wire n_13112;
wire n_10042;
wire n_10478;
wire n_16581;
wire n_981;
wire n_18597;
wire n_13163;
wire n_3702;
wire n_8754;
wire n_9847;
wire n_16968;
wire n_2233;
wire n_18098;
wire n_10367;
wire n_3233;
wire n_10867;
wire n_3310;
wire n_4061;
wire n_7460;
wire n_9519;
wire n_19735;
wire n_14814;
wire n_6367;
wire n_13564;
wire n_12671;
wire n_8714;
wire n_13260;
wire n_17302;
wire n_10085;
wire n_1051;
wire n_8182;
wire n_16165;
wire n_14090;
wire n_6056;
wire n_7200;
wire n_3206;
wire n_2363;
wire n_553;
wire n_15424;
wire n_4903;
wire n_17301;
wire n_15554;
wire n_15836;
wire n_15966;
wire n_16009;
wire n_15309;
wire n_14463;
wire n_2540;
wire n_973;
wire n_5743;
wire n_13503;
wire n_11152;
wire n_16318;
wire n_14166;
wire n_4522;
wire n_10122;
wire n_679;
wire n_9327;
wire n_16175;
wire n_5368;
wire n_4263;
wire n_14271;
wire n_7059;
wire n_915;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_11964;
wire n_3155;
wire n_7826;
wire n_19078;
wire n_5933;
wire n_7076;
wire n_4780;
wire n_11403;
wire n_2697;
wire n_6866;
wire n_17108;
wire n_2512;
wire n_9387;
wire n_3039;
wire n_14596;
wire n_6514;
wire n_9794;
wire n_1322;
wire n_16387;
wire n_11142;
wire n_1958;
wire n_17434;
wire n_1197;
wire n_17509;
wire n_4984;
wire n_3420;
wire n_10862;
wire n_4283;
wire n_8911;
wire n_900;
wire n_8248;
wire n_11476;
wire n_2659;
wire n_13633;
wire n_14538;
wire n_2116;
wire n_19534;
wire n_1013;
wire n_17999;
wire n_11367;
wire n_15478;
wire n_2183;
wire n_16797;
wire n_12676;
wire n_18755;
wire n_3392;
wire n_13913;
wire n_19166;
wire n_8733;
wire n_6050;
wire n_7976;
wire n_13080;
wire n_13403;
wire n_17444;
wire n_1581;
wire n_1357;
wire n_14952;
wire n_1853;
wire n_10386;
wire n_12128;
wire n_14060;
wire n_14018;
wire n_15959;
wire n_5563;
wire n_1348;
wire n_11026;
wire n_13309;
wire n_15292;
wire n_11467;
wire n_12672;
wire n_12063;
wire n_8330;
wire n_1009;
wire n_15560;
wire n_1160;
wire n_15065;
wire n_5717;
wire n_1247;
wire n_9696;
wire n_6017;
wire n_15771;
wire n_15508;
wire n_471;
wire n_17990;
wire n_14148;
wire n_5720;
wire n_4702;
wire n_4895;
wire n_12924;
wire n_16331;
wire n_12732;
wire n_17171;
wire n_12649;
wire n_5898;
wire n_17458;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_12843;
wire n_14279;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_17856;
wire n_2365;
wire n_19573;
wire n_15687;
wire n_8540;
wire n_2447;
wire n_11248;
wire n_9915;
wire n_5940;
wire n_6089;
wire n_7588;
wire n_18480;
wire n_4969;
wire n_10017;
wire n_11141;
wire n_5105;
wire n_11093;
wire n_19556;
wire n_17716;
wire n_5263;
wire n_2510;
wire n_6713;
wire n_18750;
wire n_15968;
wire n_17893;
wire n_4602;
wire n_13181;
wire n_18303;
wire n_1163;
wire n_16487;
wire n_17592;
wire n_15047;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_7593;
wire n_17156;
wire n_17908;
wire n_14085;
wire n_8068;
wire n_19599;
wire n_2173;
wire n_7764;
wire n_19634;
wire n_10196;
wire n_493;
wire n_14573;
wire n_17433;
wire n_19453;
wire n_2108;
wire n_8693;
wire n_6454;
wire n_12625;
wire n_12177;
wire n_7307;
wire n_14512;
wire n_1280;
wire n_6918;
wire n_16214;
wire n_13761;
wire n_19576;
wire n_3296;
wire n_19065;
wire n_16219;
wire n_17017;
wire n_14456;
wire n_13364;
wire n_11494;
wire n_14743;
wire n_10218;
wire n_18492;
wire n_3792;
wire n_4791;
wire n_19127;
wire n_14859;
wire n_8062;
wire n_11832;
wire n_6375;
wire n_12974;
wire n_13078;
wire n_1956;
wire n_7047;
wire n_6632;
wire n_4549;
wire n_17241;
wire n_15795;
wire n_10542;
wire n_16814;
wire n_4349;
wire n_10681;
wire n_15162;
wire n_9732;
wire n_16494;
wire n_13370;
wire n_11894;
wire n_10222;
wire n_10524;
wire n_6705;
wire n_17988;
wire n_8629;
wire n_818;
wire n_9517;
wire n_15237;
wire n_15862;
wire n_6591;
wire n_2207;
wire n_13643;
wire n_9780;
wire n_3482;
wire n_2198;
wire n_13607;
wire n_6289;
wire n_3272;
wire n_8524;
wire n_19355;
wire n_18907;
wire n_4393;
wire n_14114;
wire n_1068;
wire n_932;
wire n_14904;
wire n_3978;
wire n_3317;
wire n_5560;
wire n_6512;
wire n_4074;
wire n_4918;
wire n_13820;
wire n_4013;
wire n_6703;
wire n_12122;
wire n_13428;
wire n_354;
wire n_17958;
wire n_19667;
wire n_2941;
wire n_547;
wire n_17194;
wire n_19686;
wire n_6086;
wire n_16668;
wire n_4147;
wire n_4477;
wire n_18139;
wire n_3168;
wire n_12184;
wire n_10210;
wire n_1793;
wire n_5611;
wire n_12571;
wire n_6219;
wire n_11853;
wire n_19626;
wire n_16770;
wire n_4742;
wire n_9609;
wire n_10029;
wire n_1703;
wire n_6761;
wire n_8972;
wire n_11725;
wire n_13635;
wire n_10801;
wire n_9206;
wire n_3384;
wire n_18488;
wire n_15698;
wire n_1950;
wire n_6811;
wire n_16865;
wire n_18642;
wire n_11622;
wire n_4838;
wire n_12336;
wire n_18345;
wire n_19754;
wire n_12543;
wire n_16129;
wire n_347;
wire n_9705;
wire n_16585;
wire n_17490;
wire n_2965;
wire n_9624;
wire n_3861;
wire n_1977;
wire n_10389;
wire n_3891;
wire n_15688;
wire n_1655;
wire n_13677;
wire n_1886;
wire n_13757;
wire n_14036;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_8982;
wire n_17899;
wire n_13910;
wire n_4673;
wire n_7086;
wire n_3415;
wire n_2947;
wire n_9532;
wire n_18195;
wire n_6601;
wire n_16247;
wire n_13196;
wire n_17482;
wire n_5088;
wire n_19261;
wire n_8034;
wire n_484;
wire n_15824;
wire n_5856;
wire n_9836;
wire n_2497;
wire n_11525;
wire n_11999;
wire n_10837;
wire n_3545;
wire n_18921;
wire n_10554;
wire n_3993;
wire n_8994;
wire n_17827;
wire n_8413;
wire n_4685;
wire n_10149;
wire n_19473;
wire n_19393;
wire n_2663;
wire n_5825;
wire n_2938;
wire n_3780;
wire n_15791;
wire n_12190;
wire n_15484;
wire n_15152;
wire n_11847;
wire n_11976;
wire n_12511;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_8765;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_8213;
wire n_1495;
wire n_14472;
wire n_10534;
wire n_11049;
wire n_14974;
wire n_8451;
wire n_19410;
wire n_1128;
wire n_12743;
wire n_16523;
wire n_8731;
wire n_8385;
wire n_4999;
wire n_15587;
wire n_4922;
wire n_7370;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_18324;
wire n_19383;
wire n_17917;
wire n_7026;
wire n_7053;
wire n_14618;
wire n_9226;
wire n_1765;
wire n_2707;
wire n_18810;
wire n_10608;
wire n_16355;
wire n_7173;
wire n_7042;
wire n_17314;
wire n_718;
wire n_17915;
wire n_5331;
wire n_19225;
wire n_19011;
wire n_16774;
wire n_16436;
wire n_2089;
wire n_10638;
wire n_17923;
wire n_9112;
wire n_18582;
wire n_18970;
wire n_4216;
wire n_19284;
wire n_5797;
wire n_9235;
wire n_16570;
wire n_19124;
wire n_4240;
wire n_3491;
wire n_13852;
wire n_9333;
wire n_704;
wire n_4162;
wire n_17813;
wire n_14089;
wire n_15758;
wire n_1999;
wire n_2731;
wire n_622;
wire n_147;
wire n_3353;
wire n_11804;
wire n_14234;
wire n_3018;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_12809;
wire n_18770;
wire n_4785;
wire n_2002;
wire n_2138;
wire n_2414;
wire n_1771;
wire n_11052;
wire n_3148;
wire n_17350;
wire n_18598;
wire n_6671;
wire n_13470;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_19151;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_13068;
wire n_19158;
wire n_3775;
wire n_18795;
wire n_1176;
wire n_7792;
wire n_15985;
wire n_8161;
wire n_18798;
wire n_5763;
wire n_10014;
wire n_15723;
wire n_16840;
wire n_6029;
wire n_18698;
wire n_10677;
wire n_18269;
wire n_5751;
wire n_15852;
wire n_18857;
wire n_19216;
wire n_12321;
wire n_5924;
wire n_11247;
wire n_290;
wire n_18581;
wire n_8384;
wire n_6445;
wire n_18079;
wire n_13106;
wire n_14294;
wire n_17609;
wire n_6701;
wire n_14862;
wire n_7380;
wire n_8736;
wire n_11514;
wire n_4497;
wire n_1568;
wire n_12470;
wire n_18604;
wire n_12994;
wire n_10215;
wire n_18768;
wire n_14059;
wire n_4871;
wire n_10834;
wire n_17632;
wire n_17611;
wire n_1665;
wire n_19341;
wire n_154;
wire n_12064;
wire n_2127;
wire n_12696;
wire n_18024;
wire n_15735;
wire n_11133;
wire n_5449;
wire n_17143;
wire n_18341;
wire n_10871;
wire n_16405;
wire n_5926;
wire n_2354;
wire n_5398;
wire n_4573;
wire n_14624;
wire n_16600;
wire n_15036;
wire n_17695;
wire n_18193;
wire n_19489;
wire n_11571;
wire n_14120;
wire n_13147;
wire n_8844;
wire n_7641;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_14407;
wire n_14260;
wire n_16845;
wire n_18924;
wire n_17307;
wire n_7169;
wire n_10407;
wire n_19330;
wire n_14175;
wire n_11941;
wire n_4368;
wire n_15780;
wire n_18085;
wire n_1942;
wire n_3196;
wire n_15189;
wire n_8110;
wire n_5319;
wire n_9008;
wire n_12079;
wire n_15335;
wire n_399;
wire n_1440;
wire n_19147;
wire n_2063;
wire n_15227;
wire n_8805;
wire n_7209;
wire n_6014;
wire n_18908;
wire n_15026;
wire n_13895;
wire n_2475;
wire n_5181;
wire n_6979;
wire n_13222;
wire n_3144;
wire n_1268;
wire n_17284;
wire n_5583;
wire n_15987;
wire n_10462;
wire n_642;
wire n_3481;
wire n_11769;
wire n_8856;
wire n_19362;
wire n_303;
wire n_6142;
wire n_14901;
wire n_7769;
wire n_2374;
wire n_416;
wire n_17034;
wire n_10291;
wire n_4597;
wire n_18575;
wire n_18764;
wire n_3364;
wire n_17502;
wire n_14333;
wire n_7233;
wire n_8732;
wire n_13506;
wire n_7602;
wire n_9296;
wire n_18587;
wire n_7390;
wire n_10669;
wire n_19515;
wire n_8231;
wire n_13717;
wire n_5127;
wire n_2920;
wire n_7598;
wire n_12440;
wire n_19032;
wire n_8908;
wire n_1374;
wire n_2648;
wire n_16085;
wire n_1169;
wire n_6767;
wire n_12782;
wire n_3093;
wire n_10111;
wire n_19186;
wire n_19629;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_17796;
wire n_7045;
wire n_3169;
wire n_8740;
wire n_11727;
wire n_6788;
wire n_12192;
wire n_2204;
wire n_177;
wire n_2087;
wire n_17342;
wire n_14465;
wire n_13412;
wire n_4422;
wire n_11749;
wire n_11300;
wire n_6143;
wire n_13457;
wire n_12551;
wire n_18066;
wire n_12497;
wire n_15043;
wire n_4632;
wire n_3084;
wire n_16602;
wire n_2343;
wire n_5967;
wire n_4963;
wire n_16864;
wire n_16761;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_7679;
wire n_18133;
wire n_7936;
wire n_8966;
wire n_4847;
wire n_10287;
wire n_8538;
wire n_12101;
wire n_11145;
wire n_3586;
wire n_3653;
wire n_16684;
wire n_19594;
wire n_725;
wire n_10349;
wire n_4668;
wire n_5213;
wire n_16340;
wire n_7490;
wire n_7545;
wire n_1273;
wire n_9809;
wire n_7160;
wire n_10750;
wire n_617;
wire n_7295;
wire n_14338;
wire n_7348;
wire n_19071;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_17554;
wire n_16071;
wire n_3991;
wire n_15394;
wire n_3516;
wire n_16875;
wire n_15941;
wire n_610;
wire n_9558;
wire n_11594;
wire n_8715;
wire n_12474;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_16655;
wire n_12346;
wire n_517;
wire n_18167;
wire n_4182;
wire n_667;
wire n_8371;
wire n_13916;
wire n_15195;
wire n_1279;
wire n_11458;
wire n_17056;
wire n_12244;
wire n_18753;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_7681;
wire n_11504;
wire n_16850;
wire n_13981;
wire n_4637;
wire n_11516;
wire n_2412;
wire n_8392;
wire n_14659;
wire n_8095;
wire n_10830;
wire n_16868;
wire n_17644;
wire n_5118;
wire n_7503;
wire n_6854;
wire n_17254;
wire n_2757;
wire n_18733;
wire n_4977;
wire n_2716;
wire n_12953;
wire n_2452;
wire n_15224;
wire n_9215;
wire n_11406;
wire n_3043;
wire n_11047;
wire n_14963;
wire n_8050;
wire n_12817;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_16916;
wire n_13866;
wire n_3177;
wire n_12435;
wire n_10946;
wire n_18106;
wire n_7065;
wire n_9216;
wire n_1262;
wire n_4835;
wire n_11961;
wire n_6122;
wire n_7911;
wire n_17486;
wire n_17504;
wire n_14605;
wire n_7330;
wire n_9202;
wire n_2373;
wire n_13543;
wire n_10351;
wire n_13772;
wire n_4734;
wire n_7493;
wire n_12940;
wire n_10460;
wire n_15487;
wire n_19221;
wire n_10334;
wire n_2244;
wire n_11614;
wire n_4290;
wire n_1684;
wire n_1352;
wire n_5407;
wire n_15242;
wire n_8422;
wire n_12224;
wire n_7088;
wire n_9394;
wire n_2704;
wire n_8878;
wire n_7440;
wire n_17681;
wire n_260;
wire n_17676;
wire n_14797;
wire n_9622;
wire n_14177;
wire n_14093;
wire n_3318;
wire n_14607;
wire n_10191;
wire n_4888;
wire n_17919;
wire n_776;
wire n_6000;
wire n_12679;
wire n_14921;
wire n_11168;
wire n_10911;
wire n_12756;
wire n_5004;
wire n_5294;
wire n_16097;
wire n_9845;
wire n_16147;
wire n_7374;
wire n_14389;
wire n_19514;
wire n_11937;
wire n_17277;
wire n_2229;
wire n_4527;
wire n_6046;
wire n_8251;
wire n_5323;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_14621;
wire n_3184;
wire n_18864;
wire n_3075;
wire n_17875;
wire n_11192;
wire n_4949;
wire n_6852;
wire n_8677;
wire n_9091;
wire n_17206;
wire n_13914;
wire n_14663;
wire n_16921;
wire n_17559;
wire n_2536;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_18143;
wire n_16742;
wire n_18464;
wire n_13494;
wire n_5260;
wire n_9751;
wire n_5809;
wire n_10543;
wire n_7924;
wire n_17225;
wire n_560;
wire n_1321;
wire n_7659;
wire n_569;
wire n_3530;
wire n_16203;
wire n_8875;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_1235;
wire n_12662;
wire n_1292;
wire n_15697;
wire n_17879;
wire n_18140;
wire n_9293;
wire n_12503;
wire n_18510;
wire n_15202;
wire n_18218;
wire n_12871;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_18224;
wire n_16400;
wire n_2246;
wire n_4469;
wire n_431;
wire n_10809;
wire n_16934;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_15250;
wire n_17193;
wire n_6711;
wire n_1941;
wire n_11997;
wire n_8946;
wire n_13090;
wire n_18984;
wire n_13541;
wire n_16958;
wire n_4924;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_17396;
wire n_766;
wire n_1746;
wire n_7275;
wire n_8795;
wire n_7195;
wire n_11199;
wire n_17642;
wire n_11264;
wire n_19791;
wire n_2062;
wire n_4539;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_16229;
wire n_10006;
wire n_11757;
wire n_2070;
wire n_18447;
wire n_12622;
wire n_6353;
wire n_4953;
wire n_12659;
wire n_2348;
wire n_6818;
wire n_391;
wire n_2066;
wire n_7539;
wire n_1476;
wire n_12629;
wire n_12868;
wire n_19263;
wire n_10275;
wire n_3458;
wire n_7775;
wire n_11392;
wire n_3190;
wire n_7930;
wire n_7661;
wire n_5383;
wire n_16498;
wire n_19673;
wire n_14165;
wire n_17309;
wire n_19413;
wire n_13787;
wire n_875;
wire n_1678;
wire n_13674;
wire n_18311;
wire n_13912;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_11278;
wire n_14445;
wire n_3787;
wire n_7548;
wire n_16732;
wire n_4450;
wire n_6156;
wire n_12913;
wire n_7064;
wire n_19285;
wire n_16839;
wire n_16798;
wire n_12154;
wire n_8000;
wire n_14427;
wire n_5645;
wire n_3990;
wire n_18327;
wire n_6917;
wire n_6937;
wire n_1628;
wire n_9963;
wire n_988;
wire n_17211;
wire n_7324;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_17568;
wire n_1536;
wire n_6301;
wire n_18061;
wire n_16815;
wire n_18022;
wire n_1132;
wire n_15570;
wire n_15562;
wire n_17207;
wire n_1327;
wire n_19000;
wire n_7729;
wire n_246;
wire n_19622;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_16987;
wire n_18337;
wire n_2380;
wire n_6699;
wire n_12926;
wire n_14809;
wire n_4579;
wire n_14725;
wire n_16892;
wire n_4811;
wire n_19717;
wire n_6874;
wire n_6259;
wire n_9340;
wire n_16527;
wire n_17963;
wire n_6677;
wire n_12161;
wire n_3432;
wire n_11735;
wire n_4282;
wire n_1196;
wire n_8769;
wire n_6764;
wire n_11189;
wire n_10324;
wire n_8815;
wire n_12044;
wire n_748;
wire n_9303;
wire n_1785;
wire n_3057;
wire n_8261;
wire n_13104;
wire n_19730;
wire n_2287;
wire n_7139;
wire n_5727;
wire n_16819;
wire n_16612;
wire n_761;
wire n_5946;
wire n_3778;
wire n_9722;
wire n_12155;
wire n_15664;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_19376;
wire n_14579;
wire n_17930;
wire n_4569;
wire n_8665;
wire n_15847;
wire n_5097;
wire n_7751;
wire n_2234;
wire n_18763;
wire n_14718;
wire n_4384;
wire n_19253;
wire n_2741;
wire n_3114;
wire n_18298;
wire n_888;
wire n_13116;
wire n_19781;
wire n_2203;
wire n_14589;
wire n_5246;
wire n_236;
wire n_12386;
wire n_14257;
wire n_16492;
wire n_16811;
wire n_3836;
wire n_8835;
wire n_18645;
wire n_10688;
wire n_16771;
wire n_1215;
wire n_12964;
wire n_16404;
wire n_15099;
wire n_779;
wire n_2205;
wire n_7579;
wire n_16874;
wire n_4025;
wire n_11687;
wire n_4121;
wire n_8870;
wire n_7155;
wire n_4313;
wire n_6475;
wire n_7699;
wire n_15951;
wire n_6103;
wire n_5546;
wire n_232;
wire n_6394;
wire n_8781;
wire n_18618;
wire n_14102;
wire n_17196;
wire n_4246;
wire n_12267;
wire n_15803;
wire n_8365;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_13780;
wire n_16699;
wire n_7194;
wire n_4049;
wire n_6752;
wire n_6426;
wire n_984;
wire n_5626;
wire n_8025;
wire n_8502;
wire n_7612;
wire n_16999;
wire n_18843;
wire n_11120;
wire n_6350;
wire n_19702;
wire n_7736;
wire n_16040;
wire n_14259;
wire n_5921;
wire n_3596;
wire n_4537;
wire n_6159;
wire n_13360;
wire n_2429;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_3521;
wire n_802;
wire n_17306;
wire n_6235;
wire n_17996;
wire n_2360;
wire n_12647;
wire n_7662;
wire n_15340;
wire n_16061;
wire n_7773;
wire n_5340;
wire n_3947;
wire n_16776;
wire n_13048;
wire n_13563;
wire n_17905;
wire n_7555;
wire n_1194;
wire n_4506;
wire n_19764;
wire n_2742;
wire n_3695;
wire n_12060;
wire n_3976;
wire n_18254;
wire n_10199;
wire n_8658;
wire n_11910;
wire n_15377;
wire n_15583;
wire n_13347;
wire n_5925;
wire n_2909;
wire n_8866;
wire n_8061;
wire n_5730;
wire n_16623;
wire n_17186;
wire n_13111;
wire n_15563;
wire n_10117;
wire n_12716;
wire n_467;
wire n_16341;
wire n_16679;
wire n_13456;
wire n_10198;
wire n_7157;
wire n_13237;
wire n_15448;
wire n_857;
wire n_7411;
wire n_19716;
wire n_16851;
wire n_2221;
wire n_588;
wire n_7871;
wire n_12051;
wire n_1010;
wire n_6477;
wire n_15298;
wire n_11533;
wire n_8652;
wire n_534;
wire n_7198;
wire n_1578;
wire n_9904;
wire n_17891;
wire n_19182;
wire n_1557;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_10973;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_3433;
wire n_17362;
wire n_4463;
wire n_10267;
wire n_10551;
wire n_18589;
wire n_17029;
wire n_3833;
wire n_2774;
wire n_17924;
wire n_18323;
wire n_13127;
wire n_18004;
wire n_4129;
wire n_11002;
wire n_19637;
wire n_5032;
wire n_14075;
wire n_9032;
wire n_6313;
wire n_18884;
wire n_16184;
wire n_3965;
wire n_7145;
wire n_12325;
wire n_9245;
wire n_5065;
wire n_9357;
wire n_3085;
wire n_19060;
wire n_5826;
wire n_15766;
wire n_18121;
wire n_2991;
wire n_16759;
wire n_14530;
wire n_17724;
wire n_19773;
wire n_7994;
wire n_14206;
wire n_17328;
wire n_4703;
wire n_7349;
wire n_9598;
wire n_14481;
wire n_17993;
wire n_15044;
wire n_12504;
wire n_12602;
wire n_12062;
wire n_15375;
wire n_16100;
wire n_12335;
wire n_12949;
wire n_13611;
wire n_801;
wire n_4452;
wire n_15268;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_5362;
wire n_2157;
wire n_10960;
wire n_6141;
wire n_18540;
wire n_3849;
wire n_10931;
wire n_11574;
wire n_15049;
wire n_15181;
wire n_8168;
wire n_3257;
wire n_14870;
wire n_7190;
wire n_1387;
wire n_12322;
wire n_1151;
wire n_14196;
wire n_2317;
wire n_5524;
wire n_10236;
wire n_11776;
wire n_11205;
wire n_11650;
wire n_5818;
wire n_5963;
wire n_19197;
wire n_12179;
wire n_14439;
wire n_9896;
wire n_11856;
wire n_14825;
wire n_11536;
wire n_5950;
wire n_1192;
wire n_14914;
wire n_1844;
wire n_10283;
wire n_5057;
wire n_3030;
wire n_5838;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_2838;
wire n_5325;
wire n_16696;
wire n_18865;
wire n_2926;
wire n_8411;
wire n_2019;
wire n_5102;
wire n_16733;
wire n_18799;
wire n_13221;
wire n_2074;
wire n_2919;
wire n_11163;
wire n_13657;
wire n_945;
wire n_14099;
wire n_15632;
wire n_16245;
wire n_12095;
wire n_13990;
wire n_11419;
wire n_16302;
wire n_9018;
wire n_13663;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_14939;
wire n_11740;
wire n_17471;
wire n_8444;
wire n_17227;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_12392;
wire n_11979;
wire n_7596;
wire n_6280;
wire n_18090;
wire n_18626;
wire n_2786;
wire n_10759;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_18211;
wire n_8977;
wire n_15797;
wire n_9962;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_3107;
wire n_11537;
wire n_13814;
wire n_18993;
wire n_12707;
wire n_14861;
wire n_15194;
wire n_1421;
wire n_7686;
wire n_1936;
wire n_5337;
wire n_18894;
wire n_15572;
wire n_12424;
wire n_1660;
wire n_3047;
wire n_11699;
wire n_8125;
wire n_14811;
wire n_17608;
wire n_10226;
wire n_6526;
wire n_1088;
wire n_17401;
wire n_7196;
wire n_3347;
wire n_907;
wire n_14864;
wire n_4110;
wire n_17936;
wire n_16643;
wire n_1658;
wire n_12107;
wire n_10161;
wire n_9842;
wire n_9614;
wire n_3999;
wire n_16024;
wire n_10699;
wire n_4751;
wire n_7846;
wire n_5151;
wire n_8598;
wire n_7256;
wire n_281;
wire n_16078;
wire n_7331;
wire n_13509;
wire n_17637;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14791;
wire n_14485;
wire n_10606;
wire n_11164;
wire n_4296;
wire n_12203;
wire n_7147;
wire n_5902;
wire n_512;
wire n_12359;
wire n_19175;
wire n_5063;
wire n_9037;
wire n_1328;
wire n_15983;
wire n_12548;
wire n_15874;
wire n_3900;
wire n_3732;
wire n_14461;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_13958;
wire n_17619;
wire n_3980;
wire n_4366;
wire n_6863;
wire n_10012;
wire n_13754;
wire n_12985;
wire n_4445;
wire n_2692;
wire n_16191;
wire n_14171;
wire n_6768;
wire n_4456;
wire n_15212;
wire n_15977;
wire n_9128;
wire n_9872;
wire n_14380;
wire n_10310;
wire n_15896;
wire n_6151;
wire n_16843;
wire n_7110;
wire n_5476;
wire n_17273;
wire n_13920;
wire n_18119;
wire n_2922;
wire n_10097;
wire n_3882;
wire n_2068;
wire n_8915;
wire n_16509;
wire n_9866;
wire n_9858;
wire n_2072;
wire n_586;
wire n_423;
wire n_4375;
wire n_13977;
wire n_8727;
wire n_18494;
wire n_3935;
wire n_5130;
wire n_16538;
wire n_11662;
wire n_1726;
wire n_16992;
wire n_2878;
wire n_18065;
wire n_3012;
wire n_10266;
wire n_17949;
wire n_4877;
wire n_2641;
wire n_8955;
wire n_7734;
wire n_178;
wire n_17781;
wire n_12384;
wire n_15438;
wire n_11260;
wire n_3298;
wire n_11351;
wire n_4467;
wire n_195;
wire n_780;
wire n_15611;
wire n_14388;
wire n_12249;
wire n_2350;
wire n_14977;
wire n_10628;
wire n_13429;
wire n_4220;
wire n_7905;
wire n_5281;
wire n_11775;
wire n_10769;
wire n_10256;
wire n_1654;
wire n_13999;
wire n_14037;
wire n_11706;
wire n_11800;
wire n_18382;
wire n_1588;
wire n_11642;
wire n_4381;
wire n_11143;
wire n_17103;
wire n_11074;
wire n_6831;
wire n_16352;
wire n_18713;
wire n_18032;
wire n_11934;
wire n_4473;
wire n_6043;
wire n_687;
wire n_7677;
wire n_5457;
wire n_10396;
wire n_13919;
wire n_19357;
wire n_190;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_1709;
wire n_10693;
wire n_2657;
wire n_15872;
wire n_13240;
wire n_949;
wire n_3500;
wire n_12578;
wire n_4589;
wire n_12194;
wire n_2972;
wire n_7519;
wire n_7400;
wire n_15649;
wire n_9724;
wire n_9281;
wire n_10101;
wire n_15863;
wire n_6581;
wire n_19690;
wire n_2279;
wire n_161;
wire n_7013;
wire n_14150;
wire n_12125;
wire n_7290;
wire n_18830;
wire n_595;
wire n_4921;
wire n_9687;
wire n_18052;
wire n_19108;
wire n_9426;
wire n_2712;
wire n_7889;
wire n_9102;
wire n_11526;
wire n_16115;
wire n_14128;
wire n_11851;
wire n_898;
wire n_18983;
wire n_17323;
wire n_6965;
wire n_9144;
wire n_18191;
wire n_7461;
wire n_15133;
wire n_16885;
wire n_4137;
wire n_9521;
wire n_15288;
wire n_16900;
wire n_13040;
wire n_963;
wire n_7278;
wire n_6509;
wire n_7454;
wire n_11253;
wire n_17102;
wire n_15527;
wire n_12861;
wire n_17443;
wire n_16146;
wire n_16654;
wire n_3400;
wire n_1521;
wire n_12918;
wire n_1366;
wire n_18332;
wire n_5501;
wire n_5342;
wire n_4345;
wire n_18145;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_16991;
wire n_18051;
wire n_19051;
wire n_4664;
wire n_13716;
wire n_7069;
wire n_7904;
wire n_11691;
wire n_14408;
wire n_9410;
wire n_2643;
wire n_5748;
wire n_12865;
wire n_10712;
wire n_4713;
wire n_7168;
wire n_17604;
wire n_18765;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_3435;
wire n_842;
wire n_10972;
wire n_6359;
wire n_1432;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_8229;
wire n_18743;
wire n_14863;
wire n_5811;
wire n_6766;
wire n_1035;
wire n_7629;
wire n_9735;
wire n_18831;
wire n_5397;
wire n_14711;
wire n_9802;
wire n_1448;
wire n_14373;
wire n_8107;
wire n_12992;
wire n_11108;
wire n_11004;
wire n_2445;
wire n_6519;
wire n_15752;
wire n_11686;
wire n_6530;
wire n_4440;
wire n_10566;
wire n_17798;
wire n_19592;
wire n_16568;
wire n_17581;
wire n_18906;
wire n_12104;
wire n_17954;
wire n_6402;
wire n_12469;
wire n_19554;
wire n_15829;
wire n_19568;
wire n_7326;
wire n_17522;
wire n_7067;
wire n_14835;
wire n_15391;
wire n_16226;
wire n_14871;
wire n_8691;
wire n_14907;
wire n_3342;
wire n_6748;
wire n_11719;
wire n_19307;
wire n_16685;
wire n_19498;
wire n_3656;
wire n_16979;
wire n_1424;
wire n_18282;
wire n_15358;
wire n_14636;
wire n_1507;
wire n_2482;
wire n_8026;
wire n_9638;
wire n_16069;
wire n_7528;
wire n_8174;
wire n_13524;
wire n_912;
wire n_11175;
wire n_10040;
wire n_2661;
wire n_8861;
wire n_5359;
wire n_8644;
wire n_931;
wire n_1791;
wire n_12304;
wire n_15156;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_13138;
wire n_18490;
wire n_6205;
wire n_7136;
wire n_6754;
wire n_12692;
wire n_1334;
wire n_7939;
wire n_13602;
wire n_17436;
wire n_16785;
wire n_9612;
wire n_10790;
wire n_14919;
wire n_16653;
wire n_6723;
wire n_9108;
wire n_16692;
wire n_6440;
wire n_7436;
wire n_14101;
wire n_9376;
wire n_8446;
wire n_17654;
wire n_3534;
wire n_12996;
wire n_15171;
wire n_19711;
wire n_13625;
wire n_12643;
wire n_3944;
wire n_6124;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_19265;
wire n_1939;
wire n_8197;
wire n_2209;
wire n_6622;
wire n_11521;
wire n_12827;
wire n_12678;
wire n_15868;
wire n_1053;
wire n_17249;
wire n_7747;
wire n_9779;
wire n_8082;
wire n_8730;
wire n_15533;
wire n_266;
wire n_6528;
wire n_15165;
wire n_13475;
wire n_15079;
wire n_13859;
wire n_18640;
wire n_1745;
wire n_3479;
wire n_12713;
wire n_13144;
wire n_18129;
wire n_488;
wire n_19488;
wire n_10660;
wire n_7430;
wire n_18560;
wire n_9937;
wire n_5679;
wire n_7912;
wire n_5100;
wire n_16749;
wire n_5973;
wire n_8281;
wire n_4807;
wire n_1243;
wire n_301;
wire n_2928;
wire n_5166;
wire n_19437;
wire n_18876;
wire n_19430;
wire n_11428;
wire n_2822;
wire n_17626;
wire n_1281;
wire n_11677;
wire n_7281;
wire n_9717;
wire n_13577;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_18523;
wire n_1419;
wire n_19176;
wire n_5688;
wire n_13769;
wire n_18044;
wire n_4676;
wire n_13672;
wire n_19036;
wire n_17600;
wire n_6763;
wire n_8956;
wire n_7858;
wire n_663;
wire n_4880;
wire n_6542;
wire n_15681;
wire n_2781;
wire n_4126;
wire n_17262;
wire n_1696;
wire n_6556;
wire n_12374;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_8998;
wire n_10538;
wire n_1790;
wire n_4014;
wire n_13342;
wire n_18856;
wire n_9123;
wire n_17374;
wire n_6471;
wire n_5949;
wire n_15545;
wire n_4048;
wire n_14924;
wire n_4444;
wire n_11867;
wire n_12796;
wire n_3919;
wire n_16053;
wire n_19185;
wire n_15708;
wire n_19441;
wire n_11716;
wire n_8979;
wire n_7245;
wire n_18858;
wire n_6675;
wire n_6270;
wire n_18111;
wire n_6808;
wire n_2884;
wire n_16091;
wire n_11886;
wire n_7006;
wire n_16264;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_17231;
wire n_3797;
wire n_10925;
wire n_4770;
wire n_11158;
wire n_9861;
wire n_15878;
wire n_2549;
wire n_4690;
wire n_14390;
wire n_18678;
wire n_8264;
wire n_7381;
wire n_16160;
wire n_12078;
wire n_15647;
wire n_9832;
wire n_6580;
wire n_18790;
wire n_9898;
wire n_5500;
wire n_6412;
wire n_18410;
wire n_183;
wire n_13293;
wire n_3967;
wire n_6437;
wire n_14381;
wire n_2526;
wire n_15709;
wire n_18590;
wire n_8408;
wire n_3277;
wire n_10661;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_11771;
wire n_16870;
wire n_19082;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_13833;
wire n_16518;
wire n_1960;
wire n_2694;
wire n_1686;
wire n_9867;
wire n_6059;
wire n_14441;
wire n_9688;
wire n_5094;
wire n_10967;
wire n_7870;
wire n_3228;
wire n_18377;
wire n_3657;
wire n_1287;
wire n_6117;
wire n_11828;
wire n_12326;
wire n_1586;
wire n_14264;
wire n_19317;
wire n_14115;
wire n_16635;
wire n_3464;
wire n_380;
wire n_8963;
wire n_4380;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_4193;
wire n_3570;
wire n_12309;
wire n_7399;
wire n_3828;
wire n_1539;
wire n_13953;
wire n_7482;
wire n_14847;
wire n_10312;
wire n_4090;
wire n_18308;
wire n_9223;
wire n_17465;
wire n_15930;
wire n_13226;
wire n_5931;
wire n_2371;
wire n_19416;
wire n_17943;
wire n_662;
wire n_16433;
wire n_3262;
wire n_11244;
wire n_4008;
wire n_18577;
wire n_14432;
wire n_1642;
wire n_10209;
wire n_13253;
wire n_4689;
wire n_8183;
wire n_16098;
wire n_4547;
wire n_11245;
wire n_13354;
wire n_6085;
wire n_12422;
wire n_15616;
wire n_17614;
wire n_3329;
wire n_14422;
wire n_9694;
wire n_3826;
wire n_16636;
wire n_9948;
wire n_14630;
wire n_17048;
wire n_3681;
wire n_18966;
wire n_19390;
wire n_19729;
wire n_10887;
wire n_16876;
wire n_5883;
wire n_6554;
wire n_12146;
wire n_5754;
wire n_6560;
wire n_14055;
wire n_1720;
wire n_12136;
wire n_17046;
wire n_16138;
wire n_12399;
wire n_942;
wire n_12342;
wire n_9744;
wire n_7414;
wire n_9548;
wire n_8973;
wire n_6448;
wire n_1964;
wire n_12378;
wire n_19155;
wire n_12533;
wire n_5434;
wire n_7431;
wire n_5934;
wire n_12178;
wire n_18871;
wire n_11346;
wire n_17210;
wire n_2626;
wire n_5880;
wire n_18206;
wire n_14810;
wire n_8249;
wire n_12257;
wire n_3528;
wire n_15770;
wire n_13394;
wire n_13391;
wire n_14680;
wire n_8234;
wire n_16835;
wire n_1066;
wire n_18438;
wire n_16863;
wire n_9280;
wire n_18285;
wire n_13263;
wire n_14877;
wire n_5145;
wire n_15203;
wire n_1229;
wire n_11491;
wire n_14048;
wire n_2427;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_16112;
wire n_15891;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12769;
wire n_4190;
wire n_5149;
wire n_12641;
wire n_10765;
wire n_3375;
wire n_15263;
wire n_11792;
wire n_18776;
wire n_2668;
wire n_8558;
wire n_10489;
wire n_12421;
wire n_2128;
wire n_7274;
wire n_10159;
wire n_14351;
wire n_7466;
wire n_1002;
wire n_13310;
wire n_2508;
wire n_11568;
wire n_2054;
wire n_7429;
wire n_11766;
wire n_11038;
wire n_13798;
wire n_16894;
wire n_18890;
wire n_17294;
wire n_16932;
wire n_15842;
wire n_14822;
wire n_2758;
wire n_8813;
wire n_10356;
wire n_17461;
wire n_18216;
wire n_10173;
wire n_4789;
wire n_19162;
wire n_12311;
wire n_14374;
wire n_2241;
wire n_6555;
wire n_9448;
wire n_14815;
wire n_10739;
wire n_8470;
wire n_1690;
wire n_5341;
wire n_16480;
wire n_4512;
wire n_1378;
wire n_17657;
wire n_14831;
wire n_11170;
wire n_17683;
wire n_11758;
wire n_1542;
wire n_9396;
wire n_19486;
wire n_14450;
wire n_7061;
wire n_12480;
wire n_14192;
wire n_1716;
wire n_278;
wire n_9053;
wire n_15504;
wire n_11893;
wire n_10573;
wire n_3303;
wire n_4324;
wire n_10850;
wire n_384;
wire n_9185;
wire n_19697;
wire n_13376;
wire n_2905;
wire n_8092;
wire n_13864;
wire n_3954;
wire n_15279;
wire n_11456;
wire n_10546;
wire n_5622;
wire n_3160;
wire n_6574;
wire n_6571;
wire n_17484;
wire n_143;
wire n_9151;
wire n_7824;
wire n_17202;
wire n_18080;
wire n_698;
wire n_13236;
wire n_3569;
wire n_14299;
wire n_7094;
wire n_2528;
wire n_16320;
wire n_4639;
wire n_7036;
wire n_13777;
wire n_19359;
wire n_1730;
wire n_814;
wire n_5779;
wire n_2020;
wire n_6260;
wire n_7413;
wire n_16803;
wire n_17229;
wire n_6286;
wire n_8267;
wire n_4023;
wire n_18929;
wire n_721;
wire n_7175;
wire n_6019;
wire n_4344;
wire n_9978;
wire n_11914;
wire n_9670;
wire n_3154;
wire n_9334;
wire n_15131;
wire n_3898;
wire n_12531;
wire n_4391;
wire n_11302;
wire n_946;
wire n_1303;
wire n_19006;
wire n_4095;
wire n_9413;
wire n_12727;
wire n_15509;
wire n_3551;
wire n_3064;
wire n_11707;
wire n_1689;
wire n_7697;
wire n_1944;
wire n_13835;
wire n_16260;
wire n_7547;
wire n_6013;
wire n_13815;
wire n_9557;
wire n_15957;
wire n_16319;
wire n_448;
wire n_3853;
wire n_17259;
wire n_14039;
wire n_6348;
wire n_6744;
wire n_18578;
wire n_8582;
wire n_5068;
wire n_6293;
wire n_234;
wire n_6049;
wire n_1460;
wire n_9762;
wire n_8957;
wire n_18646;
wire n_15793;
wire n_6558;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_18209;
wire n_2444;
wire n_2437;
wire n_9271;
wire n_17747;
wire n_3035;
wire n_13688;
wire n_4166;
wire n_11396;
wire n_15196;
wire n_16176;
wire n_9483;
wire n_19649;
wire n_1058;
wire n_19435;
wire n_19769;
wire n_14754;
wire n_19768;
wire n_15020;
wire n_2934;
wire n_6091;
wire n_14252;
wire n_15830;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_8747;
wire n_9539;
wire n_4817;
wire n_2014;
wire n_9385;
wire n_1584;
wire n_13462;
wire n_5381;
wire n_9785;
wire n_3468;
wire n_8922;
wire n_9027;
wire n_12750;
wire n_4383;
wire n_6995;
wire n_5696;
wire n_455;
wire n_4486;
wire n_19315;
wire n_9233;
wire n_3024;
wire n_16895;
wire n_10282;
wire n_17602;
wire n_4529;
wire n_500;
wire n_15142;
wire n_291;
wire n_10913;
wire n_18803;
wire n_18409;
wire n_17838;
wire n_15991;
wire n_5823;
wire n_13388;
wire n_2800;
wire n_13731;
wire n_10703;
wire n_9666;
wire n_14503;
wire n_12248;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_17754;
wire n_14886;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_14644;
wire n_11715;
wire n_7071;
wire n_15454;
wire n_10642;
wire n_15213;
wire n_756;
wire n_18859;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_18428;
wire n_12181;
wire n_18670;
wire n_14560;
wire n_17257;
wire n_19726;
wire n_3992;
wire n_14829;
wire n_11007;
wire n_15473;
wire n_249;
wire n_15584;
wire n_3125;
wire n_10316;
wire n_9795;
wire n_18386;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_16515;
wire n_5027;
wire n_17914;
wire n_10479;
wire n_13660;
wire n_19280;
wire n_6801;
wire n_1921;
wire n_18099;
wire n_5630;
wire n_12738;
wire n_4057;
wire n_15062;
wire n_1170;
wire n_5379;
wire n_11599;
wire n_308;
wire n_3444;
wire n_6113;
wire n_10070;
wire n_16178;
wire n_1890;
wire n_18841;
wire n_2477;
wire n_17304;
wire n_18393;
wire n_14983;
wire n_2333;
wire n_8439;
wire n_18434;
wire n_9641;
wire n_1089;
wire n_12755;
wire n_18522;
wire n_12059;
wire n_18541;
wire n_18257;
wire n_15845;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_9138;
wire n_18072;
wire n_18048;
wire n_7537;
wire n_10516;
wire n_15924;
wire n_1616;
wire n_8675;
wire n_17906;
wire n_12567;
wire n_9367;
wire n_15130;
wire n_4197;
wire n_4482;
wire n_2547;
wire n_2415;
wire n_11887;
wire n_17852;
wire n_17442;
wire n_10026;
wire n_9729;
wire n_5073;
wire n_827;
wire n_12471;
wire n_12451;
wire n_17243;
wire n_15740;
wire n_9411;
wire n_3660;
wire n_3766;
wire n_12507;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_14564;
wire n_11277;
wire n_4907;
wire n_5077;
wire n_18416;
wire n_17606;
wire n_7410;
wire n_365;
wire n_8777;
wire n_2534;
wire n_4975;
wire n_13581;
wire n_2451;
wire n_12972;
wire n_13789;
wire n_4815;
wire n_14511;
wire n_13286;
wire n_9951;
wire n_396;
wire n_19023;
wire n_9424;
wire n_480;
wire n_4134;
wire n_10507;
wire n_11968;
wire n_19003;
wire n_1238;
wire n_4092;
wire n_10045;
wire n_11335;
wire n_18606;
wire n_13988;
wire n_4755;
wire n_4960;
wire n_1700;
wire n_15272;
wire n_4933;
wire n_17169;
wire n_13609;
wire n_4591;
wire n_5528;
wire n_16886;
wire n_5111;
wire n_13679;
wire n_11785;
wire n_873;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_12855;
wire n_17370;
wire n_15834;
wire n_13276;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_16058;
wire n_2509;
wire n_11801;
wire n_16994;
wire n_16519;
wire n_3757;
wire n_17810;
wire n_1704;
wire n_250;
wire n_4884;
wire n_14830;
wire n_7867;
wire n_14281;
wire n_14594;
wire n_18213;
wire n_6135;
wire n_17303;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_8669;
wire n_7525;
wire n_19219;
wire n_7257;
wire n_9372;
wire n_4692;
wire n_6791;
wire n_616;
wire n_3165;
wire n_11915;
wire n_13704;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_1902;
wire n_1735;
wire n_3890;
wire n_641;
wire n_3750;
wire n_7650;
wire n_17297;
wire n_13043;
wire n_4311;
wire n_4722;
wire n_17260;
wire n_12620;
wire n_12632;
wire n_6309;
wire n_19618;
wire n_11303;
wire n_405;
wire n_213;
wire n_6733;
wire n_19047;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_9902;
wire n_4820;
wire n_9900;
wire n_17367;
wire n_18937;
wire n_15521;
wire n_18415;
wire n_7202;
wire n_12416;
wire n_8265;
wire n_4619;
wire n_5762;
wire n_11609;
wire n_1961;
wire n_18287;
wire n_16464;
wire n_5036;
wire n_4221;
wire n_19597;
wire n_3297;
wire n_12494;
wire n_10327;
wire n_13826;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_10437;
wire n_10021;
wire n_16673;
wire n_9146;
wire n_15753;
wire n_2996;
wire n_8131;
wire n_8941;
wire n_5014;
wire n_17093;
wire n_17685;
wire n_16357;
wire n_12623;
wire n_11444;
wire n_659;
wire n_6269;
wire n_5233;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_3164;
wire n_9565;
wire n_8257;
wire n_13072;
wire n_18120;
wire n_7726;
wire n_5436;
wire n_17026;
wire n_13839;
wire n_594;
wire n_6120;
wire n_6068;
wire n_4141;
wire n_13954;
wire n_8799;
wire n_2850;
wire n_572;
wire n_6641;
wire n_5789;
wire n_2104;
wire n_19215;
wire n_10124;
wire n_19595;
wire n_14689;
wire n_10245;
wire n_14132;
wire n_10905;
wire n_11235;
wire n_19020;
wire n_6399;
wire n_4499;
wire n_5195;
wire n_9563;
wire n_17077;
wire n_17702;
wire n_11166;
wire n_7031;
wire n_9285;
wire n_263;
wire n_18093;
wire n_16595;
wire n_7763;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_15172;
wire n_4458;
wire n_19470;
wire n_19720;
wire n_5103;
wire n_8393;
wire n_16561;
wire n_10784;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_10944;
wire n_10211;
wire n_18554;
wire n_18077;
wire n_12431;
wire n_11855;
wire n_6790;
wire n_3099;
wire n_17628;
wire n_13799;
wire n_16084;
wire n_13854;
wire n_18250;
wire n_15380;
wire n_2457;
wire n_6686;
wire n_15956;
wire n_4119;
wire n_18835;
wire n_11787;
wire n_5958;
wire n_16059;
wire n_8103;
wire n_2971;
wire n_715;
wire n_4526;
wire n_14752;
wire n_5792;
wire n_6183;
wire n_11544;
wire n_15447;
wire n_10730;
wire n_2028;
wire n_1069;
wire n_10564;
wire n_8682;
wire n_7655;
wire n_18276;
wire n_4485;
wire n_1504;
wire n_11509;
wire n_19191;
wire n_11960;
wire n_1801;
wire n_3917;
wire n_7878;
wire n_9514;
wire n_6210;
wire n_6500;
wire n_12465;
wire n_2206;
wire n_13532;
wire n_11029;
wire n_13118;
wire n_17390;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_19415;
wire n_6785;
wire n_10454;
wire n_15401;
wire n_13339;
wire n_4940;
wire n_8039;
wire n_5757;
wire n_19323;
wire n_8916;
wire n_10087;
wire n_3510;
wire n_10146;
wire n_12959;
wire n_9946;
wire n_9885;
wire n_6849;
wire n_8162;
wire n_18263;
wire n_7457;
wire n_8744;
wire n_5488;
wire n_10701;
wire n_3827;
wire n_891;
wire n_2067;
wire n_7752;
wire n_15775;
wire n_4245;
wire n_17346;
wire n_8286;
wire n_9015;
wire n_6452;
wire n_16408;
wire n_1008;
wire n_6611;
wire n_4560;
wire n_18828;
wire n_4899;
wire n_18297;
wire n_5471;
wire n_11433;
wire n_10592;
wire n_5164;
wire n_18130;
wire n_7207;
wire n_8218;
wire n_17978;
wire n_1767;
wire n_8537;
wire n_10126;
wire n_14421;
wire n_15890;
wire n_4663;
wire n_2893;
wire n_13653;
wire n_5484;
wire n_12566;
wire n_6227;
wire n_13680;
wire n_3421;
wire n_16077;
wire n_9066;
wire n_10302;
wire n_12546;
wire n_13058;
wire n_18342;
wire n_12036;
wire n_17650;
wire n_8782;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_12911;
wire n_15715;
wire n_9857;
wire n_12781;
wire n_10057;
wire n_10882;
wire n_894;
wire n_9338;
wire n_353;
wire n_8144;
wire n_10435;
wire n_9542;
wire n_10921;
wire n_7171;
wire n_12061;
wire n_3922;
wire n_14585;
wire n_11085;
wire n_16541;
wire n_7068;
wire n_13649;
wire n_10609;
wire n_14804;
wire n_2554;
wire n_9783;
wire n_13806;
wire n_19542;
wire n_4934;
wire n_9404;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_18351;
wire n_16198;
wire n_14466;
wire n_7777;
wire n_12138;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_7652;
wire n_10220;
wire n_3150;
wire n_11347;
wire n_17635;
wire n_4479;
wire n_2608;
wire n_10550;
wire n_14673;
wire n_12365;
wire n_1959;
wire n_3133;
wire n_13738;
wire n_14972;
wire n_765;
wire n_1492;
wire n_16996;
wire n_9306;
wire n_14138;
wire n_1340;
wire n_10232;
wire n_10461;
wire n_14586;
wire n_7966;
wire n_8591;
wire n_8811;
wire n_19188;
wire n_1277;
wire n_14031;
wire n_5242;
wire n_10326;
wire n_8417;
wire n_2675;
wire n_5631;
wire n_6008;
wire n_3887;
wire n_12487;
wire n_7997;
wire n_6420;
wire n_4587;
wire n_1577;
wire n_12288;
wire n_17300;
wire n_1117;
wire n_12130;
wire n_13120;
wire n_3223;
wire n_16299;
wire n_12271;
wire n_12704;
wire n_7680;
wire n_15190;
wire n_16909;
wire n_12958;
wire n_8172;
wire n_19559;
wire n_9502;
wire n_6447;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_14761;
wire n_6751;
wire n_2718;
wire n_15243;
wire n_1384;
wire n_11087;
wire n_11477;
wire n_3325;
wire n_2238;
wire n_8375;
wire n_8612;
wire n_4624;
wire n_8345;
wire n_13725;
wire n_3600;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_6741;
wire n_5015;
wire n_1178;
wire n_2338;
wire n_19414;
wire n_17551;
wire n_19417;
wire n_9164;
wire n_7183;
wire n_13197;
wire n_10878;
wire n_18408;
wire n_7140;
wire n_14860;
wire n_10450;
wire n_623;
wire n_19609;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_10529;
wire n_8515;
wire n_1502;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_12254;
wire n_9392;
wire n_1250;
wire n_14531;
wire n_3615;
wire n_11538;
wire n_3087;
wire n_2121;
wire n_9698;
wire n_13435;
wire n_15408;
wire n_15173;
wire n_4015;
wire n_477;
wire n_9644;
wire n_11353;
wire n_18745;
wire n_2213;
wire n_2389;
wire n_9499;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_14771;
wire n_1564;
wire n_5296;
wire n_3718;
wire n_7750;
wire n_11597;
wire n_537;
wire n_15902;
wire n_6277;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_546;
wire n_10920;
wire n_14398;
wire n_3582;
wire n_11126;
wire n_4223;
wire n_5674;
wire n_18453;
wire n_5282;
wire n_9409;
wire n_18629;
wire n_1060;
wire n_1951;
wire n_17814;
wire n_12555;
wire n_11646;
wire n_1223;
wire n_5121;
wire n_9768;
wire n_6070;
wire n_1286;
wire n_12980;
wire n_9881;
wire n_5013;
wire n_6807;
wire n_7251;
wire n_4489;
wire n_7254;
wire n_18178;
wire n_12973;
wire n_3163;
wire n_17313;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_12234;
wire n_10776;
wire n_7882;
wire n_16348;
wire n_16514;
wire n_17704;
wire n_10848;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_11482;
wire n_1625;
wire n_5006;
wire n_7816;
wire n_2226;
wire n_2801;
wire n_10164;
wire n_15809;
wire n_1901;
wire n_3869;
wire n_15579;
wire n_18549;
wire n_18084;
wire n_15585;
wire n_3753;
wire n_12033;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_14376;
wire n_3260;
wire n_9595;
wire n_18978;
wire n_15555;
wire n_13923;
wire n_13051;
wire n_11524;
wire n_17220;
wire n_9265;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_2159;
wire n_2315;
wire n_11228;
wire n_5273;
wire n_7898;
wire n_18286;
wire n_9789;
wire n_5936;
wire n_7646;
wire n_17537;
wire n_3220;
wire n_14627;
wire n_13699;
wire n_6069;
wire n_171;
wire n_169;
wire n_7665;
wire n_9354;
wire n_10501;
wire n_14026;
wire n_2379;
wire n_17782;
wire n_19687;
wire n_9436;
wire n_18157;
wire n_8489;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_12730;
wire n_6887;
wire n_18926;
wire n_16123;
wire n_13152;
wire n_17221;
wire n_4374;
wire n_6637;
wire n_9238;
wire n_358;
wire n_6633;
wire n_2420;
wire n_11031;
wire n_3722;
wire n_186;
wire n_4400;
wire n_17365;
wire n_9839;
wire n_18479;
wire n_15704;
wire n_7900;
wire n_6569;
wire n_10807;
wire n_12478;
wire n_2538;
wire n_724;
wire n_3250;
wire n_17265;
wire n_13545;
wire n_557;
wire n_13760;
wire n_1871;
wire n_13883;
wire n_10511;
wire n_7576;
wire n_19499;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_2102;
wire n_10873;
wire n_14484;
wire n_7676;
wire n_18956;
wire n_9017;
wire n_4304;
wire n_15726;
wire n_14307;
wire n_2544;
wire n_8865;
wire n_15302;
wire n_10337;
wire n_7779;
wire n_8999;
wire n_1206;
wire n_11626;
wire n_12148;
wire n_16872;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_16312;
wire n_16204;
wire n_8820;
wire n_16793;
wire n_16443;
wire n_6090;
wire n_18456;
wire n_5515;
wire n_3131;
wire n_18281;
wire n_12132;
wire n_1298;
wire n_10593;
wire n_5862;
wire n_16801;
wire n_2088;
wire n_12182;
wire n_12043;
wire n_10636;
wire n_16478;
wire n_18489;
wire n_5697;
wire n_2401;
wire n_18723;
wire n_8992;
wire n_8880;
wire n_8690;
wire n_2900;
wire n_6234;
wire n_3994;
wire n_1497;
wire n_7818;
wire n_11721;
wire n_13573;
wire n_19019;
wire n_6608;
wire n_9109;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_7896;
wire n_12482;
wire n_18839;
wire n_15208;
wire n_6860;
wire n_12137;
wire n_12306;
wire n_11328;
wire n_2988;
wire n_1350;
wire n_11200;
wire n_14442;
wire n_15210;
wire n_4109;
wire n_16536;
wire n_13418;
wire n_5175;
wire n_7996;
wire n_986;
wire n_10533;
wire n_460;
wire n_5987;
wire n_16681;
wire n_10176;
wire n_19707;
wire n_7517;
wire n_8080;
wire n_450;
wire n_4150;
wire n_12345;
wire n_13551;
wire n_19135;
wire n_19178;
wire n_16060;
wire n_8772;
wire n_8786;
wire n_15597;
wire n_4643;
wire n_12694;
wire n_8083;
wire n_10155;
wire n_1332;
wire n_9805;
wire n_19799;
wire n_13593;
wire n_8157;
wire n_2346;
wire n_19660;
wire n_936;
wire n_3821;
wire n_13902;
wire n_19792;
wire n_3676;
wire n_4896;
wire n_3675;
wire n_9110;
wire n_18358;
wire n_5904;
wire n_599;
wire n_14468;
wire n_6062;
wire n_12550;
wire n_13861;
wire n_13350;
wire n_10051;
wire n_4209;
wire n_10414;
wire n_8344;
wire n_17597;
wire n_1341;
wire n_8120;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_18882;
wire n_11496;
wire n_4128;
wire n_12225;
wire n_4271;
wire n_2258;
wire n_8621;
wire n_12884;
wire n_325;
wire n_5845;
wire n_19171;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_4716;
wire n_12207;
wire n_9975;
wire n_1782;
wire n_5600;
wire n_12011;
wire n_707;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_6843;
wire n_4715;
wire n_10626;
wire n_6901;
wire n_19014;
wire n_13273;
wire n_4694;
wire n_18855;
wire n_8101;
wire n_19751;
wire n_5448;
wire n_6489;
wire n_7402;
wire n_737;
wire n_3517;
wire n_3893;
wire n_19552;
wire n_11273;
wire n_138;
wire n_19089;
wire n_16954;
wire n_12472;
wire n_19526;
wire n_14035;
wire n_13218;
wire n_9081;
wire n_333;
wire n_4084;
wire n_11762;
wire n_9236;
wire n_6844;
wire n_459;
wire n_4850;
wire n_10156;
wire n_9607;
wire n_2840;
wire n_6779;
wire n_10774;
wire n_12332;
wire n_7216;
wire n_3855;
wire n_15990;
wire n_15364;
wire n_3091;
wire n_6543;
wire n_19585;
wire n_6178;
wire n_9621;
wire n_3398;
wire n_5685;
wire n_18075;
wire n_2793;
wire n_4235;
wire n_16117;
wire n_10398;
wire n_17947;
wire n_16459;
wire n_774;
wire n_17987;
wire n_18165;
wire n_15661;
wire n_17932;
wire n_7706;
wire n_1860;
wire n_5016;
wire n_479;
wire n_6458;
wire n_7642;
wire n_1777;
wire n_12506;
wire n_18356;
wire n_3308;
wire n_12718;
wire n_1600;
wire n_2253;
wire n_12638;
wire n_14116;
wire n_4799;
wire n_2261;
wire n_18710;
wire n_2516;
wire n_16453;
wire n_16645;
wire n_1177;
wire n_10470;
wire n_15034;
wire n_19808;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_12747;
wire n_10625;
wire n_12561;
wire n_18420;
wire n_5514;
wire n_8388;
wire n_18469;
wire n_14730;
wire n_18732;
wire n_9589;
wire n_4543;
wire n_10445;
wire n_15110;
wire n_8988;
wire n_15025;
wire n_19329;
wire n_18161;
wire n_12900;
wire n_18761;
wire n_8569;
wire n_14598;
wire n_3255;
wire n_1401;
wire n_10679;
wire n_1516;
wire n_11323;
wire n_10799;
wire n_2029;
wire n_5890;
wire n_17228;
wire n_1394;
wire n_10585;
wire n_18519;
wire n_13696;
wire n_12948;
wire n_13322;
wire n_7931;
wire n_9092;
wire n_10034;
wire n_935;
wire n_9451;
wire n_11148;
wire n_18729;
wire n_13934;
wire n_6899;
wire n_7373;
wire n_7895;
wire n_676;
wire n_15331;
wire n_17109;
wire n_832;
wire n_13254;
wire n_3049;
wire n_15191;
wire n_17617;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_18783;
wire n_15676;
wire n_17044;
wire n_9011;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_14440;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_372;
wire n_314;
wire n_13875;
wire n_17319;
wire n_17774;
wire n_338;
wire n_19255;
wire n_14076;
wire n_506;
wire n_11220;
wire n_17709;
wire n_9012;
wire n_2396;
wire n_18150;
wire n_2450;
wire n_14638;
wire n_2284;
wire n_19803;
wire n_7238;
wire n_2769;
wire n_14936;
wire n_16469;
wire n_8047;
wire n_11596;
wire n_6273;
wire n_7572;
wire n_5663;
wire n_525;
wire n_11955;
wire n_1677;
wire n_18818;
wire n_16156;
wire n_11654;
wire n_18361;
wire n_12982;
wire n_4160;
wire n_4231;
wire n_11619;
wire n_10649;
wire n_2779;
wire n_5203;
wire n_19638;
wire n_6311;
wire n_7590;
wire n_5162;
wire n_1464;
wire n_5285;
wire n_2721;
wire n_12275;
wire n_13742;
wire n_270;
wire n_15177;
wire n_12376;
wire n_563;
wire n_13114;
wire n_8583;
wire n_4521;
wire n_10447;
wire n_15063;
wire n_7176;
wire n_9353;
wire n_13054;
wire n_8948;
wire n_5715;
wire n_8295;
wire n_498;
wire n_5395;
wire n_10522;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_1693;
wire n_16618;
wire n_10278;
wire n_15384;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_2915;
wire n_15686;
wire n_9263;
wire n_11082;
wire n_1989;
wire n_15950;
wire n_2802;
wire n_19724;
wire n_6181;
wire n_7447;
wire n_17998;
wire n_19156;
wire n_18928;
wire n_12721;
wire n_18301;
wire n_5672;
wire n_16008;
wire n_11730;
wire n_3098;
wire n_6924;
wire n_9804;
wire n_1851;
wire n_9304;
wire n_5799;
wire n_8380;
wire n_12039;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_10377;
wire n_9926;
wire n_570;
wire n_15161;
wire n_620;
wire n_2523;
wire n_10858;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_16303;
wire n_9843;
wire n_3130;
wire n_16559;
wire n_1710;
wire n_13320;
wire n_1301;
wire n_6683;
wire n_10683;
wire n_2282;
wire n_9921;
wire n_19606;
wire n_6229;
wire n_1609;
wire n_13488;
wire n_15907;
wire n_7286;
wire n_13668;
wire n_13016;
wire n_6177;
wire n_16961;
wire n_14708;
wire n_2867;
wire n_2726;
wire n_17293;
wire n_12048;
wire n_5982;
wire n_10930;
wire n_17972;
wire n_8749;
wire n_18264;
wire n_2662;
wire n_12057;
wire n_6696;
wire n_17590;
wire n_9527;
wire n_16450;
wire n_19651;
wire n_2795;
wire n_18352;
wire n_14875;
wire n_3472;
wire n_15056;
wire n_15860;
wire n_19460;
wire n_17288;
wire n_5376;
wire n_16197;
wire n_14003;
wire n_5106;
wire n_9511;
wire n_6730;
wire n_17822;
wire n_13670;
wire n_11254;
wire n_15023;
wire n_11617;
wire n_18184;
wire n_5561;
wire n_404;
wire n_158;
wire n_18436;
wire n_6170;
wire n_9459;
wire n_14185;
wire n_6094;
wire n_9098;
wire n_14953;
wire n_15604;
wire n_4826;
wire n_16000;
wire n_3903;
wire n_12360;
wire n_9268;
wire n_17116;
wire n_15431;
wire n_3854;
wire n_3235;
wire n_8673;
wire n_18702;
wire n_19174;
wire n_5378;
wire n_10456;
wire n_3673;
wire n_13186;
wire n_18824;
wire n_5916;
wire n_15655;
wire n_11907;
wire n_3094;
wire n_10627;
wire n_10475;
wire n_965;
wire n_1428;
wire n_15430;
wire n_1576;
wire n_2077;
wire n_8581;
wire n_15732;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_4951;
wire n_17772;
wire n_540;
wire n_14170;
wire n_3070;
wire n_13496;
wire n_8058;
wire n_9308;
wire n_3504;
wire n_11838;
wire n_10508;
wire n_18008;
wire n_10811;
wire n_18696;
wire n_8333;
wire n_17152;
wire n_7619;
wire n_6985;
wire n_18551;
wire n_7170;
wire n_13853;
wire n_8823;
wire n_11457;
wire n_12751;
wire n_15284;
wire n_3054;
wire n_5399;
wire n_4620;
wire n_5421;
wire n_4127;
wire n_17901;
wire n_15443;
wire n_5206;
wire n_18228;
wire n_17833;
wire n_18471;
wire n_4517;
wire n_16852;
wire n_18817;
wire n_6916;
wire n_15524;
wire n_2260;
wire n_10725;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_18354;
wire n_8290;
wire n_7536;
wire n_1743;
wire n_18152;
wire n_6230;
wire n_16108;
wire n_11107;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_12757;
wire n_14379;
wire n_8840;
wire n_16284;
wire n_16001;
wire n_18873;
wire n_13189;
wire n_5881;
wire n_18915;
wire n_2382;
wire n_3754;
wire n_19492;
wire n_12328;
wire n_415;
wire n_9083;
wire n_17271;
wire n_383;
wire n_2974;
wire n_4213;
wire n_200;
wire n_6483;
wire n_10994;
wire n_14004;
wire n_17023;
wire n_5863;
wire n_2645;
wire n_16221;
wire n_3904;
wire n_8036;
wire n_11485;
wire n_1444;
wire n_7300;
wire n_6975;
wire n_14666;
wire n_1263;
wire n_13605;
wire n_17387;
wire n_11048;
wire n_4733;
wire n_14237;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_11240;
wire n_13841;
wire n_3080;
wire n_11634;
wire n_12580;
wire n_10013;
wire n_17166;
wire n_2865;
wire n_16119;
wire n_6076;
wire n_8933;
wire n_19344;
wire n_15876;
wire n_18819;
wire n_15231;
wire n_11287;
wire n_943;
wire n_9774;
wire n_4879;
wire n_6390;
wire n_13409;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_9720;
wire n_15727;
wire n_10169;
wire n_12690;
wire n_7563;
wire n_12475;
wire n_1345;
wire n_4556;
wire n_11765;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_19510;
wire n_4117;
wire n_14414;
wire n_15565;
wire n_5995;
wire n_17823;
wire n_2378;
wire n_5905;
wire n_9149;
wire n_2655;
wire n_7035;
wire n_6193;
wire n_1467;
wire n_4250;
wire n_16858;
wire n_16980;
wire n_224;
wire n_3963;
wire n_9345;
wire n_11550;
wire n_17315;
wire n_7527;
wire n_13061;
wire n_9682;
wire n_2214;
wire n_17719;
wire n_6582;
wire n_18432;
wire n_12545;
wire n_18320;
wire n_1230;
wire n_3850;
wire n_18078;
wire n_9924;
wire n_14744;
wire n_15091;
wire n_5525;
wire n_17527;
wire n_163;
wire n_1644;
wire n_12753;
wire n_2277;
wire n_7090;
wire n_9254;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_11641;
wire n_7415;
wire n_11211;
wire n_13375;
wire n_13691;
wire n_824;
wire n_6745;
wire n_6972;
wire n_18526;
wire n_16913;
wire n_16663;
wire n_11857;
wire n_395;
wire n_6240;
wire n_13482;
wire n_18069;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_9469;
wire n_15869;
wire n_2961;
wire n_15598;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_483;
wire n_16604;
wire n_2546;
wire n_13873;
wire n_15805;
wire n_476;
wire n_1957;
wire n_17836;
wire n_4732;
wire n_18769;
wire n_11201;
wire n_10531;
wire n_14964;
wire n_8918;
wire n_12878;
wire n_19273;
wire n_8932;
wire n_17756;
wire n_4581;
wire n_16603;
wire n_9249;
wire n_2143;
wire n_8180;
wire n_15580;
wire n_9444;
wire n_10772;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_15984;
wire n_6770;
wire n_17730;
wire n_15151;
wire n_16626;
wire n_5639;
wire n_487;
wire n_8943;
wire n_14767;
wire n_18463;
wire n_4503;
wire n_14773;
wire n_10127;
wire n_13654;
wire n_5361;
wire n_11814;
wire n_12255;
wire n_4199;
wire n_1912;
wire n_9723;
wire n_19446;
wire n_19669;
wire n_1982;
wire n_3872;
wire n_1312;
wire n_19577;
wire n_5330;
wire n_7199;
wire n_10039;
wire n_11358;
wire n_10854;
wire n_13366;
wire n_247;
wire n_5892;
wire n_7940;
wire n_16467;
wire n_6782;
wire n_18746;
wire n_2008;
wire n_2192;
wire n_328;
wire n_17669;
wire n_1386;
wire n_6503;
wire n_19423;
wire n_12017;
wire n_17357;
wire n_15381;
wire n_18477;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_16103;
wire n_19041;
wire n_16460;
wire n_690;
wire n_8271;
wire n_4800;
wire n_1157;
wire n_12728;
wire n_1752;
wire n_16651;
wire n_4958;
wire n_6783;
wire n_12259;
wire n_8699;
wire n_16305;
wire n_19409;
wire n_2963;
wire n_15861;
wire n_3873;
wire n_8225;
wire n_9536;
wire n_14250;
wire n_16818;
wire n_16573;
wire n_18671;
wire n_16562;
wire n_6296;
wire n_7708;
wire n_11671;
wire n_10328;
wire n_5968;
wire n_2644;
wire n_3326;
wire n_6497;
wire n_15705;
wire n_2411;
wire n_16816;
wire n_7333;
wire n_15376;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_18035;
wire n_7371;
wire n_17547;
wire n_8152;
wire n_15050;
wire n_10826;
wire n_7463;
wire n_8525;
wire n_17767;
wire n_18680;
wire n_283;
wire n_12160;
wire n_590;
wire n_9620;
wire n_1990;
wire n_3805;
wire n_5205;
wire n_17145;
wire n_11119;
wire n_7954;
wire n_1465;
wire n_2622;
wire n_7951;
wire n_8096;
wire n_13901;
wire n_7231;
wire n_5080;
wire n_3128;
wire n_15252;
wire n_18043;
wire n_16238;
wire n_5372;
wire n_14050;
wire n_15763;
wire n_17983;
wire n_2691;
wire n_15317;
wire n_7772;
wire n_2690;
wire n_14197;
wire n_18159;
wire n_19364;
wire n_8996;
wire n_12070;
wire n_9714;
wire n_3078;
wire n_14898;
wire n_15672;
wire n_3793;
wire n_15920;
wire n_11928;
wire n_5071;
wire n_14395;
wire n_5801;
wire n_13528;
wire n_6047;
wire n_8292;
wire n_8601;
wire n_9377;
wire n_11932;
wire n_6970;
wire n_19328;
wire n_1308;
wire n_13027;
wire n_12607;
wire n_7272;
wire n_15782;
wire n_19553;
wire n_12075;
wire n_4540;
wire n_13489;
wire n_2097;
wire n_18887;
wire n_3499;
wire n_19693;
wire n_19797;
wire n_13877;
wire n_1005;
wire n_6209;
wire n_11922;
wire n_14020;
wire n_1469;
wire n_12358;
wire n_7408;
wire n_2650;
wire n_10488;
wire n_8969;
wire n_14187;
wire n_11577;
wire n_17840;
wire n_16914;
wire n_18513;
wire n_153;
wire n_3348;
wire n_19165;
wire n_17907;
wire n_11475;
wire n_9048;
wire n_5228;
wire n_10274;
wire n_1723;
wire n_189;
wire n_6694;
wire n_15318;
wire n_9168;
wire n_14220;
wire n_13837;
wire n_2335;
wire n_18570;
wire n_529;
wire n_5507;
wire n_5569;
wire n_15559;
wire n_16871;
wire n_14221;
wire n_13964;
wire n_10832;
wire n_3173;
wire n_18829;
wire n_6856;
wire n_1049;
wire n_6466;
wire n_16039;
wire n_7864;
wire n_18295;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_1717;
wire n_2449;
wire n_3880;
wire n_13601;
wire n_17457;
wire n_17115;
wire n_19281;
wire n_18155;
wire n_4545;
wire n_272;
wire n_6820;
wire n_2896;
wire n_2639;
wire n_17083;
wire n_458;
wire n_5490;
wire n_19007;
wire n_4771;
wire n_13392;
wire n_5836;
wire n_17563;
wire n_9169;
wire n_252;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_3561;
wire n_19008;
wire n_18401;
wire n_6469;
wire n_6700;
wire n_3032;
wire n_6223;
wire n_11398;
wire n_8798;
wire n_9600;
wire n_2877;
wire n_11274;
wire n_8085;
wire n_1021;
wire n_8123;
wire n_811;
wire n_17997;
wire n_12512;
wire n_9927;
wire n_5497;
wire n_16973;
wire n_15657;
wire n_17571;
wire n_3598;
wire n_7127;
wire n_831;
wire n_15513;
wire n_8666;
wire n_2435;
wire n_12284;
wire n_18322;
wire n_1382;
wire n_7801;
wire n_9155;
wire n_1483;
wire n_10416;
wire n_15837;
wire n_1372;
wire n_14370;
wire n_1719;
wire n_7959;
wire n_13430;
wire n_1427;
wire n_2745;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_10583;
wire n_10806;
wire n_2323;
wire n_162;
wire n_5234;
wire n_7546;
wire n_6272;
wire n_14274;
wire n_6588;
wire n_3265;
wire n_3755;
wire n_4042;
wire n_18125;
wire n_15403;
wire n_13081;
wire n_15602;
wire n_12252;
wire n_16743;
wire n_10439;
wire n_12627;
wire n_19378;
wire n_16730;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_2410;
wire n_18868;
wire n_6222;
wire n_15012;
wire n_1783;
wire n_4176;
wire n_14551;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_7521;
wire n_12968;
wire n_10663;
wire n_15517;
wire n_3894;
wire n_13974;
wire n_12277;
wire n_14917;
wire n_3127;
wire n_3623;
wire n_5312;
wire n_16075;
wire n_6625;
wire n_15680;
wire n_2502;
wire n_3646;
wire n_17441;
wire n_14855;
wire n_16757;
wire n_2783;
wire n_8487;
wire n_4034;
wire n_18601;
wire n_1470;
wire n_8141;
wire n_4887;
wire n_14058;
wire n_11020;
wire n_13141;
wire n_16461;
wire n_14065;
wire n_11920;
wire n_19756;
wire n_17299;
wire n_3862;
wire n_14366;
wire n_10481;
wire n_19250;
wire n_6876;
wire n_16022;
wire n_5049;
wire n_19001;
wire n_19627;
wire n_9573;
wire n_5846;
wire n_17235;
wire n_7636;
wire n_9799;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_1855;
wire n_3051;
wire n_15143;
wire n_11198;
wire n_18932;
wire n_18346;
wire n_18238;
wire n_385;
wire n_1439;
wire n_2859;
wire n_1331;
wire n_19794;
wire n_5157;
wire n_3525;
wire n_2100;
wire n_11840;
wire n_13157;
wire n_1134;
wire n_10261;
wire n_4003;
wire n_5708;
wire n_3751;
wire n_4894;
wire n_14084;
wire n_4113;
wire n_5649;
wire n_9827;
wire n_13334;
wire n_10907;
wire n_4983;
wire n_14002;
wire n_419;
wire n_7214;
wire n_3907;
wire n_16205;
wire n_13399;
wire n_1254;
wire n_7075;
wire n_19503;
wire n_14697;
wire n_7124;
wire n_13967;
wire n_3291;
wire n_2304;
wire n_7799;
wire n_5698;
wire n_11092;
wire n_14310;
wire n_5084;
wire n_15792;
wire n_15281;
wire n_15675;
wire n_8917;
wire n_9647;
wire n_15515;
wire n_15106;
wire n_4710;
wire n_12067;
wire n_9214;
wire n_17030;
wire n_19537;
wire n_4101;
wire n_7776;
wire n_19621;
wire n_14309;
wire n_9864;
wire n_16256;
wire n_3236;
wire n_17416;
wire n_16741;
wire n_923;
wire n_11770;
wire n_19201;
wire n_13996;
wire n_17944;
wire n_17679;
wire n_9000;
wire n_18442;
wire n_18505;
wire n_10864;
wire n_18412;
wire n_14704;
wire n_8307;
wire n_9383;
wire n_17692;
wire n_4611;
wire n_15258;
wire n_2337;
wire n_12174;
wire n_16322;
wire n_15220;
wire n_19611;
wire n_6400;
wire n_16304;
wire n_18417;
wire n_13504;
wire n_7543;
wire n_16787;
wire n_13169;
wire n_7877;
wire n_9672;
wire n_15291;
wire n_18375;
wire n_8855;
wire n_8885;
wire n_5486;
wire n_15345;
wire n_137;
wire n_1596;
wire n_5092;
wire n_14721;
wire n_1734;
wire n_3172;
wire n_13265;
wire n_4832;
wire n_2902;
wire n_12153;
wire n_7284;
wire n_7264;
wire n_13666;
wire n_19192;
wire n_6537;
wire n_10702;
wire n_13730;
wire n_3536;
wire n_12405;
wire n_2894;
wire n_3710;
wire n_4195;
wire n_10319;
wire n_9654;
wire n_8802;
wire n_9859;
wire n_5240;
wire n_2225;
wire n_6092;
wire n_6241;
wire n_1692;
wire n_8667;
wire n_18996;
wire n_2006;
wire n_3402;
wire n_8121;
wire n_9645;
wire n_7754;
wire n_15549;
wire n_18777;
wire n_2789;
wire n_12792;
wire n_1828;
wire n_19661;
wire n_9796;
wire n_8320;
wire n_18219;
wire n_18231;
wire n_4862;
wire n_15889;
wire n_2376;
wire n_12438;
wire n_11830;
wire n_8766;
wire n_16665;
wire n_16173;
wire n_9165;
wire n_2700;
wire n_19555;
wire n_1041;
wire n_12539;
wire n_565;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_18461;
wire n_14369;
wire n_1062;
wire n_7240;
wire n_15354;
wire n_10476;
wire n_9966;
wire n_16794;
wire n_1222;
wire n_2635;
wire n_11486;
wire n_15999;
wire n_15280;
wire n_12677;
wire n_4321;
wire n_7237;
wire n_17867;
wire n_16456;
wire n_6877;
wire n_12873;
wire n_16364;
wire n_6949;
wire n_19356;
wire n_17036;
wire n_19698;
wire n_806;
wire n_13401;
wire n_584;
wire n_12276;
wire n_9893;
wire n_14122;
wire n_17565;
wire n_8126;
wire n_15819;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4757;
wire n_15603;
wire n_12352;
wire n_17267;
wire n_2809;
wire n_18528;
wire n_787;
wire n_10099;
wire n_9961;
wire n_16833;
wire n_14895;
wire n_7163;
wire n_1528;
wire n_1146;
wire n_16582;
wire n_18028;
wire n_2021;
wire n_15270;
wire n_17964;
wire n_10181;
wire n_15670;
wire n_4604;
wire n_5724;
wire n_7201;
wire n_3157;
wire n_16825;
wire n_2422;
wire n_10949;
wire n_3457;
wire n_3762;
wire n_18197;
wire n_3411;
wire n_4519;
wire n_5355;
wire n_13969;
wire n_16548;
wire n_5186;
wire n_1498;
wire n_12693;
wire n_6792;
wire n_1210;
wire n_9316;
wire n_5438;
wire n_13259;
wire n_1269;
wire n_19164;
wire n_14954;
wire n_12648;
wire n_655;
wire n_4726;
wire n_6045;
wire n_1872;
wire n_9914;
wire n_8132;
wire n_19541;
wire n_10917;
wire n_16050;
wire n_3761;
wire n_18006;
wire n_7821;
wire n_12407;
wire n_11284;
wire n_14668;
wire n_14776;
wire n_10458;
wire n_2041;
wire n_11656;
wire n_13134;
wire n_10271;
wire n_15415;
wire n_16808;
wire n_18902;
wire n_1098;
wire n_5746;
wire n_6673;
wire n_18207;
wire n_11909;
wire n_12637;
wire n_7887;
wire n_398;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_3726;
wire n_12009;
wire n_2369;
wire n_13612;
wire n_19388;
wire n_10648;
wire n_2587;
wire n_7550;
wire n_17498;
wire n_15077;
wire n_3199;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_15733;
wire n_15864;
wire n_14207;
wire n_1953;
wire n_19080;
wire n_19736;
wire n_13863;
wire n_14305;
wire n_9863;
wire n_15330;
wire n_10500;
wire n_5432;
wire n_15261;
wire n_11929;
wire n_11075;
wire n_7851;
wire n_16605;
wire n_9791;
wire n_19228;
wire n_5453;
wire n_4900;
wire n_11177;
wire n_19761;
wire n_13667;
wire n_18056;
wire n_5842;
wire n_13126;
wire n_7798;
wire n_5253;
wire n_10857;
wire n_18491;
wire n_11310;
wire n_13275;
wire n_11165;
wire n_14411;
wire n_12823;
wire n_2953;
wire n_15412;
wire n_4295;
wire n_5943;
wire n_12193;
wire n_2500;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_15257;
wire n_19701;
wire n_8528;
wire n_8204;
wire n_11733;
wire n_15646;
wire n_1389;
wire n_18214;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_18347;
wire n_14738;
wire n_12242;
wire n_5610;
wire n_3015;
wire n_13796;
wire n_10502;
wire n_15522;
wire n_17577;
wire n_17874;
wire n_6722;
wire n_17892;
wire n_7622;
wire n_11123;
wire n_8512;
wire n_14464;
wire n_387;
wire n_744;
wire n_971;
wire n_8635;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_1205;
wire n_15535;
wire n_16633;
wire n_7831;
wire n_10227;
wire n_10574;
wire n_19271;
wire n_2180;
wire n_16323;
wire n_2858;
wire n_18624;
wire n_6201;
wire n_12218;
wire n_5737;
wire n_3604;
wire n_12343;
wire n_4373;
wire n_8919;
wire n_17014;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_4711;
wire n_11478;
wire n_16067;
wire n_3068;
wire n_15650;
wire n_12236;
wire n_12902;
wire n_16230;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_13038;
wire n_2465;
wire n_12892;
wire n_17768;
wire n_3811;
wire n_11294;
wire n_910;
wire n_15667;
wire n_3486;
wire n_4086;
wire n_10289;
wire n_6565;
wire n_6942;
wire n_11819;
wire n_19389;
wire n_2032;
wire n_4812;
wire n_13420;
wire n_6862;
wire n_5858;
wire n_17200;
wire n_15053;
wire n_13005;
wire n_708;
wire n_14805;
wire n_6037;
wire n_2312;
wire n_11844;
wire n_1266;
wire n_15390;
wire n_6635;
wire n_185;
wire n_13184;
wire n_1276;
wire n_13535;
wire n_14982;
wire n_12247;
wire n_14770;
wire n_11100;
wire n_298;
wire n_1582;
wire n_5588;
wire n_3286;
wire n_19350;
wire n_7167;
wire n_6480;
wire n_15105;
wire n_5075;
wire n_3682;
wire n_18927;
wire n_3771;
wire n_18383;
wire n_12765;
wire n_7865;
wire n_15690;
wire n_9289;
wire n_11315;
wire n_6561;
wire n_12706;
wire n_11153;
wire n_17128;
wire n_859;
wire n_406;
wire n_6875;
wire n_10934;
wire n_1770;
wire n_10197;
wire n_18999;
wire n_3285;
wire n_19584;
wire n_11949;
wire n_8402;
wire n_9690;
wire n_2071;
wire n_11746;
wire n_9371;
wire n_19689;
wire n_16837;
wire n_7267;
wire n_4599;
wire n_12315;
wire n_18668;
wire n_5222;
wire n_7850;
wire n_14100;
wire n_12998;
wire n_7812;
wire n_13143;
wire n_9080;
wire n_14549;
wire n_8133;
wire n_6176;
wire n_14717;
wire n_3881;
wire n_16426;
wire n_14459;
wire n_4508;
wire n_11530;
wire n_13411;
wire n_7056;
wire n_8193;
wire n_12445;
wire n_12856;
wire n_19520;
wire n_7813;
wire n_7514;
wire n_7649;
wire n_18734;
wire n_12525;
wire n_16116;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_15823;
wire n_5832;
wire n_13758;
wire n_1305;
wire n_7688;
wire n_4562;
wire n_16820;
wire n_3383;
wire n_8707;
wire n_12357;
wire n_9208;
wire n_11791;
wire n_19525;
wire n_7611;
wire n_19778;
wire n_17218;
wire n_15216;
wire n_11848;
wire n_3610;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_12180;
wire n_2065;
wire n_15608;
wire n_10935;
wire n_2001;
wire n_7723;
wire n_11621;
wire n_19448;
wire n_225;
wire n_16171;
wire n_3555;
wire n_7450;
wire n_11667;
wire n_17311;
wire n_7362;
wire n_17455;
wire n_12208;
wire n_1131;
wire n_3110;
wire n_14565;
wire n_17248;
wire n_11298;
wire n_15796;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_13314;
wire n_670;
wire n_11741;
wire n_3908;
wire n_15537;
wire n_3467;
wire n_12773;
wire n_9044;
wire n_12381;
wire n_19302;
wire n_18174;
wire n_14883;
wire n_17024;
wire n_6451;
wire n_9813;
wire n_1226;
wire n_3740;
wire n_18482;
wire n_3186;
wire n_640;
wire n_17322;
wire n_9244;
wire n_15304;
wire n_7049;
wire n_15271;
wire n_2632;
wire n_14865;
wire n_8278;
wire n_11644;
wire n_6345;
wire n_15893;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_364;
wire n_5782;
wire n_5041;
wire n_13170;
wire n_1915;
wire n_4275;
wire n_14471;
wire n_11357;
wire n_19387;
wire n_4425;
wire n_9985;
wire n_4449;
wire n_12089;
wire n_7057;
wire n_17888;
wire n_11959;
wire n_19586;
wire n_1612;
wire n_4809;
wire n_12987;
wire n_8529;
wire n_625;
wire n_10254;
wire n_18625;
wire n_14715;
wire n_15970;
wire n_11208;
wire n_15978;
wire n_12452;
wire n_15961;
wire n_8574;
wire n_1038;
wire n_12292;
wire n_4241;
wire n_12818;
wire n_11420;
wire n_12500;
wire n_8044;
wire n_16330;
wire n_9439;
wire n_1380;
wire n_15239;
wire n_2557;
wire n_11630;
wire n_2405;
wire n_19759;
wire n_15444;
wire n_15289;
wire n_13172;
wire n_2336;
wire n_16234;
wire n_2521;
wire n_9120;
wire n_17335;
wire n_17610;
wire n_19522;
wire n_424;
wire n_12168;
wire n_16496;
wire n_8903;
wire n_141;
wire n_1985;
wire n_16057;
wire n_16401;
wire n_4531;
wire n_3282;
wire n_15781;
wire n_14448;
wire n_1532;
wire n_11017;
wire n_7247;
wire n_14622;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_14739;
wire n_16649;
wire n_12613;
wire n_14365;
wire n_9325;
wire n_16448;
wire n_4555;
wire n_17173;
wire n_9384;
wire n_6216;
wire n_7340;
wire n_12695;
wire n_15467;
wire n_4308;
wire n_14219;
wire n_3463;
wire n_11576;
wire n_1954;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_3998;
wire n_12006;
wire n_2495;
wire n_10128;
wire n_371;
wire n_18319;
wire n_12246;
wire n_18220;
wire n_9955;
wire n_19477;
wire n_3829;
wire n_9007;
wire n_10143;
wire n_1471;
wire n_18715;
wire n_3655;
wire n_17884;
wire n_3825;
wire n_2880;
wire n_13085;
wire n_19260;
wire n_7780;
wire n_8452;
wire n_11518;
wire n_5670;
wire n_8557;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_18892;
wire n_11252;
wire n_8012;
wire n_1445;
wire n_1526;
wire n_17055;
wire n_1978;
wire n_6472;
wire n_18067;
wire n_574;
wire n_8114;
wire n_4202;
wire n_16227;
wire n_5879;
wire n_14563;
wire n_4403;
wire n_5238;
wire n_16329;
wire n_11256;
wire n_6166;
wire n_12370;
wire n_9136;
wire n_12860;
wire n_16278;
wire n_473;
wire n_17404;
wire n_559;
wire n_19635;
wire n_7063;
wire n_14768;
wire n_4139;
wire n_13885;
wire n_1986;
wire n_13631;
wire n_18103;
wire n_6081;
wire n_16746;
wire n_15929;
wire n_6724;
wire n_813;
wire n_11336;
wire n_12758;
wire n_17410;
wire n_19248;
wire n_11849;
wire n_3910;
wire n_9204;
wire n_9476;
wire n_12142;
wire n_9689;
wire n_16711;
wire n_10659;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_6946;
wire n_3319;
wire n_12983;
wire n_3748;
wire n_6424;
wire n_11210;
wire n_7599;
wire n_16271;
wire n_15541;
wire n_13980;
wire n_16366;
wire n_982;
wire n_11191;
wire n_10547;
wire n_6778;
wire n_17359;
wire n_13205;
wire n_1697;
wire n_979;
wire n_5544;
wire n_5067;
wire n_15283;
wire n_12396;
wire n_15407;
wire n_7614;
wire n_19381;
wire n_1278;
wire n_7839;
wire n_9837;
wire n_634;
wire n_10896;
wire n_136;
wire n_17761;
wire n_4130;
wire n_10562;
wire n_16042;
wire n_5941;
wire n_2009;
wire n_14417;
wire n_6340;
wire n_3601;
wire n_10355;
wire n_10054;
wire n_1289;
wire n_16893;
wire n_3055;
wire n_6706;
wire n_3966;
wire n_13034;
wire n_1014;
wire n_16828;
wire n_10007;
wire n_882;
wire n_11751;
wire n_17550;
wire n_3746;
wire n_17185;
wire n_14637;
wire n_11495;
wire n_4478;
wire n_1662;
wire n_17015;
wire n_7372;
wire n_19617;
wire n_2818;
wire n_17980;
wire n_674;
wire n_3921;
wire n_17535;
wire n_16822;
wire n_10704;
wire n_11520;
wire n_1927;
wire n_19614;
wire n_12169;
wire n_16788;
wire n_15088;
wire n_17976;
wire n_702;
wire n_4965;
wire n_16383;
wire n_17538;
wire n_11012;
wire n_6111;
wire n_11502;
wire n_15348;
wire n_11631;
wire n_13588;
wire n_13570;
wire n_2193;
wire n_4523;
wire n_6011;
wire n_11842;
wire n_14710;
wire n_3153;
wire n_877;
wire n_13737;
wire n_16590;
wire n_728;
wire n_18188;
wire n_4607;
wire n_16640;
wire n_11389;
wire n_7226;
wire n_9013;
wire n_18373;
wire n_4041;
wire n_9634;
wire n_17846;
wire n_5876;
wire n_10916;
wire n_8584;
wire n_11557;
wire n_17113;
wire n_16748;
wire n_15363;
wire n_7810;
wire n_14955;
wire n_9364;
wire n_8228;
wire n_1825;
wire n_16015;
wire n_170;
wire n_15642;
wire n_1412;
wire n_10929;
wire n_18854;
wire n_19372;
wire n_13862;
wire n_8100;
wire n_13446;
wire n_13086;
wire n_8091;
wire n_5837;
wire n_148;
wire n_4675;
wire n_17155;
wire n_5491;
wire n_2987;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_12787;
wire n_12799;
wire n_4002;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_15205;
wire n_8158;
wire n_1295;
wire n_8469;
wire n_18718;
wire n_18481;
wire n_10102;
wire n_5983;
wire n_3146;
wire n_1438;
wire n_3953;
wire n_11825;
wire n_1100;
wire n_14354;
wire n_7684;
wire n_15532;
wire n_5604;
wire n_673;
wire n_16083;
wire n_10589;
wire n_11611;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_865;
wire n_4191;
wire n_18221;
wire n_12408;
wire n_16287;
wire n_16169;
wire n_19314;
wire n_17556;
wire n_2341;
wire n_10110;
wire n_11230;
wire n_11688;
wire n_4350;
wire n_12715;
wire n_12434;
wire n_11709;
wire n_14328;
wire n_6095;
wire n_17049;
wire n_18938;
wire n_16540;
wire n_14429;
wire n_12979;
wire n_16901;
wire n_6559;
wire n_3924;
wire n_15799;
wire n_19733;
wire n_17195;
wire n_19050;
wire n_4621;
wire n_510;
wire n_1488;
wire n_2148;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_2339;
wire n_10190;
wire n_19656;
wire n_5984;
wire n_6287;
wire n_13614;
wire n_8347;
wire n_17703;
wire n_19440;
wire n_1766;
wire n_1776;
wire n_14208;
wire n_9330;
wire n_4021;
wire n_3014;
wire n_15693;
wire n_12029;
wire n_4103;
wire n_9523;
wire n_14584;
wire n_4022;
wire n_19636;
wire n_10060;
wire n_18192;
wire n_9686;
wire n_4481;
wire n_17130;
wire n_19375;
wire n_1304;
wire n_10162;
wire n_4669;
wire n_15002;
wire n_9964;
wire n_17515;
wire n_13842;
wire n_7510;
wire n_6662;
wire n_11291;
wire n_9154;
wire n_5603;
wire n_13107;
wire n_14501;
wire n_3312;
wire n_7109;
wire n_2936;
wire n_3224;
wire n_8822;
wire n_14790;
wire n_1087;
wire n_17204;
wire n_12187;
wire n_657;
wire n_19662;
wire n_18772;
wire n_1505;
wire n_7253;
wire n_3129;
wire n_17201;
wire n_8476;
wire n_17745;
wire n_11927;
wire n_16674;
wire n_16326;
wire n_16571;
wire n_8359;
wire n_4484;
wire n_15808;
wire n_16497;
wire n_16752;
wire n_14574;
wire n_526;
wire n_14451;
wire n_2251;
wire n_9455;
wire n_8708;
wire n_14092;
wire n_2837;
wire n_4883;
wire n_14509;
wire n_11882;
wire n_17649;
wire n_11647;
wire n_15027;
wire n_15404;
wire n_10706;
wire n_3341;
wire n_19129;
wire n_8872;
wire n_19746;
wire n_3559;
wire n_8238;
wire n_15465;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_5146;
wire n_3056;
wire n_745;
wire n_15858;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_18946;
wire n_2589;
wire n_4535;
wire n_14765;
wire n_7704;
wire n_18893;
wire n_16170;
wire n_14995;
wire n_6302;
wire n_2442;
wire n_17479;
wire n_7203;
wire n_11259;
wire n_7670;
wire n_18258;
wire n_16010;
wire n_9673;
wire n_14434;
wire n_2545;
wire n_8642;
wire n_11875;
wire n_18567;
wire n_12111;
wire n_8912;
wire n_19067;
wire n_1314;
wire n_864;
wire n_14275;
wire n_19309;
wire n_12903;
wire n_6343;
wire n_12593;
wire n_5270;
wire n_1534;
wire n_17849;
wire n_11602;
wire n_15689;
wire n_12413;
wire n_17474;
wire n_723;
wire n_13813;
wire n_16190;
wire n_8111;
wire n_18315;
wire n_10432;
wire n_19227;
wire n_16888;
wire n_8056;
wire n_18376;
wire n_3287;
wire n_9674;
wire n_2357;
wire n_6433;
wire n_18253;
wire n_15469;
wire n_17140;
wire n_18407;
wire n_1681;
wire n_520;
wire n_18816;
wire n_4020;
wire n_13636;
wire n_19332;
wire n_19456;
wire n_5220;
wire n_18920;
wire n_11341;
wire n_10787;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_16308;
wire n_6279;
wire n_13905;
wire n_12290;
wire n_7881;
wire n_9369;
wire n_18896;
wire n_16986;
wire n_17872;
wire n_6071;
wire n_9583;
wire n_19422;
wire n_15119;
wire n_19117;
wire n_12150;
wire n_1617;
wire n_3370;
wire n_335;
wire n_15256;
wire n_18366;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_15982;
wire n_274;
wire n_19643;
wire n_18647;
wire n_15452;
wire n_1267;
wire n_1806;
wire n_13615;
wire n_15625;
wire n_2023;
wire n_12633;
wire n_14779;
wire n_496;
wire n_15114;
wire n_4614;
wire n_3360;
wire n_10277;
wire n_17934;
wire n_3956;
wire n_8163;
wire n_16632;
wire n_16028;
wire n_10948;
wire n_10525;
wire n_14287;
wire n_9507;
wire n_11528;
wire n_15296;
wire n_15828;
wire n_18107;
wire n_19211;
wire n_3870;
wire n_16126;
wire n_18102;
wire n_19699;
wire n_18545;
wire n_16168;
wire n_15915;
wire n_793;
wire n_10049;
wire n_3749;
wire n_15551;
wire n_9457;
wire n_5780;
wire n_5037;
wire n_16738;
wire n_316;
wire n_6084;
wire n_11039;
wire n_14342;
wire n_2555;
wire n_13693;
wire n_18992;
wire n_12606;
wire n_10900;
wire n_2201;
wire n_14107;
wire n_14781;
wire n_13333;
wire n_13229;
wire n_994;
wire n_17336;
wire n_11380;
wire n_15737;
wire n_19567;
wire n_10792;
wire n_15573;
wire n_13296;
wire n_14611;
wire n_3448;
wire n_17863;
wire n_1036;
wire n_1661;
wire n_5360;
wire n_17088;
wire n_19100;
wire n_15051;
wire n_6548;
wire n_3926;
wire n_6993;
wire n_1095;
wire n_15916;
wire n_4405;
wire n_16468;
wire n_10241;
wire n_19598;
wire n_15639;
wire n_3670;
wire n_179;
wire n_4667;
wire n_8702;
wire n_17158;
wire n_8116;
wire n_1115;
wire n_7946;
wire n_8195;
wire n_14069;
wire n_18452;
wire n_19786;
wire n_1409;
wire n_9991;
wire n_11366;
wire n_11872;
wire n_10823;
wire n_19685;
wire n_14766;
wire n_11106;
wire n_1126;
wire n_14592;
wire n_15109;
wire n_11132;
wire n_17625;
wire n_18546;
wire n_18034;
wire n_3635;
wire n_18181;
wire n_17126;
wire n_10824;
wire n_4155;
wire n_19566;
wire n_16216;
wire n_19398;
wire n_14277;
wire n_19565;
wire n_13493;
wire n_16389;
wire n_9047;
wire n_12842;
wire n_18569;
wire n_12481;
wire n_18168;
wire n_11316;
wire n_9599;
wire n_11559;
wire n_9072;
wire n_4929;
wire n_9428;
wire n_10340;
wire n_17463;
wire n_15817;
wire n_15344;
wire n_2220;
wire n_2577;
wire n_13669;
wire n_17245;
wire n_3529;
wire n_17179;
wire n_11109;
wire n_13840;
wire n_16601;
wire n_11591;
wire n_19710;
wire n_14251;
wire n_11225;
wire n_6765;
wire n_4565;
wire n_4159;
wire n_8883;
wire n_10634;
wire n_4586;
wire n_11058;
wire n_15888;
wire n_1608;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_3628;
wire n_14679;
wire n_10961;
wire n_7357;
wire n_1491;
wire n_17064;
wire n_8737;
wire n_13925;
wire n_18334;
wire n_10379;
wire n_16704;
wire n_2586;
wire n_18223;
wire n_13368;
wire n_14507;
wire n_9484;
wire n_10989;
wire n_17725;
wire n_10939;
wire n_19557;
wire n_1046;
wire n_2560;
wire n_1145;
wire n_11144;
wire n_14857;
wire n_6406;
wire n_14034;
wire n_10962;
wire n_11128;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_12007;
wire n_11025;
wire n_5062;
wire n_15901;
wire n_321;
wire n_13481;
wire n_12018;
wire n_3588;
wire n_18040;
wire n_17393;
wire n_14457;
wire n_16931;
wire n_12872;
wire n_18189;
wire n_6492;
wire n_14517;
wire n_2288;
wire n_11460;
wire n_13713;
wire n_12372;
wire n_13608;
wire n_7046;
wire n_19059;
wire n_10956;
wire n_2642;
wire n_7468;
wire n_2383;
wire n_18785;
wire n_14934;
wire n_19663;
wire n_2351;
wire n_18844;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_2986;
wire n_19752;
wire n_17870;
wire n_139;
wire n_15652;
wire n_3489;
wire n_19466;
wire n_16713;
wire n_14578;
wire n_15653;
wire n_5914;
wire n_12955;
wire n_9321;
wire n_16856;
wire n_18555;
wire n_1282;
wire n_15016;
wire n_2567;
wire n_18493;
wire n_275;
wire n_3377;
wire n_9161;
wire n_2869;
wire n_7836;
wire n_10737;
wire n_17910;
wire n_17750;
wire n_346;
wire n_15865;
wire n_13448;
wire n_16928;
wire n_5813;
wire n_13767;
wire n_790;
wire n_2611;
wire n_2901;
wire n_11055;
wire n_4358;
wire n_16616;
wire n_14832;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_17599;
wire n_14571;
wire n_6631;
wire n_12369;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_8927;
wire n_17985;
wire n_16396;
wire n_17531;
wire n_15155;
wire n_12686;
wire n_6228;
wire n_19336;
wire n_5416;
wire n_14881;
wire n_18588;
wire n_14527;
wire n_12822;
wire n_13307;
wire n_7279;
wire n_17460;
wire n_13312;
wire n_11761;
wire n_9984;
wire n_8474;
wire n_3524;
wire n_489;
wire n_2885;
wire n_10600;
wire n_6102;
wire n_636;
wire n_10833;
wire n_18329;
wire n_18649;
wire n_13023;
wire n_19343;
wire n_1607;
wire n_1454;
wire n_15315;
wire n_19210;
wire n_11185;
wire n_13440;
wire n_869;
wire n_1154;
wire n_13436;
wire n_19615;
wire n_19133;
wire n_16982;
wire n_846;
wire n_841;
wire n_508;
wire n_11081;
wire n_16687;
wire n_1562;
wire n_14858;
wire n_8787;
wire n_13911;
wire n_5051;
wire n_17544;
wire n_5587;
wire n_10941;
wire n_14617;
wire n_9816;
wire n_17132;
wire n_14263;
wire n_661;
wire n_8605;
wire n_10358;
wire n_3565;
wire n_17593;
wire n_9944;
wire n_6998;
wire n_16158;
wire n_4173;
wire n_12338;
wire n_7615;
wire n_5651;
wire n_9605;
wire n_1217;
wire n_7591;
wire n_11404;
wire n_16488;
wire n_15994;
wire n_15685;
wire n_9788;
wire n_16273;
wire n_10785;
wire n_18262;
wire n_13872;
wire n_17646;
wire n_12341;
wire n_18389;
wire n_5412;
wire n_14475;
wire n_10815;
wire n_1120;
wire n_555;
wire n_8784;
wire n_7382;
wire n_2048;
wire n_13955;
wire n_176;
wire n_17708;
wire n_14400;
wire n_4857;
wire n_16725;
wire n_16904;
wire n_16432;
wire n_12085;
wire n_2883;
wire n_18190;
wire n_13554;
wire n_18421;
wire n_863;
wire n_6780;
wire n_11582;
wire n_3268;
wire n_1147;
wire n_1754;
wire n_11705;
wire n_3701;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_17391;
wire n_19782;
wire n_17682;
wire n_7282;
wire n_9968;
wire n_11474;
wire n_10657;
wire n_13595;
wire n_5997;
wire n_2492;
wire n_10687;
wire n_13283;
wire n_19543;
wire n_15615;
wire n_12110;
wire n_8363;
wire n_5119;
wire n_19445;
wire n_17802;
wire n_9669;
wire n_17775;
wire n_6510;
wire n_8282;
wire n_5938;
wire n_15972;
wire n_6237;
wire n_12216;
wire n_11752;
wire n_12040;
wire n_17446;
wire n_2117;
wire n_18573;
wire n_14975;
wire n_7581;
wire n_6360;
wire n_17960;
wire n_15217;
wire n_4858;
wire n_13308;
wire n_19049;
wire n_9952;
wire n_15323;
wire n_12183;
wire n_10668;
wire n_9256;
wire n_5750;
wire n_4823;
wire n_4309;
wire n_839;
wire n_14007;
wire n_7346;
wire n_1537;
wire n_13373;
wire n_4243;
wire n_7428;
wire n_12221;
wire n_5666;
wire n_9195;
wire n_16236;
wire n_17787;
wire n_7283;
wire n_4142;
wire n_6314;
wire n_10632;
wire n_18861;
wire n_9623;
wire n_3796;
wire n_6964;
wire n_3408;
wire n_19027;
wire n_19561;
wire n_1184;
wire n_18912;
wire n_19322;
wire n_16702;
wire n_1525;
wire n_2594;
wire n_11329;
wire n_5994;
wire n_6495;
wire n_17280;
wire n_9516;
wire n_4244;
wire n_2147;
wire n_13241;
wire n_16027;
wire n_2503;
wire n_8976;
wire n_17844;
wire n_18136;
wire n_10130;
wire n_11661;
wire n_9222;
wire n_8435;
wire n_8882;
wire n_16391;
wire n_4787;
wire n_15949;
wire n_10622;
wire n_5633;
wire n_5664;
wire n_6797;
wire n_15673;
wire n_14012;
wire n_8759;
wire n_16941;
wire n_7177;
wire n_357;
wire n_13066;
wire n_13665;
wire n_12993;
wire n_19604;
wire n_11314;
wire n_17784;
wire n_2681;
wire n_15678;
wire n_8235;
wire n_13083;
wire n_3764;
wire n_19093;
wire n_16164;
wire n_6152;
wire n_16444;
wire n_4075;
wire n_9820;
wire n_14071;
wire n_12749;
wire n_2303;
wire n_1619;
wire n_8448;
wire n_4538;
wire n_12066;
wire n_6513;
wire n_2367;
wire n_1034;
wire n_15908;
wire n_754;
wire n_11184;
wire n_11945;
wire n_11368;
wire n_6330;
wire n_17842;
wire n_19628;
wire n_8457;
wire n_19200;
wire n_18605;
wire n_18837;
wire n_9339;
wire n_14312;
wire n_9601;
wire n_15045;
wire n_11409;
wire n_18995;
wire n_2107;
wire n_2040;
wire n_18737;
wire n_12437;
wire n_5624;
wire n_10840;
wire n_6263;
wire n_10515;
wire n_15501;
wire n_6490;
wire n_15751;
wire n_11605;
wire n_1861;
wire n_10242;
wire n_10144;
wire n_9684;
wire n_15741;
wire n_16195;
wire n_14793;
wire n_18754;
wire n_13472;
wire n_2162;
wire n_15596;
wire n_207;
wire n_4763;
wire n_3587;
wire n_205;
wire n_18316;
wire n_6038;
wire n_15379;
wire n_16272;
wire n_14884;
wire n_3162;
wire n_8964;
wire n_16629;
wire n_1899;
wire n_9814;
wire n_4804;
wire n_5619;
wire n_5859;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_4500;
wire n_13443;
wire n_4433;
wire n_5644;
wire n_2813;
wire n_14626;
wire n_2027;
wire n_2091;
wire n_8960;
wire n_5030;
wire n_15402;
wire n_4194;
wire n_18026;
wire n_8443;
wire n_7715;
wire n_2419;
wire n_8683;
wire n_18558;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_3182;
wire n_5756;
wire n_15306;
wire n_15981;
wire n_16367;

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_29),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_8),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_49),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_40),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_83),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_21),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_42),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_72),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_3),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_25),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_27),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_54),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_59),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_16),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_119),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_70),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_52),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_0),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_6),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_67),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_45),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_92),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_58),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_69),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_41),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_51),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_39),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_23),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_61),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_93),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_18),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_65),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_81),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_33),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_0),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_77),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_44),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_47),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_132),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_28),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_73),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_60),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_37),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_35),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_38),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_80),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_112),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_63),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_32),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_99),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_68),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_7),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_94),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_76),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_110),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_31),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_15),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_84),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_56),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_86),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_109),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_122),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_50),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_30),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_91),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_146),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_148),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_185),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_154),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_135),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_155),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_136),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_156),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_138),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_165),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_137),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_12),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_157),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_166),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_170),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_140),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_141),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_183),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_142),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_144),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_184),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_153),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_169),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_145),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_182),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_193),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_177),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_169),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_205),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_211),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_224),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_280),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_272),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_297),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_267),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_273),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_188),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_278),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_270),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_281),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_286),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_287),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_289),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_290),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_291),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_295),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_306),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_206),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_239),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_254),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_307),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_267),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_267),
.B(n_221),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_280),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_348),
.A2(n_178),
.B(n_195),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_225),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_158),
.B(n_256),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_149),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_346),
.B(n_191),
.Y(n_368)
);

OAI22x1_ASAP7_75t_SL g369 ( 
.A1(n_335),
.A2(n_264),
.B1(n_263),
.B2(n_204),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

AND2x2_ASAP7_75t_SL g371 ( 
.A(n_329),
.B(n_147),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_177),
.Y(n_373)
);

OA22x2_ASAP7_75t_SL g374 ( 
.A1(n_325),
.A2(n_247),
.B1(n_231),
.B2(n_241),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_198),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_209),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

OAI22x1_ASAP7_75t_SL g386 ( 
.A1(n_310),
.A2(n_223),
.B1(n_253),
.B2(n_240),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_191),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_340),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_322),
.A2(n_257),
.B1(n_252),
.B2(n_251),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_150),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_325),
.A2(n_236),
.B(n_230),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_347),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_347),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_324),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_265),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_318),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_314),
.B(n_246),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_309),
.Y(n_420)
);

CKINVDCx6p67_ASAP7_75t_R g421 ( 
.A(n_329),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_309),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_329),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_325),
.A2(n_232),
.B(n_262),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_309),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_317),
.B(n_212),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_314),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_325),
.A2(n_208),
.B(n_260),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_314),
.B(n_207),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_309),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_314),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_317),
.B(n_212),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_317),
.B(n_202),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_314),
.B(n_201),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_353),
.B(n_214),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_325),
.A2(n_210),
.B(n_259),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_320),
.B(n_200),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_331),
.B(n_197),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_314),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_318),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_309),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_318),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_329),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_346),
.A2(n_213),
.B1(n_258),
.B2(n_255),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_320),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_309),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_346),
.A2(n_192),
.B1(n_249),
.B2(n_245),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_309),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_309),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_320),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_329),
.B(n_214),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_309),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_309),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_346),
.B(n_189),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_318),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_331),
.B(n_187),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_318),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_324),
.B(n_196),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_347),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_335),
.A2(n_180),
.B1(n_244),
.B2(n_243),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_331),
.B(n_179),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_347),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_317),
.B(n_261),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_309),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_309),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_347),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_309),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_317),
.B(n_176),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_318),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_317),
.B(n_242),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_317),
.B(n_175),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_318),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_314),
.B(n_174),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_318),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_317),
.B(n_238),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_309),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_318),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_318),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_173),
.B1(n_235),
.B2(n_234),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_357),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_366),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_172),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_380),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_406),
.B(n_171),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_365),
.B(n_237),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_362),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_390),
.B(n_168),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_361),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_477),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_480),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_375),
.B(n_214),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_428),
.B(n_167),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_412),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_SL g523 ( 
.A(n_398),
.B(n_215),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_164),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_444),
.B(n_216),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_360),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_370),
.B(n_163),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_429),
.B(n_436),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_469),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_363),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_377),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_393),
.B(n_96),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_376),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_407),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_377),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_438),
.B(n_217),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_359),
.B(n_218),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_382),
.B(n_162),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_382),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_429),
.B(n_219),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_423),
.B(n_161),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_379),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_392),
.B(n_220),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_411),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_471),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_358),
.A2(n_160),
.B(n_228),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_396),
.B(n_106),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_434),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_453),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_467),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_394),
.B(n_123),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_456),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_459),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_385),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_475),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_470),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_389),
.B(n_152),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_474),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_385),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_484),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_431),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_395),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_478),
.B(n_159),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_479),
.B(n_222),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_419),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_430),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_408),
.B(n_439),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_442),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_374),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_457),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_443),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_441),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_483),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_367),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_454),
.A2(n_226),
.B(n_229),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_481),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_458),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_400),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_404),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_465),
.B(n_436),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_451),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_445),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_373),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_445),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_373),
.B(n_368),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_401),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_397),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_402),
.B(n_399),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_371),
.B(n_468),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_403),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_416),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_415),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_421),
.A2(n_386),
.B(n_369),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_378),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_391),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_381),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_405),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_357),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_417),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_365),
.B(n_428),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_417),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_435),
.B(n_461),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_370),
.B(n_381),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_370),
.B(n_381),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_461),
.B(n_435),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_365),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_417),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_381),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_461),
.B(n_435),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_357),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_365),
.B(n_428),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_357),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_381),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_357),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_398),
.B(n_368),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_357),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_381),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_357),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_357),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_357),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_381),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_417),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_365),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_357),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g652 ( 
.A(n_398),
.B(n_368),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_357),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_405),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_375),
.B(n_393),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_381),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_461),
.B(n_435),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_357),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_357),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_417),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_405),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_435),
.B(n_461),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_381),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_370),
.B(n_381),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_357),
.Y(n_665)
);

BUFx8_ASAP7_75t_L g666 ( 
.A(n_403),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_405),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_381),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_357),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_357),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_381),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_381),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_461),
.B(n_435),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_365),
.B(n_428),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_381),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_357),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_417),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_357),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_381),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_357),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_381),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_357),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_357),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_365),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_381),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_405),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_365),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_405),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_405),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_357),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_398),
.B(n_368),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_381),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_357),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_365),
.B(n_428),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_405),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_405),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_357),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_381),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_357),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_435),
.A2(n_461),
.B1(n_390),
.B2(n_359),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_435),
.B(n_390),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_381),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_405),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_357),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_381),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_381),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_381),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_461),
.B(n_435),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_375),
.B(n_393),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_357),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_370),
.B(n_381),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_357),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_417),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_381),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_405),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_358),
.A2(n_410),
.B(n_364),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_381),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_461),
.A2(n_375),
.B1(n_435),
.B2(n_359),
.Y(n_718)
);

XNOR2xp5_ASAP7_75t_L g719 ( 
.A(n_416),
.B(n_310),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_405),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_357),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_365),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_461),
.B(n_435),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_417),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_405),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_405),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_381),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_357),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_405),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_435),
.B(n_461),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_365),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_435),
.B(n_390),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_357),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_405),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_357),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_357),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_357),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_423),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_461),
.B(n_435),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_405),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_417),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_357),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_381),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_461),
.B(n_435),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_370),
.B(n_381),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_405),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_461),
.B(n_435),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_357),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_365),
.B(n_428),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_405),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_405),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_381),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_423),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_398),
.B(n_368),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_381),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_365),
.B(n_428),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_381),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_370),
.B(n_381),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_381),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_357),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_365),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_405),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_357),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_357),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_381),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_381),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_357),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_357),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_370),
.B(n_381),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_370),
.B(n_381),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_357),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_357),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_435),
.B(n_461),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_357),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_357),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_357),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_365),
.B(n_428),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_405),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_357),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_435),
.B(n_461),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_417),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_405),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_461),
.A2(n_375),
.B1(n_435),
.B2(n_359),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_357),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_381),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_357),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_357),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_357),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_370),
.B(n_381),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_405),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_SL g791 ( 
.A1(n_400),
.A2(n_293),
.B1(n_297),
.B2(n_280),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_357),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_487),
.Y(n_793)
);

BUFx4f_ASAP7_75t_L g794 ( 
.A(n_487),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_490),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_629),
.B(n_662),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_730),
.A2(n_780),
.B1(n_773),
.B2(n_530),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_590),
.B(n_592),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_493),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_R g800 ( 
.A(n_738),
.B(n_753),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_491),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_608),
.A2(n_595),
.B1(n_600),
.B2(n_632),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_495),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_636),
.B(n_657),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_514),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_491),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_515),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_498),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_R g809 ( 
.A(n_604),
.B(n_583),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_673),
.B(n_708),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_503),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_624),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_739),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_624),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_504),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_661),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_661),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_655),
.B(n_709),
.Y(n_818)
);

AND2x6_ASAP7_75t_L g819 ( 
.A(n_594),
.B(n_627),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_505),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_SL g821 ( 
.A1(n_791),
.A2(n_605),
.B1(n_719),
.B2(n_618),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_744),
.B(n_747),
.Y(n_822)
);

AND2x2_ASAP7_75t_SL g823 ( 
.A(n_613),
.B(n_654),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_686),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_686),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_SL g826 ( 
.A1(n_506),
.A2(n_510),
.B(n_509),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_512),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_513),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_516),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_688),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_688),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_650),
.B(n_761),
.C(n_684),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_529),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_625),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_637),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_689),
.Y(n_836)
);

BUFx8_ASAP7_75t_SL g837 ( 
.A(n_613),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_689),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_718),
.A2(n_783),
.B1(n_616),
.B2(n_599),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_703),
.Y(n_841)
);

OAI21xp33_ASAP7_75t_L g842 ( 
.A1(n_519),
.A2(n_524),
.B(n_638),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_639),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_720),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_641),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_557),
.B(n_585),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_643),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_645),
.Y(n_848)
);

BUFx6f_ASAP7_75t_SL g849 ( 
.A(n_720),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_646),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_647),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_651),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_499),
.B(n_700),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_532),
.B(n_538),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_725),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_501),
.B(n_596),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_734),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_653),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_633),
.B(n_687),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_658),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_722),
.B(n_731),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_734),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_659),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_667),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_750),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_665),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_526),
.B(n_540),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_588),
.B(n_589),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_750),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_669),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_670),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_674),
.B(n_694),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_532),
.B(n_538),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_676),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_782),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_680),
.A2(n_683),
.B1(n_690),
.B2(n_682),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_782),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_666),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_693),
.Y(n_880)
);

INVx5_ASAP7_75t_L g881 ( 
.A(n_790),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_541),
.B(n_749),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_597),
.A2(n_792),
.B1(n_697),
.B2(n_699),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_756),
.B(n_777),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_621),
.B(n_695),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_704),
.B(n_710),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_494),
.B(n_701),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_712),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_721),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_728),
.B(n_733),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_735),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_732),
.B(n_615),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_547),
.B(n_574),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_696),
.B(n_715),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_736),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_547),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_726),
.B(n_729),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_737),
.B(n_742),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_740),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_751),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_554),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_748),
.A2(n_771),
.B1(n_788),
.B2(n_787),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_760),
.B(n_763),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_764),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_574),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_581),
.B(n_606),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_767),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_768),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_772),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_774),
.B(n_775),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_776),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_746),
.B(n_762),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_779),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_784),
.Y(n_915)
);

OAI22xp33_ASAP7_75t_L g916 ( 
.A1(n_786),
.A2(n_612),
.B1(n_603),
.B2(n_601),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_581),
.B(n_614),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_489),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_492),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_488),
.B(n_500),
.C(n_523),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_496),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_778),
.B(n_619),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_655),
.B(n_709),
.Y(n_923)
);

XOR2x2_ASAP7_75t_L g924 ( 
.A(n_550),
.B(n_607),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_617),
.B(n_622),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_623),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_635),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_640),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_655),
.B(n_709),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_644),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_554),
.Y(n_931)
);

BUFx4f_ASAP7_75t_L g932 ( 
.A(n_587),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_648),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_656),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_518),
.A2(n_672),
.B1(n_671),
.B2(n_668),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_642),
.B(n_691),
.C(n_652),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_561),
.B(n_587),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_518),
.A2(n_707),
.B1(n_785),
.B2(n_766),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_630),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_598),
.A2(n_579),
.B1(n_586),
.B2(n_525),
.Y(n_940)
);

AND2x6_ASAP7_75t_L g941 ( 
.A(n_610),
.B(n_591),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_663),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_544),
.Y(n_943)
);

AND2x6_ASAP7_75t_L g944 ( 
.A(n_609),
.B(n_611),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_518),
.B(n_552),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_626),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_628),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_602),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_631),
.B(n_664),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_675),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_711),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_754),
.B(n_745),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_SL g953 ( 
.A1(n_551),
.A2(n_533),
.B1(n_560),
.B2(n_528),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_679),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_681),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_634),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_593),
.B(n_502),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_685),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_649),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_692),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_698),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_702),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_705),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_706),
.Y(n_964)
);

OA22x2_ASAP7_75t_L g965 ( 
.A1(n_620),
.A2(n_789),
.B1(n_758),
.B2(n_770),
.Y(n_965)
);

AND2x2_ASAP7_75t_SL g966 ( 
.A(n_549),
.B(n_769),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_714),
.B(n_755),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_717),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_727),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_743),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_752),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_757),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_759),
.Y(n_973)
);

AND2x6_ASAP7_75t_L g974 ( 
.A(n_517),
.B(n_562),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_660),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_677),
.Y(n_976)
);

NOR2x1p5_ASAP7_75t_L g977 ( 
.A(n_713),
.B(n_781),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_765),
.B(n_497),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_584),
.B(n_548),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_527),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_520),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_531),
.B(n_555),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_536),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_724),
.B(n_741),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_580),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_537),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_539),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_542),
.B(n_556),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_543),
.A2(n_573),
.B1(n_559),
.B2(n_569),
.Y(n_989)
);

INVxp33_ASAP7_75t_L g990 ( 
.A(n_521),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_565),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_570),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_571),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_572),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_576),
.A2(n_577),
.B1(n_582),
.B2(n_511),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_533),
.B(n_560),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_507),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_508),
.B(n_522),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_534),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_535),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_546),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_553),
.B(n_566),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_563),
.B(n_567),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_533),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_564),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_575),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_578),
.B(n_545),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_716),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_568),
.B(n_560),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_558),
.B(n_629),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_629),
.B(n_662),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_632),
.B(n_636),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_629),
.B(n_662),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_629),
.B(n_662),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_L g1015 ( 
.A(n_654),
.B(n_421),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_490),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_487),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_487),
.Y(n_1018)
);

INVx8_ASAP7_75t_L g1019 ( 
.A(n_554),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_632),
.B(n_636),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_654),
.B(n_554),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_514),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_487),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_490),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_514),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_629),
.B(n_730),
.C(n_662),
.Y(n_1026)
);

BUFx8_ASAP7_75t_SL g1027 ( 
.A(n_738),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_490),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_SL g1029 ( 
.A1(n_608),
.A2(n_662),
.B(n_629),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_738),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_487),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_487),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_514),
.Y(n_1033)
);

BUFx4f_ASAP7_75t_L g1034 ( 
.A(n_487),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_632),
.B(n_636),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_487),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_629),
.B(n_662),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_514),
.Y(n_1038)
);

BUFx4f_ASAP7_75t_L g1039 ( 
.A(n_487),
.Y(n_1039)
);

INVx6_ASAP7_75t_L g1040 ( 
.A(n_554),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_632),
.B(n_636),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_629),
.B(n_662),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_632),
.B(n_636),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_514),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_487),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_490),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_514),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_629),
.B(n_662),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_R g1049 ( 
.A(n_604),
.B(n_583),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_490),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_SL g1051 ( 
.A1(n_629),
.A2(n_730),
.B1(n_773),
.B2(n_662),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_629),
.B(n_662),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_514),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_629),
.B(n_662),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_583),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_514),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_487),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_514),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_487),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_632),
.B(n_636),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_487),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_487),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_629),
.B(n_662),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_487),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_514),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_SL g1066 ( 
.A(n_616),
.B(n_415),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_514),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_632),
.B(n_636),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_490),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_514),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_490),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_490),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_487),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_490),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_487),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_654),
.B(n_415),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_613),
.B(n_654),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_629),
.B(n_662),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_487),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_487),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_490),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_490),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_490),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_655),
.B(n_709),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_738),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_514),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_490),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_514),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_514),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_629),
.A2(n_662),
.B1(n_773),
.B2(n_730),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_487),
.Y(n_1091)
);

NOR2x1p5_ASAP7_75t_L g1092 ( 
.A(n_654),
.B(n_421),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_629),
.A2(n_662),
.B1(n_773),
.B2(n_730),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_487),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_632),
.B(n_636),
.Y(n_1095)
);

AND2x6_ASAP7_75t_L g1096 ( 
.A(n_590),
.B(n_592),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_487),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_490),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_629),
.A2(n_662),
.B1(n_773),
.B2(n_730),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_487),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_632),
.B(n_636),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_632),
.A2(n_708),
.B1(n_636),
.B2(n_673),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_487),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_487),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_487),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_632),
.B(n_636),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_654),
.B(n_554),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_SL g1108 ( 
.A(n_613),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_629),
.B(n_662),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_583),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_490),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_487),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_583),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_490),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_514),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_487),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_487),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_514),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_629),
.A2(n_662),
.B1(n_773),
.B2(n_730),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_632),
.B(n_636),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_514),
.Y(n_1121)
);

AND2x6_ASAP7_75t_L g1122 ( 
.A(n_590),
.B(n_592),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_490),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_490),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_487),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_629),
.B(n_662),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_490),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_490),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_613),
.B(n_654),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_629),
.B(n_662),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_490),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_487),
.Y(n_1132)
);

AO22x1_ASAP7_75t_L g1133 ( 
.A1(n_629),
.A2(n_730),
.B1(n_773),
.B2(n_662),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_629),
.B(n_662),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_490),
.Y(n_1135)
);

BUFx10_ASAP7_75t_L g1136 ( 
.A(n_529),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_490),
.Y(n_1137)
);

INVx8_ASAP7_75t_L g1138 ( 
.A(n_554),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_632),
.B(n_636),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_613),
.B(n_654),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_629),
.B(n_662),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_529),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_514),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_490),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_487),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_629),
.B(n_662),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_487),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_629),
.B(n_662),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_490),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_490),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_629),
.B(n_662),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_583),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_490),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_514),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_487),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_514),
.Y(n_1156)
);

AND2x6_ASAP7_75t_L g1157 ( 
.A(n_590),
.B(n_592),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_490),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_490),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_487),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_514),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_514),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_514),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_629),
.A2(n_662),
.B1(n_773),
.B2(n_730),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_490),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_514),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_632),
.B(n_636),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_514),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_514),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_514),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_487),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_487),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_490),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_487),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_490),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_487),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_514),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_490),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_487),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_487),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_490),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_490),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_487),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_490),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_514),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_490),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_629),
.B(n_662),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_514),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_487),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_487),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_487),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_629),
.B(n_662),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_514),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_629),
.B(n_662),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_490),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_490),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_616),
.B(n_415),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_490),
.Y(n_1198)
);

XNOR2xp5_ASAP7_75t_L g1199 ( 
.A(n_719),
.B(n_310),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_629),
.B(n_730),
.C(n_662),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_514),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_514),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_629),
.B(n_662),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_514),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_583),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_629),
.B(n_662),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_629),
.B(n_662),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_629),
.B(n_662),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_629),
.A2(n_730),
.B1(n_773),
.B2(n_662),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_514),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_487),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_490),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_L g1213 ( 
.A(n_629),
.B(n_730),
.C(n_662),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_654),
.B(n_554),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_487),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_514),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_514),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_487),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_487),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_487),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_490),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_629),
.B(n_662),
.Y(n_1222)
);

AND2x2_ASAP7_75t_SL g1223 ( 
.A(n_613),
.B(n_329),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_629),
.B(n_662),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_514),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_490),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_490),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_629),
.B(n_662),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_514),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_632),
.B(n_636),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_487),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_514),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_632),
.B(n_636),
.Y(n_1233)
);

AND2x2_ASAP7_75t_SL g1234 ( 
.A(n_613),
.B(n_329),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_490),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_629),
.B(n_662),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_490),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_487),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_632),
.B(n_636),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_629),
.B(n_662),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_632),
.B(n_636),
.Y(n_1241)
);

INVx6_ASAP7_75t_L g1242 ( 
.A(n_554),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1102),
.B(n_797),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_813),
.B(n_1013),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_859),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_810),
.B(n_822),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1109),
.B(n_1192),
.C(n_1148),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_796),
.B(n_1078),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_795),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1051),
.B(n_1041),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1194),
.B(n_1207),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_808),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_799),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1209),
.B(n_1090),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1208),
.B(n_1236),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_L g1256 ( 
.A(n_853),
.B(n_1213),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1240),
.B(n_1011),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_803),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1014),
.B(n_1037),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1110),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1261)
);

AO221x1_ASAP7_75t_L g1262 ( 
.A1(n_1119),
.A2(n_839),
.B1(n_916),
.B2(n_883),
.C(n_940),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1026),
.B(n_1200),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1076),
.B(n_932),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_881),
.B(n_1036),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1052),
.B(n_1054),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1063),
.B(n_1126),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1141),
.B(n_1151),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1187),
.B(n_1206),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1093),
.B(n_1164),
.C(n_1099),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1222),
.B(n_1224),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_868),
.B(n_1228),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1130),
.B(n_1134),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_815),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_893),
.B(n_888),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1146),
.B(n_1203),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1133),
.B(n_804),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1012),
.B(n_1020),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1035),
.B(n_1043),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_820),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1060),
.B(n_1068),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_811),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_872),
.B(n_885),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_SL g1285 ( 
.A(n_1223),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_828),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_861),
.Y(n_1287)
);

NOR3xp33_ASAP7_75t_L g1288 ( 
.A(n_821),
.B(n_842),
.C(n_1066),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1106),
.A2(n_1120),
.B1(n_1167),
.B2(n_1139),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_827),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_902),
.B(n_881),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1230),
.B(n_1233),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1239),
.B(n_1241),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_867),
.B(n_1029),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_802),
.B(n_882),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_887),
.B(n_891),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_L g1297 ( 
.A(n_923),
.B(n_929),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_856),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_829),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1197),
.A2(n_957),
.B1(n_920),
.B2(n_846),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_823),
.B(n_1004),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_812),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1108),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_SL g1304 ( 
.A(n_1234),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_812),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_899),
.B(n_904),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_834),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_847),
.A2(n_863),
.B1(n_871),
.B2(n_848),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_817),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_911),
.B(n_835),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1004),
.B(n_925),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1036),
.B(n_1059),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_843),
.B(n_845),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1019),
.B(n_1138),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_850),
.B(n_851),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_922),
.B(n_953),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_832),
.B(n_903),
.C(n_877),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_852),
.B(n_858),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_860),
.B(n_866),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_870),
.B(n_876),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_874),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_895),
.B(n_913),
.C(n_898),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_880),
.B(n_889),
.Y(n_1323)
);

INVxp33_ASAP7_75t_L g1324 ( 
.A(n_1152),
.Y(n_1324)
);

NOR3xp33_ASAP7_75t_L g1325 ( 
.A(n_952),
.B(n_1113),
.C(n_1055),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_892),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_896),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1205),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_910),
.B(n_912),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_890),
.B(n_905),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_908),
.B(n_909),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1016),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1024),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_809),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1059),
.B(n_1021),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_864),
.B(n_900),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_SL g1337 ( 
.A(n_837),
.B(n_1027),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1028),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1049),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1077),
.B(n_1129),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_886),
.Y(n_1341)
);

AO221x1_ASAP7_75t_L g1342 ( 
.A1(n_869),
.A2(n_1176),
.B1(n_824),
.B2(n_830),
.C(n_814),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_914),
.B(n_915),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1046),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_805),
.A2(n_1022),
.B1(n_1025),
.B2(n_807),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1077),
.B(n_1129),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_794),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1050),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_SL g1349 ( 
.A(n_1107),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_928),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_901),
.B(n_990),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1005),
.B(n_1199),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1030),
.B(n_1085),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1069),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_826),
.B(n_989),
.C(n_1071),
.Y(n_1355)
);

BUFx5_ASAP7_75t_L g1356 ( 
.A(n_798),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1081),
.B(n_1083),
.C(n_1082),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1040),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1023),
.B(n_1031),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1094),
.B(n_1100),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1087),
.B(n_1098),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_SL g1363 ( 
.A(n_1019),
.B(n_1138),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_L g1364 ( 
.A(n_1214),
.B(n_936),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_SL g1365 ( 
.A(n_937),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_817),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_930),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_933),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_934),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_939),
.B(n_951),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1111),
.B(n_1114),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_950),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_960),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1123),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1105),
.B(n_1179),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_L g1376 ( 
.A(n_819),
.B(n_941),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_949),
.B(n_1218),
.C(n_1183),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1116),
.B(n_1172),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1124),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_964),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1131),
.B(n_1135),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1242),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1137),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_939),
.B(n_951),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_966),
.B(n_937),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_943),
.B(n_946),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_L g1388 ( 
.A(n_819),
.B(n_941),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_947),
.B(n_956),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1150),
.B(n_1153),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_857),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1140),
.B(n_977),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1034),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1165),
.B(n_1173),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1175),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_836),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1178),
.B(n_1181),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_968),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1186),
.B(n_1195),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1196),
.B(n_1198),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_959),
.B(n_985),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1212),
.B(n_1221),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_836),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1226),
.B(n_1227),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1039),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1140),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1235),
.B(n_1237),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_L g1411 ( 
.A(n_819),
.B(n_941),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_857),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_978),
.B(n_1033),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_984),
.B(n_981),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_SL g1415 ( 
.A(n_833),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_969),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1001),
.B(n_1231),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_840),
.B(n_841),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_965),
.A2(n_849),
.B1(n_996),
.B2(n_1155),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1056),
.B(n_1058),
.Y(n_1422)
);

BUFx5_ASAP7_75t_L g1423 ( 
.A(n_798),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1065),
.B(n_1067),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1007),
.B(n_1084),
.C(n_818),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_840),
.B(n_841),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1070),
.B(n_1086),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_970),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_865),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_971),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1009),
.A2(n_982),
.B1(n_988),
.B2(n_1229),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_865),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_L g1433 ( 
.A(n_801),
.B(n_838),
.C(n_831),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1010),
.A2(n_945),
.B1(n_1121),
.B2(n_1232),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1088),
.B(n_1089),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_875),
.B(n_1017),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_875),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1017),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1045),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_972),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1045),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1143),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1064),
.B(n_1097),
.Y(n_1444)
);

XOR2xp5_ASAP7_75t_L g1445 ( 
.A(n_879),
.B(n_924),
.Y(n_1445)
);

BUFx5_ASAP7_75t_L g1446 ( 
.A(n_798),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1064),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1154),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1097),
.B(n_1145),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1156),
.B(n_1161),
.Y(n_1450)
);

NOR3xp33_ASAP7_75t_L g1451 ( 
.A(n_844),
.B(n_1180),
.C(n_1174),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1162),
.B(n_1163),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1166),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_992),
.Y(n_1454)
);

INVxp33_ASAP7_75t_L g1455 ( 
.A(n_800),
.Y(n_1455)
);

XOR2xp5_ASAP7_75t_L g1456 ( 
.A(n_995),
.B(n_1238),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1145),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_967),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1168),
.B(n_1169),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_SL g1460 ( 
.A(n_931),
.B(n_806),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1155),
.B(n_1220),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1170),
.B(n_1177),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1185),
.Y(n_1463)
);

NOR3xp33_ASAP7_75t_L g1464 ( 
.A(n_862),
.B(n_1171),
.C(n_1132),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1188),
.B(n_1193),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1201),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1202),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1204),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1210),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1216),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1220),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_SL g1472 ( 
.A(n_816),
.B(n_825),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_855),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1217),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1225),
.B(n_980),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1238),
.B(n_884),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_983),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_878),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_986),
.A2(n_987),
.B1(n_991),
.B2(n_994),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_993),
.B(n_918),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_997),
.B(n_919),
.Y(n_1481)
);

NOR3xp33_ASAP7_75t_L g1482 ( 
.A(n_1018),
.B(n_1219),
.C(n_1061),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1032),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1062),
.B(n_1215),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1002),
.B(n_1190),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_921),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_926),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1075),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1073),
.B(n_1189),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_927),
.B(n_955),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_942),
.B(n_973),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_954),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_958),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_961),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_962),
.B(n_963),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1079),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1003),
.B(n_979),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1006),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1080),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_999),
.B(n_1000),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_998),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_907),
.B(n_935),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_974),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1160),
.Y(n_1504)
);

NOR2x1p5_ASAP7_75t_L g1505 ( 
.A(n_1191),
.B(n_1112),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_SL g1506 ( 
.A(n_1136),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_938),
.B(n_944),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_L g1508 ( 
.A(n_944),
.B(n_974),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1104),
.B(n_1125),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1008),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_974),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_917),
.B(n_976),
.C(n_975),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_L g1513 ( 
.A(n_1117),
.B(n_906),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1096),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_793),
.B(n_1057),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1091),
.B(n_1211),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1096),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_897),
.B(n_1103),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1147),
.B(n_854),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_873),
.B(n_894),
.Y(n_1520)
);

NOR3xp33_ASAP7_75t_L g1521 ( 
.A(n_1142),
.B(n_1015),
.C(n_1092),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_975),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_944),
.B(n_1096),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1122),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1157),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_976),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1009),
.B(n_948),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_795),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_808),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1076),
.B(n_415),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_796),
.B(n_1078),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_808),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_813),
.B(n_1109),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1102),
.B(n_797),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_813),
.B(n_1109),
.Y(n_1540)
);

INVxp33_ASAP7_75t_L g1541 ( 
.A(n_856),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_813),
.B(n_1109),
.Y(n_1542)
);

AO221x1_ASAP7_75t_L g1543 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1102),
.B2(n_400),
.C(n_839),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1545)
);

BUFx5_ASAP7_75t_L g1546 ( 
.A(n_798),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_813),
.B(n_1109),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_795),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_795),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_813),
.B(n_1109),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1076),
.B(n_415),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_813),
.B(n_1109),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1102),
.B(n_797),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1102),
.B(n_797),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_837),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_881),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_808),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_808),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_813),
.B(n_1109),
.Y(n_1562)
);

NOR2xp67_ASAP7_75t_L g1563 ( 
.A(n_902),
.B(n_554),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_808),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1102),
.B(n_797),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_813),
.B(n_1109),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1102),
.B(n_797),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_813),
.B(n_1109),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_881),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1055),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_795),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_808),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_795),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_808),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_813),
.B(n_1109),
.Y(n_1575)
);

AO221x1_ASAP7_75t_L g1576 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1102),
.B2(n_400),
.C(n_839),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_808),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_902),
.B(n_554),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_813),
.B(n_1109),
.Y(n_1579)
);

NOR2x1p5_ASAP7_75t_L g1580 ( 
.A(n_902),
.B(n_397),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_796),
.B(n_1078),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_808),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1041),
.B(n_810),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_813),
.B(n_1109),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_813),
.B(n_1109),
.Y(n_1586)
);

INVxp33_ASAP7_75t_L g1587 ( 
.A(n_856),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1110),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1102),
.B(n_797),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_813),
.B(n_1109),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_813),
.B(n_1109),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_813),
.B(n_1109),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_795),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_796),
.B(n_1078),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_813),
.B(n_1109),
.Y(n_1596)
);

NOR2xp67_ASAP7_75t_L g1597 ( 
.A(n_902),
.B(n_554),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_813),
.B(n_1109),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_813),
.B(n_1109),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_837),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_795),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_808),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_796),
.B(n_1078),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_813),
.B(n_1109),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_808),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_L g1606 ( 
.A(n_902),
.B(n_554),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_813),
.B(n_1109),
.Y(n_1607)
);

NOR3xp33_ASAP7_75t_L g1608 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_795),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1102),
.B(n_797),
.Y(n_1611)
);

NAND2x1_ASAP7_75t_L g1612 ( 
.A(n_798),
.B(n_1096),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_813),
.B(n_1109),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_808),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1102),
.B(n_797),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1013),
.A2(n_1148),
.B1(n_1192),
.B2(n_1109),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_808),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1618)
);

NAND3xp33_ASAP7_75t_SL g1619 ( 
.A(n_1209),
.B(n_1099),
.C(n_1093),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_796),
.B(n_1078),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_796),
.B(n_1078),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1102),
.B(n_797),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_795),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_856),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_853),
.B(n_1213),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1076),
.B(n_415),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_859),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_932),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_L g1629 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_881),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_808),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_813),
.B(n_1109),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_881),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_932),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1102),
.B(n_797),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_795),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_796),
.B(n_1078),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_795),
.Y(n_1638)
);

NOR2xp67_ASAP7_75t_L g1639 ( 
.A(n_902),
.B(n_554),
.Y(n_1639)
);

INVxp33_ASAP7_75t_L g1640 ( 
.A(n_856),
.Y(n_1640)
);

NOR2xp67_ASAP7_75t_L g1641 ( 
.A(n_902),
.B(n_554),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_L g1642 ( 
.A(n_853),
.B(n_1213),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1102),
.B(n_797),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_813),
.B(n_1109),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_808),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_808),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_808),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_932),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_795),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_813),
.B(n_1109),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_795),
.Y(n_1652)
);

BUFx5_ASAP7_75t_L g1653 ( 
.A(n_798),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_795),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_813),
.B(n_1109),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_813),
.B(n_1109),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_813),
.B(n_1109),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1102),
.B(n_797),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_813),
.B(n_1109),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_795),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_881),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_813),
.B(n_1109),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_808),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_813),
.B(n_1109),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_795),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_813),
.B(n_1109),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_795),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_813),
.B(n_1109),
.Y(n_1670)
);

NOR2xp67_ASAP7_75t_L g1671 ( 
.A(n_902),
.B(n_554),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1013),
.B2(n_1148),
.C(n_1109),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_902),
.B(n_654),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_813),
.B(n_1109),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_813),
.B(n_1109),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_808),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_813),
.B(n_1109),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_813),
.B(n_1109),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_813),
.B(n_1109),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_932),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_881),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_796),
.B(n_1078),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_SL g1685 ( 
.A(n_1223),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_808),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_813),
.B(n_1109),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_932),
.Y(n_1688)
);

BUFx5_ASAP7_75t_L g1689 ( 
.A(n_798),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_795),
.Y(n_1690)
);

NOR2xp67_ASAP7_75t_L g1691 ( 
.A(n_902),
.B(n_554),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_808),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_813),
.B(n_1109),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1019),
.B(n_1138),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_813),
.B(n_1109),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_795),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1013),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1013),
.B2(n_1148),
.C(n_1109),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1699)
);

NOR3xp33_ASAP7_75t_L g1700 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_813),
.B(n_1109),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_808),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_813),
.B(n_1109),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1102),
.B(n_797),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1019),
.B(n_1138),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_808),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_796),
.B(n_1078),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1102),
.B(n_797),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1102),
.B(n_797),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_808),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_881),
.B(n_1036),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_813),
.B(n_1109),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1013),
.A2(n_1109),
.B1(n_1192),
.B2(n_1148),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_808),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_813),
.B(n_1109),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_795),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_813),
.B(n_1109),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_L g1719 ( 
.A(n_853),
.B(n_1213),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1102),
.B(n_797),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1110),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_813),
.B(n_1109),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1723)
);

AO221x1_ASAP7_75t_L g1724 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1102),
.B2(n_400),
.C(n_839),
.Y(n_1724)
);

AND2x6_ASAP7_75t_L g1725 ( 
.A(n_923),
.B(n_595),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_808),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_813),
.B(n_1109),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_808),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_932),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_808),
.Y(n_1731)
);

AND2x2_ASAP7_75t_SL g1732 ( 
.A(n_1213),
.B(n_1223),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_932),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_932),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_813),
.B(n_1109),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_932),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_813),
.B(n_1109),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_808),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_795),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_902),
.B(n_554),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_813),
.B(n_1109),
.Y(n_1743)
);

NOR2xp67_ASAP7_75t_L g1744 ( 
.A(n_902),
.B(n_554),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1102),
.B(n_797),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_808),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_932),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_813),
.B(n_1109),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_837),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_808),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1102),
.B(n_797),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_795),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1055),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_808),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1102),
.B(n_797),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_813),
.B(n_1109),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_795),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_796),
.B(n_1078),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_881),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_795),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_813),
.B(n_1109),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1110),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_837),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1102),
.B(n_797),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_813),
.B(n_1109),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_808),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_795),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_859),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_795),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_796),
.B(n_1078),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_808),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_932),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1102),
.B(n_797),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1102),
.B(n_797),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_796),
.B(n_1078),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_808),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1013),
.A2(n_1148),
.B1(n_1192),
.B2(n_1109),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_837),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_796),
.B(n_1078),
.Y(n_1779)
);

INVxp33_ASAP7_75t_L g1780 ( 
.A(n_856),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_813),
.B(n_1109),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1102),
.B(n_797),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_813),
.B(n_1109),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1008),
.A2(n_716),
.B(n_590),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1102),
.B(n_797),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1013),
.A2(n_1148),
.B1(n_1192),
.B2(n_1109),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_881),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1213),
.A2(n_1013),
.B1(n_1148),
.B2(n_1109),
.Y(n_1789)
);

NAND2x1p5_ASAP7_75t_L g1790 ( 
.A(n_881),
.B(n_1036),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_881),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_813),
.B(n_1109),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_808),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_808),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_795),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_796),
.B(n_1078),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_813),
.B(n_1109),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_SL g1799 ( 
.A(n_1209),
.B(n_1099),
.C(n_1093),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_808),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_808),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_808),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_795),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_795),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_808),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_808),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_813),
.B(n_1109),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_808),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_795),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1102),
.B(n_797),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_813),
.B(n_1109),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_808),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_R g1815 ( 
.A(n_1030),
.B(n_310),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_813),
.B(n_1109),
.Y(n_1816)
);

BUFx2_ASAP7_75t_R g1817 ( 
.A(n_837),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_795),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_813),
.B(n_1109),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1102),
.B(n_797),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_813),
.B(n_1109),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_813),
.B(n_1109),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_795),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1102),
.B(n_797),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_795),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_795),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_795),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_795),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_808),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_813),
.B(n_1109),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1102),
.B(n_797),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_813),
.B(n_1109),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_L g1834 ( 
.A(n_853),
.B(n_1213),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1027),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_808),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1102),
.B(n_797),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_932),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_813),
.B(n_1109),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_795),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_859),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1102),
.B(n_797),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_795),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1102),
.B(n_797),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_L g1846 ( 
.A(n_853),
.B(n_1213),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_932),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_932),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_859),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_795),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_796),
.B(n_1078),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1102),
.B(n_797),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_813),
.B(n_1109),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_813),
.B(n_1109),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_796),
.B(n_1078),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_808),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_795),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_813),
.B(n_1109),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_SL g1861 ( 
.A(n_1223),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_808),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1013),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_795),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_813),
.B(n_1109),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_808),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_795),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_813),
.B(n_1109),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1102),
.B(n_797),
.Y(n_1870)
);

OA21x2_ASAP7_75t_L g1871 ( 
.A1(n_1008),
.A2(n_716),
.B(n_590),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_SL g1872 ( 
.A(n_1223),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_808),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_795),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_797),
.A2(n_1209),
.B1(n_1099),
.B2(n_1164),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_932),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_881),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_813),
.B(n_1109),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_813),
.B(n_1109),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1102),
.B(n_797),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_813),
.B(n_1109),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_813),
.B(n_1109),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1102),
.B(n_797),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_813),
.B(n_1109),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_813),
.B(n_1109),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_932),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_932),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_813),
.B(n_1109),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_795),
.Y(n_1890)
);

NOR3xp33_ASAP7_75t_L g1891 ( 
.A(n_1090),
.B(n_1119),
.C(n_1109),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_795),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1102),
.B(n_797),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_813),
.B(n_1109),
.Y(n_1894)
);

INVxp67_ASAP7_75t_SL g1895 ( 
.A(n_1013),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1102),
.B(n_797),
.Y(n_1896)
);

INVx3_ASAP7_75t_R g1897 ( 
.A(n_1021),
.Y(n_1897)
);

BUFx5_ASAP7_75t_L g1898 ( 
.A(n_798),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1102),
.B(n_797),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_813),
.B(n_1109),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1102),
.B(n_797),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1102),
.B(n_797),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_813),
.B(n_1109),
.Y(n_1905)
);

NAND2x1p5_ASAP7_75t_L g1906 ( 
.A(n_881),
.B(n_1036),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_808),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_808),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_808),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_881),
.B(n_1036),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_808),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1102),
.B(n_797),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_813),
.B(n_1109),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_795),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_813),
.B(n_1109),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_881),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1090),
.A2(n_1119),
.B1(n_1013),
.B2(n_1148),
.C(n_1109),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_881),
.B(n_1036),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_813),
.B(n_1109),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1102),
.B(n_797),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_813),
.B(n_1109),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_837),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_L g1926 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_SL g1927 ( 
.A(n_1004),
.B(n_397),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_795),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_813),
.B(n_1109),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_813),
.B(n_1109),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1013),
.A2(n_1109),
.B1(n_1192),
.B2(n_1148),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1102),
.B(n_797),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_813),
.B(n_1109),
.Y(n_1934)
);

NAND3xp33_ASAP7_75t_L g1935 ( 
.A(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_795),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_796),
.B(n_1078),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1102),
.B(n_797),
.Y(n_1938)
);

OR2x6_ASAP7_75t_L g1939 ( 
.A(n_1019),
.B(n_1138),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_808),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1013),
.A2(n_1148),
.B1(n_1192),
.B2(n_1109),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1102),
.B(n_797),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1944)
);

AND2x6_ASAP7_75t_L g1945 ( 
.A(n_1514),
.B(n_1524),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1532),
.B(n_1551),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1612),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1302),
.Y(n_1948)
);

NOR2xp67_ASAP7_75t_L g1949 ( 
.A(n_1322),
.B(n_1334),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1396),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1711),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1626),
.B(n_1584),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1244),
.B(n_1538),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1249),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1248),
.B(n_1534),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1336),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1251),
.B(n_1255),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1537),
.A2(n_1608),
.B1(n_1649),
.B2(n_1629),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1253),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1547),
.B(n_1550),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1552),
.B(n_1562),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1294),
.A2(n_1306),
.B(n_1296),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1533),
.B(n_1536),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_SL g1965 ( 
.A(n_1340),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1258),
.Y(n_1966)
);

INVx4_ASAP7_75t_L g1967 ( 
.A(n_1711),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1672),
.B(n_1698),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1283),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1364),
.B(n_1346),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1575),
.B(n_1579),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1713),
.B(n_1545),
.C(n_1544),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1290),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1585),
.B(n_1586),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1299),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1560),
.A2(n_1583),
.B1(n_1660),
.B2(n_1618),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1593),
.A2(n_1598),
.B(n_1599),
.C(n_1596),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1604),
.B(n_1607),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1679),
.A2(n_1700),
.B1(n_1723),
.B2(n_1680),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1891),
.A2(n_1619),
.B1(n_1799),
.B2(n_1920),
.Y(n_1983)
);

INVx8_ASAP7_75t_L g1984 ( 
.A(n_1921),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1699),
.A2(n_1729),
.B1(n_1788),
.B2(n_1734),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1921),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1328),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1613),
.B(n_1632),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1644),
.B(n_1651),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1656),
.B(n_1657),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1658),
.B(n_1661),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1664),
.B(n_1666),
.Y(n_1992)
);

AOI22x1_ASAP7_75t_SL g1993 ( 
.A1(n_1836),
.A2(n_1863),
.B1(n_1895),
.B2(n_1697),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1668),
.B(n_1670),
.Y(n_1994)
);

AO22x1_ASAP7_75t_L g1995 ( 
.A1(n_1796),
.A2(n_1809),
.B1(n_1825),
.B2(n_1805),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1674),
.B(n_1675),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1677),
.B(n_1678),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1681),
.B(n_1687),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1307),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1332),
.Y(n_2000)
);

NAND2x1p5_ASAP7_75t_L g2001 ( 
.A(n_1927),
.B(n_1340),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1693),
.B(n_1695),
.Y(n_2002)
);

NOR2xp67_ASAP7_75t_L g2003 ( 
.A(n_1339),
.B(n_1245),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1333),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1701),
.B(n_1703),
.Y(n_2005)
);

OR2x6_ASAP7_75t_L g2006 ( 
.A(n_1314),
.B(n_1694),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1712),
.B(n_1716),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1817),
.B(n_1264),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1718),
.B(n_1722),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1338),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1815),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1727),
.B(n_1737),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1739),
.B(n_1743),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1852),
.B(n_1860),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1942),
.B(n_1616),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1733),
.Y(n_2016)
);

INVx8_ASAP7_75t_L g2017 ( 
.A(n_1365),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1748),
.B(n_1756),
.Y(n_2018)
);

OAI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1777),
.A2(n_1786),
.B1(n_1765),
.B2(n_1781),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1302),
.Y(n_2020)
);

INVx2_ASAP7_75t_SL g2021 ( 
.A(n_1772),
.Y(n_2021)
);

NAND2x1_ASAP7_75t_L g2022 ( 
.A(n_1517),
.B(n_1527),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1937),
.B(n_1581),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1761),
.B(n_1783),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1792),
.B(n_1798),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1808),
.B(n_1813),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1816),
.B(n_1819),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1821),
.B(n_1822),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1869),
.B(n_1879),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1351),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1831),
.B(n_1833),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1344),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1875),
.A2(n_1270),
.B1(n_1254),
.B2(n_1899),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1348),
.Y(n_2034)
);

INVx5_ASAP7_75t_L g2035 ( 
.A(n_1725),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1354),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1840),
.B(n_1854),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1876),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1901),
.A2(n_1907),
.B(n_1916),
.C(n_1912),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1303),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1855),
.B(n_1859),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1865),
.B(n_1868),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1374),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1932),
.B(n_1940),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1944),
.B(n_1878),
.Y(n_2045)
);

INVxp67_ASAP7_75t_L g2046 ( 
.A(n_1260),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1880),
.B(n_1882),
.Y(n_2047)
);

AND2x6_ASAP7_75t_SL g2048 ( 
.A(n_1353),
.B(n_1314),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1379),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1883),
.B(n_1885),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1543),
.A2(n_1724),
.B1(n_1576),
.B2(n_1789),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1356),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1247),
.A2(n_1610),
.B1(n_1654),
.B2(n_1588),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1384),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1397),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1628),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1275),
.A2(n_1539),
.B(n_1243),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1886),
.B(n_1889),
.Y(n_2058)
);

BUFx5_ASAP7_75t_L g2059 ( 
.A(n_1725),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1530),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_SL g2061 ( 
.A1(n_1894),
.A2(n_1905),
.B1(n_1915),
.B2(n_1902),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1548),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1918),
.B(n_1922),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_1393),
.B(n_1505),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1393),
.B(n_1386),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1924),
.B(n_1929),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_1595),
.B(n_1603),
.Y(n_2067)
);

BUFx12f_ASAP7_75t_L g2068 ( 
.A(n_1303),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1549),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1714),
.A2(n_1736),
.B1(n_1926),
.B2(n_1835),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1930),
.B(n_1934),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1931),
.B(n_1935),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_1553),
.A2(n_1554),
.B1(n_1567),
.B2(n_1565),
.Y(n_2073)
);

A2O1A1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_1256),
.A2(n_1642),
.B(n_1719),
.C(n_1625),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1571),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1573),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1620),
.B(n_1621),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1594),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1259),
.B(n_1261),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1257),
.A2(n_1267),
.B1(n_1271),
.B2(n_1269),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1601),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1609),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1266),
.B(n_1268),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1590),
.A2(n_1615),
.B(n_1611),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1637),
.B(n_1684),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1707),
.B(n_1758),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1770),
.B(n_1775),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1623),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1636),
.Y(n_2089)
);

AND2x6_ASAP7_75t_SL g2090 ( 
.A(n_1694),
.B(n_1705),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1779),
.B(n_1797),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1287),
.B(n_1627),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1851),
.B(n_1856),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1284),
.B(n_1273),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1288),
.A2(n_1834),
.B1(n_1846),
.B2(n_1250),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1276),
.B(n_1246),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1768),
.B(n_1842),
.Y(n_2097)
);

AND2x6_ASAP7_75t_SL g2098 ( 
.A(n_1705),
.B(n_1939),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_1622),
.A2(n_1635),
.B1(n_1659),
.B2(n_1643),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1638),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1497),
.A2(n_1708),
.B1(n_1709),
.B2(n_1704),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1849),
.B(n_1352),
.Y(n_2102)
);

NAND2xp33_ASAP7_75t_L g2103 ( 
.A(n_1425),
.B(n_1725),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1589),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1650),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_1720),
.A2(n_1745),
.B1(n_1755),
.B2(n_1751),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1652),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1272),
.B(n_1292),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_1721),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1263),
.B(n_1310),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1732),
.A2(n_1764),
.B1(n_1774),
.B2(n_1773),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1277),
.B(n_1782),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1295),
.B(n_1785),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1655),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1662),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1628),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_1812),
.B(n_1820),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_1824),
.A2(n_1832),
.B1(n_1843),
.B2(n_1838),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1414),
.B(n_1541),
.Y(n_2119)
);

BUFx8_ASAP7_75t_L g2120 ( 
.A(n_1349),
.Y(n_2120)
);

NAND2x1p5_ASAP7_75t_L g2121 ( 
.A(n_1301),
.B(n_1316),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_1381),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1845),
.B(n_1853),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1870),
.B(n_1881),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1285),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1884),
.B(n_1893),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1896),
.B(n_1900),
.Y(n_2127)
);

INVx8_ASAP7_75t_L g2128 ( 
.A(n_1939),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1356),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1356),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1903),
.B(n_1904),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1667),
.Y(n_2132)
);

NOR2xp67_ASAP7_75t_L g2133 ( 
.A(n_1341),
.B(n_1359),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1914),
.A2(n_1933),
.B1(n_1938),
.B2(n_1923),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1587),
.B(n_1624),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_1390),
.B(n_1391),
.Y(n_2136)
);

NAND2xp33_ASAP7_75t_L g2137 ( 
.A(n_1943),
.B(n_1356),
.Y(n_2137)
);

INVxp67_ASAP7_75t_L g2138 ( 
.A(n_1762),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1634),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1289),
.B(n_1278),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1279),
.B(n_1281),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1282),
.B(n_1293),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1458),
.B(n_1395),
.Y(n_2143)
);

INVx8_ASAP7_75t_L g2144 ( 
.A(n_1634),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1399),
.B(n_1413),
.Y(n_2145)
);

INVx4_ASAP7_75t_L g2146 ( 
.A(n_1648),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1648),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1300),
.B(n_1640),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1669),
.Y(n_2149)
);

NOR2x1p5_ASAP7_75t_L g2150 ( 
.A(n_1408),
.B(n_1555),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1427),
.B(n_1450),
.Y(n_2151)
);

NAND2xp33_ASAP7_75t_L g2152 ( 
.A(n_1423),
.B(n_1446),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1313),
.B(n_1315),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1780),
.B(n_1298),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1317),
.B(n_1324),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1570),
.B(n_1753),
.Y(n_2157)
);

AOI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_1355),
.A2(n_1431),
.B(n_1297),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1690),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1325),
.B(n_1419),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1423),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1308),
.A2(n_1358),
.B1(n_1479),
.B2(n_1323),
.Y(n_2162)
);

BUFx8_ASAP7_75t_L g2163 ( 
.A(n_1304),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1682),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1472),
.B(n_1460),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1696),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1320),
.B(n_1330),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1717),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1455),
.B(n_1456),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1741),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1331),
.B(n_1357),
.Y(n_2171)
);

INVx1_ASAP7_75t_SL g2172 ( 
.A(n_1473),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_1392),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1362),
.B(n_1371),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1382),
.B(n_1403),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1405),
.B(n_1407),
.Y(n_2176)
);

INVx5_ASAP7_75t_L g2177 ( 
.A(n_1682),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_1465),
.B(n_1410),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_1688),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_1688),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1752),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1757),
.B(n_1760),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1421),
.B(n_1435),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1767),
.B(n_1769),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1795),
.B(n_1803),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1804),
.B(n_1811),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1818),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1520),
.B(n_1401),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1823),
.B(n_1826),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1685),
.A2(n_1872),
.B1(n_1861),
.B2(n_1311),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_1402),
.B(n_1329),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1376),
.A2(n_1411),
.B(n_1388),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_1476),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1827),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1828),
.B(n_1829),
.Y(n_2195)
);

OR2x6_ASAP7_75t_L g2196 ( 
.A(n_1265),
.B(n_1790),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_1343),
.B(n_1485),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1435),
.B(n_1312),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1841),
.B(n_1844),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1850),
.B(n_1858),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1378),
.A2(n_1377),
.B1(n_1262),
.B2(n_1445),
.Y(n_2201)
);

NAND2xp33_ASAP7_75t_L g2202 ( 
.A(n_1423),
.B(n_1446),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1502),
.A2(n_1507),
.B(n_1784),
.Y(n_2203)
);

OR2x6_ASAP7_75t_L g2204 ( 
.A(n_1906),
.B(n_1911),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1252),
.B(n_1274),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_1423),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1864),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_1730),
.Y(n_2208)
);

NAND2x1p5_ASAP7_75t_L g2209 ( 
.A(n_1867),
.B(n_1874),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1890),
.B(n_1892),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1917),
.B(n_1928),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1936),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1409),
.B(n_1730),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1454),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_1345),
.A2(n_1529),
.B1(n_1280),
.B2(n_1321),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_1305),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1286),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1326),
.B(n_1327),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1531),
.B(n_1535),
.Y(n_2219)
);

NOR2x1p5_ASAP7_75t_L g2220 ( 
.A(n_1600),
.B(n_1749),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1558),
.B(n_1561),
.Y(n_2221)
);

O2A1O1Ixp5_ASAP7_75t_L g2222 ( 
.A1(n_1525),
.A2(n_1526),
.B(n_1491),
.C(n_1481),
.Y(n_2222)
);

AOI22xp33_ASAP7_75t_L g2223 ( 
.A1(n_1342),
.A2(n_1492),
.B1(n_1487),
.B2(n_1486),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1564),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1572),
.B(n_1574),
.Y(n_2225)
);

INVx8_ASAP7_75t_L g2226 ( 
.A(n_1735),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1577),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1582),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1602),
.B(n_1605),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1614),
.B(n_1617),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1735),
.Y(n_2231)
);

OAI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_1521),
.A2(n_1370),
.B1(n_1385),
.B2(n_1434),
.C(n_1519),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1631),
.B(n_1645),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1646),
.B(n_1647),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1665),
.B(n_1676),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1360),
.A2(n_1375),
.B1(n_1361),
.B2(n_1464),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1490),
.Y(n_2237)
);

NAND2x1p5_ASAP7_75t_L g2238 ( 
.A(n_1503),
.B(n_1511),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1495),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_SL g2240 ( 
.A1(n_1337),
.A2(n_1363),
.B1(n_1888),
.B2(n_1747),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1433),
.A2(n_1482),
.B1(n_1451),
.B2(n_1580),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1480),
.Y(n_2242)
);

A2O1A1Ixp33_ASAP7_75t_L g2243 ( 
.A1(n_1501),
.A2(n_1475),
.B(n_1913),
.C(n_1910),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1686),
.B(n_1692),
.Y(n_2244)
);

AND2x6_ASAP7_75t_SL g2245 ( 
.A(n_1515),
.B(n_1484),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_1493),
.A2(n_1494),
.B1(n_1909),
.B2(n_1908),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1702),
.B(n_1706),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1738),
.B(n_1747),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1710),
.B(n_1715),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1738),
.B(n_1839),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_1305),
.Y(n_2251)
);

OR2x6_ASAP7_75t_L g2252 ( 
.A(n_1839),
.B(n_1847),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1726),
.B(n_1728),
.Y(n_2253)
);

INVx4_ASAP7_75t_L g2254 ( 
.A(n_1847),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1731),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1740),
.B(n_1746),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_1504),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1750),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1754),
.B(n_1766),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_1771),
.B(n_1776),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_1848),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_L g2262 ( 
.A(n_1446),
.B(n_1546),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1793),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1794),
.B(n_1800),
.Y(n_2264)
);

OR2x6_ASAP7_75t_L g2265 ( 
.A(n_1848),
.B(n_1887),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_1801),
.B(n_1802),
.Y(n_2266)
);

BUFx8_ASAP7_75t_L g2267 ( 
.A(n_1415),
.Y(n_2267)
);

NOR3xp33_ASAP7_75t_L g2268 ( 
.A(n_1512),
.B(n_1422),
.C(n_1418),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1806),
.B(n_1807),
.Y(n_2269)
);

OAI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_1810),
.A2(n_1941),
.B1(n_1866),
.B2(n_1857),
.Y(n_2270)
);

O2A1O1Ixp5_ASAP7_75t_L g2271 ( 
.A1(n_1523),
.A2(n_1498),
.B(n_1510),
.C(n_1477),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_1887),
.B(n_1888),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1814),
.B(n_1830),
.Y(n_2273)
);

BUFx6f_ASAP7_75t_L g2274 ( 
.A(n_1309),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_1489),
.A2(n_1837),
.B1(n_1873),
.B2(n_1862),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1463),
.B(n_1467),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_1504),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_1469),
.B(n_1474),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1443),
.Y(n_2279)
);

AOI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_1448),
.A2(n_1468),
.B1(n_1470),
.B2(n_1466),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1453),
.B(n_1350),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_1417),
.A2(n_1459),
.B1(n_1452),
.B2(n_1462),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_1309),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1367),
.B(n_1368),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_1369),
.B(n_1372),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1424),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1440),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1373),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_1478),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_1380),
.B(n_1400),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1416),
.B(n_1428),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_1404),
.A2(n_1347),
.B1(n_1394),
.B2(n_1387),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1430),
.B(n_1441),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1500),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1509),
.B(n_1518),
.Y(n_2295)
);

AOI22x1_ASAP7_75t_L g2296 ( 
.A1(n_1412),
.A2(n_1528),
.B1(n_1442),
.B2(n_1522),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1389),
.B(n_1483),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_1432),
.B(n_1461),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1446),
.Y(n_2299)
);

AND2x2_ASAP7_75t_SL g2300 ( 
.A(n_1508),
.B(n_1784),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_1499),
.B(n_1496),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1488),
.B(n_1513),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_1438),
.B(n_1439),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1420),
.B(n_1444),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_1366),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1546),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1426),
.B(n_1449),
.Y(n_2307)
);

INVxp67_ASAP7_75t_SL g2308 ( 
.A(n_1546),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_1335),
.B(n_1366),
.Y(n_2309)
);

INVx2_ASAP7_75t_SL g2310 ( 
.A(n_1398),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1871),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1436),
.B(n_1457),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_L g2313 ( 
.A(n_1546),
.B(n_1653),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1471),
.B(n_1673),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1653),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1516),
.B(n_1429),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1653),
.Y(n_2317)
);

NAND2x1_ASAP7_75t_L g2318 ( 
.A(n_1871),
.B(n_1663),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1398),
.B(n_1406),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_1447),
.B(n_1437),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1653),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_1689),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_1383),
.B(n_1437),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_1689),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1406),
.B(n_1429),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1689),
.B(n_1898),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_1563),
.B(n_1606),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1689),
.B(n_1898),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_1556),
.B(n_1630),
.Y(n_2329)
);

OR2x6_ASAP7_75t_L g2330 ( 
.A(n_1763),
.B(n_1925),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_1569),
.B(n_1919),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1898),
.B(n_1291),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_1578),
.A2(n_1742),
.B1(n_1597),
.B2(n_1744),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_1778),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_1639),
.A2(n_1691),
.B1(n_1641),
.B2(n_1671),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_1633),
.B(n_1791),
.Y(n_2336)
);

NOR2x2_ASAP7_75t_L g2337 ( 
.A(n_1897),
.B(n_1683),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1898),
.B(n_1759),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1787),
.B(n_1877),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1506),
.B(n_1532),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1396),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_1612),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_1336),
.Y(n_2344)
);

BUFx4_ASAP7_75t_L g2345 ( 
.A(n_1817),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2350)
);

AOI22xp33_ASAP7_75t_SL g2351 ( 
.A1(n_1931),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1396),
.Y(n_2354)
);

AOI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1612),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_1711),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2362)
);

AND2x6_ASAP7_75t_SL g2363 ( 
.A(n_1353),
.B(n_937),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1396),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2367)
);

O2A1O1Ixp5_ASAP7_75t_L g2368 ( 
.A1(n_1243),
.A2(n_1539),
.B(n_1554),
.C(n_1553),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_1612),
.Y(n_2373)
);

OAI221xp5_ASAP7_75t_L g2374 ( 
.A1(n_1713),
.A2(n_1099),
.B1(n_1164),
.B2(n_1093),
.C(n_1051),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2375)
);

OAI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_1713),
.A2(n_1099),
.B1(n_1164),
.B2(n_1093),
.C(n_1051),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1396),
.Y(n_2379)
);

INVx2_ASAP7_75t_SL g2380 ( 
.A(n_1711),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1396),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_1815),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1396),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1396),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1396),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1396),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2394)
);

O2A1O1Ixp5_ASAP7_75t_L g2395 ( 
.A1(n_1243),
.A2(n_1539),
.B(n_1554),
.C(n_1553),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1396),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1396),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2402)
);

OR2x6_ASAP7_75t_L g2403 ( 
.A(n_1340),
.B(n_937),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_1711),
.Y(n_2405)
);

NOR2xp67_ASAP7_75t_SL g2406 ( 
.A(n_1628),
.B(n_554),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1396),
.Y(n_2411)
);

AOI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1396),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1396),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1396),
.Y(n_2418)
);

INVx5_ASAP7_75t_L g2419 ( 
.A(n_1725),
.Y(n_2419)
);

OR2x6_ASAP7_75t_L g2420 ( 
.A(n_1340),
.B(n_937),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1815),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2423)
);

AND2x6_ASAP7_75t_L g2424 ( 
.A(n_1514),
.B(n_1524),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2425)
);

OAI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2427)
);

INVx4_ASAP7_75t_L g2428 ( 
.A(n_1711),
.Y(n_2428)
);

BUFx4f_ASAP7_75t_L g2429 ( 
.A(n_1628),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_1260),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1396),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1396),
.Y(n_2437)
);

NOR2xp67_ASAP7_75t_L g2438 ( 
.A(n_1322),
.B(n_554),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1396),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_1336),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2443)
);

O2A1O1Ixp33_ASAP7_75t_L g2444 ( 
.A1(n_1244),
.A2(n_1119),
.B(n_1090),
.C(n_1109),
.Y(n_2444)
);

AOI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1396),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1396),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2448)
);

AOI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_1711),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1396),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1396),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2455)
);

INVxp67_ASAP7_75t_L g2456 ( 
.A(n_1336),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_L g2458 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_L g2459 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2459)
);

OAI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2460)
);

NAND3xp33_ASAP7_75t_L g2461 ( 
.A(n_1713),
.B(n_1109),
.C(n_1013),
.Y(n_2461)
);

NAND2xp33_ASAP7_75t_L g2462 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_1612),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1396),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1396),
.Y(n_2470)
);

NAND2xp33_ASAP7_75t_L g2471 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2472)
);

NAND2xp33_ASAP7_75t_L g2473 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2473)
);

NAND2xp33_ASAP7_75t_L g2474 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_1612),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_1815),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_1711),
.Y(n_2478)
);

INVx4_ASAP7_75t_L g2479 ( 
.A(n_1711),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1396),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_1396),
.Y(n_2486)
);

OAI22xp33_ASAP7_75t_SL g2487 ( 
.A1(n_1244),
.A2(n_1540),
.B1(n_1542),
.B2(n_1538),
.Y(n_2487)
);

NOR2x1p5_ASAP7_75t_L g2488 ( 
.A(n_1733),
.B(n_421),
.Y(n_2488)
);

NOR2xp33_ASAP7_75t_L g2489 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1396),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_1612),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_1612),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_1396),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2501)
);

INVxp67_ASAP7_75t_L g2502 ( 
.A(n_1336),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_1396),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1396),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_1711),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1396),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_1396),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2518)
);

NOR2xp33_ASAP7_75t_L g2519 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_1815),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_1612),
.Y(n_2523)
);

INVx2_ASAP7_75t_SL g2524 ( 
.A(n_1711),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_1396),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1396),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2529)
);

A2O1A1Ixp33_ASAP7_75t_L g2530 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_2530)
);

NAND3xp33_ASAP7_75t_L g2531 ( 
.A(n_1713),
.B(n_1109),
.C(n_1013),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_1396),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1396),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2537)
);

AOI22xp33_ASAP7_75t_L g2538 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2538)
);

BUFx8_ASAP7_75t_L g2539 ( 
.A(n_1365),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2542)
);

AND2x4_ASAP7_75t_SL g2543 ( 
.A(n_1628),
.B(n_613),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1396),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_1396),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_1396),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2550)
);

AND2x2_ASAP7_75t_SL g2551 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2551)
);

BUFx3_ASAP7_75t_L g2552 ( 
.A(n_1711),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_1396),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_1711),
.Y(n_2556)
);

CKINVDCx20_ASAP7_75t_R g2557 ( 
.A(n_1815),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2559)
);

INVx2_ASAP7_75t_SL g2560 ( 
.A(n_1711),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_SL g2561 ( 
.A(n_1817),
.B(n_1532),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_1396),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_1396),
.Y(n_2563)
);

NAND2xp33_ASAP7_75t_L g2564 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_1396),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_1260),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_SL g2572 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2572)
);

INVxp67_ASAP7_75t_L g2573 ( 
.A(n_1336),
.Y(n_2573)
);

AOI21x1_ASAP7_75t_L g2574 ( 
.A1(n_1294),
.A2(n_1539),
.B(n_1243),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2577)
);

NOR3xp33_ASAP7_75t_L g2578 ( 
.A(n_1672),
.B(n_1119),
.C(n_1090),
.Y(n_2578)
);

AOI22xp33_ASAP7_75t_L g2579 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_1396),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_1396),
.Y(n_2582)
);

OR2x2_ASAP7_75t_L g2583 ( 
.A(n_1584),
.B(n_1041),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_1711),
.Y(n_2585)
);

OAI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_1713),
.A2(n_1099),
.B1(n_1164),
.B2(n_1093),
.C(n_1051),
.Y(n_2586)
);

NAND2x1p5_ASAP7_75t_L g2587 ( 
.A(n_1612),
.B(n_1004),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2588)
);

INVx4_ASAP7_75t_L g2589 ( 
.A(n_1711),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_1396),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_1711),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_1612),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_1396),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_1612),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_1396),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_1612),
.Y(n_2607)
);

A2O1A1Ixp33_ASAP7_75t_L g2608 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2609)
);

INVx2_ASAP7_75t_SL g2610 ( 
.A(n_1711),
.Y(n_2610)
);

AND2x6_ASAP7_75t_L g2611 ( 
.A(n_1514),
.B(n_1524),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1396),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2616)
);

NAND2x1p5_ASAP7_75t_L g2617 ( 
.A(n_1612),
.B(n_1004),
.Y(n_2617)
);

OR2x6_ASAP7_75t_L g2618 ( 
.A(n_1340),
.B(n_937),
.Y(n_2618)
);

INVx4_ASAP7_75t_L g2619 ( 
.A(n_1711),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_1396),
.Y(n_2620)
);

INVxp67_ASAP7_75t_L g2621 ( 
.A(n_1336),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_SL g2624 ( 
.A1(n_1931),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_2624)
);

NOR2xp67_ASAP7_75t_SL g2625 ( 
.A(n_1628),
.B(n_554),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_SL g2626 ( 
.A(n_1817),
.B(n_1532),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2630)
);

BUFx4f_ASAP7_75t_L g2631 ( 
.A(n_1628),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_1396),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_1396),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_1612),
.Y(n_2637)
);

NAND2xp33_ASAP7_75t_L g2638 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2639)
);

OAI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_1396),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_1396),
.Y(n_2644)
);

AOI22xp33_ASAP7_75t_L g2645 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_1396),
.Y(n_2647)
);

OR2x6_ASAP7_75t_L g2648 ( 
.A(n_1340),
.B(n_937),
.Y(n_2648)
);

OR2x6_ASAP7_75t_L g2649 ( 
.A(n_1340),
.B(n_937),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2651)
);

INVx2_ASAP7_75t_SL g2652 ( 
.A(n_1711),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_R g2654 ( 
.A(n_1532),
.B(n_310),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2656)
);

BUFx6f_ASAP7_75t_L g2657 ( 
.A(n_1612),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2661)
);

NAND2x1p5_ASAP7_75t_L g2662 ( 
.A(n_1612),
.B(n_1004),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2664)
);

NAND2x1p5_ASAP7_75t_L g2665 ( 
.A(n_1612),
.B(n_1004),
.Y(n_2665)
);

INVx4_ASAP7_75t_L g2666 ( 
.A(n_1711),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_1396),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2668)
);

INVx4_ASAP7_75t_L g2669 ( 
.A(n_1711),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2670)
);

INVx2_ASAP7_75t_SL g2671 ( 
.A(n_1711),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_1396),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_1396),
.Y(n_2676)
);

OA22x2_ASAP7_75t_L g2677 ( 
.A1(n_1616),
.A2(n_1209),
.B1(n_1786),
.B2(n_1777),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_1396),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_SL g2679 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_1396),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_1396),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2687)
);

AOI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_1396),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2691)
);

AOI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_1396),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2699)
);

INVx2_ASAP7_75t_SL g2700 ( 
.A(n_1711),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_1711),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_1584),
.B(n_1041),
.Y(n_2702)
);

NAND2xp33_ASAP7_75t_L g2703 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2705)
);

OAI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_SL g2710 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_1612),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_1336),
.Y(n_2715)
);

OR2x6_ASAP7_75t_L g2716 ( 
.A(n_1340),
.B(n_937),
.Y(n_2716)
);

NOR2xp67_ASAP7_75t_L g2717 ( 
.A(n_1322),
.B(n_554),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2718)
);

NOR3x1_ASAP7_75t_L g2719 ( 
.A(n_1247),
.B(n_1133),
.C(n_1119),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_SL g2721 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2721)
);

AND2x6_ASAP7_75t_SL g2722 ( 
.A(n_1353),
.B(n_937),
.Y(n_2722)
);

OR2x6_ASAP7_75t_L g2723 ( 
.A(n_1340),
.B(n_937),
.Y(n_2723)
);

AOI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2724)
);

INVx8_ASAP7_75t_L g2725 ( 
.A(n_1711),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2726)
);

BUFx3_ASAP7_75t_L g2727 ( 
.A(n_1711),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_1396),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2730)
);

NAND3xp33_ASAP7_75t_L g2731 ( 
.A(n_1713),
.B(n_1109),
.C(n_1013),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_1396),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_1396),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_1396),
.Y(n_2738)
);

INVx5_ASAP7_75t_L g2739 ( 
.A(n_1725),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_1396),
.Y(n_2740)
);

INVx3_ASAP7_75t_L g2741 ( 
.A(n_1612),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_1396),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_1396),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_1396),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2747)
);

NOR3xp33_ASAP7_75t_L g2748 ( 
.A(n_1672),
.B(n_1119),
.C(n_1090),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_1396),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_1396),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_1815),
.Y(n_2757)
);

NOR3xp33_ASAP7_75t_L g2758 ( 
.A(n_1672),
.B(n_1119),
.C(n_1090),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_1260),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_1815),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2766)
);

AOI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2768)
);

BUFx3_ASAP7_75t_L g2769 ( 
.A(n_1711),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2770)
);

BUFx3_ASAP7_75t_L g2771 ( 
.A(n_1711),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2772)
);

AND2x6_ASAP7_75t_SL g2773 ( 
.A(n_1353),
.B(n_937),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_1396),
.Y(n_2778)
);

INVxp67_ASAP7_75t_L g2779 ( 
.A(n_1336),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2780)
);

NOR2xp33_ASAP7_75t_L g2781 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_1612),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_1396),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_1815),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_SL g2787 ( 
.A1(n_1713),
.A2(n_1051),
.B1(n_1255),
.B2(n_1251),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_1711),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_SL g2789 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2793)
);

AND2x6_ASAP7_75t_SL g2794 ( 
.A(n_1353),
.B(n_937),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_SL g2796 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2796)
);

AND2x6_ASAP7_75t_SL g2797 ( 
.A(n_1353),
.B(n_937),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1396),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_1396),
.Y(n_2802)
);

AOI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2803)
);

NOR3xp33_ASAP7_75t_SL g2804 ( 
.A(n_1619),
.B(n_1119),
.C(n_1090),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_R g2806 ( 
.A(n_1532),
.B(n_310),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2807)
);

INVxp67_ASAP7_75t_L g2808 ( 
.A(n_1336),
.Y(n_2808)
);

AND2x4_ASAP7_75t_SL g2809 ( 
.A(n_1628),
.B(n_613),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2811)
);

OR2x6_ASAP7_75t_L g2812 ( 
.A(n_1340),
.B(n_937),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_1396),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2814)
);

A2O1A1Ixp33_ASAP7_75t_SL g2815 ( 
.A1(n_1537),
.A2(n_1010),
.B(n_1109),
.C(n_1013),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_1396),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2817)
);

AND2x2_ASAP7_75t_SL g2818 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_1396),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_1396),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2823)
);

NOR2xp67_ASAP7_75t_L g2824 ( 
.A(n_1322),
.B(n_554),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_1815),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_1396),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_1396),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_1396),
.Y(n_2830)
);

AND2x6_ASAP7_75t_L g2831 ( 
.A(n_1514),
.B(n_1524),
.Y(n_2831)
);

O2A1O1Ixp33_ASAP7_75t_L g2832 ( 
.A1(n_1244),
.A2(n_1119),
.B(n_1090),
.C(n_1109),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2833)
);

NAND3xp33_ASAP7_75t_SL g2834 ( 
.A(n_1616),
.B(n_1209),
.C(n_1051),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2835)
);

OAI22xp5_ASAP7_75t_SL g2836 ( 
.A1(n_1713),
.A2(n_1051),
.B1(n_1255),
.B2(n_1251),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_SL g2837 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_1396),
.Y(n_2839)
);

OR2x2_ASAP7_75t_L g2840 ( 
.A(n_1584),
.B(n_1041),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1396),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_1396),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_1396),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_1244),
.A2(n_797),
.B1(n_1209),
.B2(n_1099),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_1396),
.Y(n_2849)
);

A2O1A1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_2850)
);

AOI22xp33_ASAP7_75t_L g2851 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_1396),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_1396),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_1396),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_R g2856 ( 
.A(n_1532),
.B(n_310),
.Y(n_2856)
);

NAND2x1p5_ASAP7_75t_L g2857 ( 
.A(n_1612),
.B(n_1004),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_L g2858 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2858)
);

INVxp67_ASAP7_75t_L g2859 ( 
.A(n_1336),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2861)
);

AND2x6_ASAP7_75t_SL g2862 ( 
.A(n_1353),
.B(n_937),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2863)
);

INVx8_ASAP7_75t_L g2864 ( 
.A(n_1711),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_1396),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2870)
);

O2A1O1Ixp5_ASAP7_75t_L g2871 ( 
.A1(n_1243),
.A2(n_1539),
.B(n_1554),
.C(n_1553),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_1584),
.B(n_1041),
.Y(n_2872)
);

INVx4_ASAP7_75t_L g2873 ( 
.A(n_1711),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_1396),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_1672),
.B(n_1698),
.Y(n_2876)
);

AOI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2877)
);

O2A1O1Ixp5_ASAP7_75t_L g2878 ( 
.A1(n_1243),
.A2(n_1539),
.B(n_1554),
.C(n_1553),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2879)
);

A2O1A1Ixp33_ASAP7_75t_L g2880 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_2880)
);

INVx8_ASAP7_75t_L g2881 ( 
.A(n_1711),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_1612),
.Y(n_2883)
);

AOI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2884)
);

AO22x1_ASAP7_75t_L g2885 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_1396),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2892)
);

OR2x2_ASAP7_75t_L g2893 ( 
.A(n_1584),
.B(n_1041),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_2895)
);

NAND2x1_ASAP7_75t_L g2896 ( 
.A(n_1514),
.B(n_798),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2900)
);

INVx8_ASAP7_75t_L g2901 ( 
.A(n_1711),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_1711),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2903)
);

OAI21xp5_ASAP7_75t_L g2904 ( 
.A1(n_1243),
.A2(n_853),
.B(n_1539),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_1396),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_1815),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2913)
);

NAND2x1_ASAP7_75t_L g2914 ( 
.A(n_1514),
.B(n_798),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2915)
);

CKINVDCx6p67_ASAP7_75t_R g2916 ( 
.A(n_1408),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_1396),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_1396),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2921)
);

OAI22xp33_ASAP7_75t_L g2922 ( 
.A1(n_1616),
.A2(n_1786),
.B1(n_1942),
.B2(n_1777),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_1396),
.Y(n_2925)
);

O2A1O1Ixp5_ASAP7_75t_L g2926 ( 
.A1(n_1243),
.A2(n_1539),
.B(n_1554),
.C(n_1553),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2927)
);

NOR2xp33_ASAP7_75t_L g2928 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_1396),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_1396),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_1396),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_1396),
.Y(n_2934)
);

OAI22xp33_ASAP7_75t_L g2935 ( 
.A1(n_1616),
.A2(n_1786),
.B1(n_1942),
.B2(n_1777),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_1396),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_R g2937 ( 
.A(n_1532),
.B(n_310),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_SL g2938 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2939)
);

NOR2xp33_ASAP7_75t_L g2940 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_1396),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_1396),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2949)
);

OAI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_1243),
.A2(n_853),
.B(n_1539),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_1396),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2952)
);

AND2x2_ASAP7_75t_SL g2953 ( 
.A(n_1537),
.B(n_1608),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_1396),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_1396),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_1396),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_1396),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2966)
);

INVx3_ASAP7_75t_L g2967 ( 
.A(n_1612),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_1248),
.B(n_1534),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_SL g2971 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2971)
);

AND2x6_ASAP7_75t_SL g2972 ( 
.A(n_1353),
.B(n_937),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2973)
);

OA22x2_ASAP7_75t_L g2974 ( 
.A1(n_1616),
.A2(n_1209),
.B1(n_1786),
.B2(n_1777),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2975)
);

AND2x4_ASAP7_75t_L g2976 ( 
.A(n_1364),
.B(n_1393),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_1396),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_1396),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_R g2985 ( 
.A(n_1532),
.B(n_310),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_1251),
.B(n_1255),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_1396),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_1532),
.B(n_1551),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_1396),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_1396),
.Y(n_2991)
);

AOI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_1244),
.B(n_1538),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_2998)
);

AND2x6_ASAP7_75t_SL g2999 ( 
.A(n_1353),
.B(n_937),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_1396),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_SL g3001 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_SL g3004 ( 
.A1(n_1713),
.A2(n_1051),
.B1(n_1255),
.B2(n_1251),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_1396),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3007)
);

INVx2_ASAP7_75t_SL g3008 ( 
.A(n_1711),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_1294),
.A2(n_530),
.B(n_867),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_1396),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_1396),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_1396),
.Y(n_3012)
);

AOI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_1396),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_1364),
.B(n_1393),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_1251),
.B(n_1255),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_1251),
.B(n_1255),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_1396),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_1396),
.Y(n_3022)
);

AND2x2_ASAP7_75t_SL g3023 ( 
.A(n_1537),
.B(n_1608),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_1396),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_1396),
.Y(n_3029)
);

AO22x1_ASAP7_75t_L g3030 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_1396),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_SL g3033 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_1396),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_1251),
.B(n_1255),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_1248),
.B(n_1534),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_3042)
);

AOI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_3043)
);

AOI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_1396),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_1260),
.Y(n_3047)
);

NAND3xp33_ASAP7_75t_L g3048 ( 
.A(n_1713),
.B(n_1109),
.C(n_1013),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_1711),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3050)
);

INVx2_ASAP7_75t_SL g3051 ( 
.A(n_1711),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_1396),
.Y(n_3052)
);

HB1xp67_ASAP7_75t_L g3053 ( 
.A(n_1260),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_1251),
.B(n_1255),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_1251),
.B(n_1255),
.Y(n_3055)
);

BUFx3_ASAP7_75t_L g3056 ( 
.A(n_1711),
.Y(n_3056)
);

INVx4_ASAP7_75t_L g3057 ( 
.A(n_1711),
.Y(n_3057)
);

AOI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_1251),
.A2(n_1109),
.B1(n_1148),
.B2(n_1013),
.Y(n_3058)
);

A2O1A1Ixp33_ASAP7_75t_L g3059 ( 
.A1(n_1251),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_1248),
.B(n_1534),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_1396),
.Y(n_3065)
);

HB1xp67_ASAP7_75t_L g3066 ( 
.A(n_1260),
.Y(n_3066)
);

AOI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_1537),
.A2(n_1629),
.B1(n_1649),
.B2(n_1608),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_SL g3069 ( 
.A(n_1817),
.B(n_1532),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_1532),
.B(n_1551),
.Y(n_3070)
);

INVx4_ASAP7_75t_L g3071 ( 
.A(n_1711),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_1244),
.B(n_1538),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_1396),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3074)
);

OAI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3076)
);

A2O1A1Ixp33_ASAP7_75t_L g3077 ( 
.A1(n_2444),
.A2(n_2832),
.B(n_2461),
.C(n_2731),
.Y(n_3077)
);

NOR3xp33_ASAP7_75t_L g3078 ( 
.A(n_2834),
.B(n_3048),
.C(n_2531),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2052),
.Y(n_3079)
);

OAI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2371),
.A2(n_2385),
.B(n_2375),
.Y(n_3080)
);

OAI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_2375),
.A2(n_2389),
.B(n_2385),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2389),
.B(n_2509),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2311),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2509),
.B(n_2513),
.Y(n_3086)
);

O2A1O1Ixp33_ASAP7_75t_SL g3087 ( 
.A1(n_2513),
.A2(n_2604),
.B(n_2613),
.C(n_2606),
.Y(n_3087)
);

INVx3_ASAP7_75t_L g3088 ( 
.A(n_2052),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2578),
.A2(n_2758),
.B(n_2748),
.C(n_2608),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2467),
.A2(n_2522),
.B(n_2511),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2604),
.A2(n_2606),
.B1(n_2615),
.B2(n_2613),
.Y(n_3091)
);

A2O1A1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2578),
.A2(n_2758),
.B(n_2748),
.C(n_2634),
.Y(n_3092)
);

OAI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2615),
.A2(n_2712),
.B(n_2630),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2554),
.A2(n_2692),
.B(n_2684),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2630),
.A2(n_2714),
.B1(n_2721),
.B2(n_2712),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2756),
.A2(n_2777),
.B(n_2760),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_1958),
.B(n_1964),
.Y(n_3097)
);

AND2x4_ASAP7_75t_L g3098 ( 
.A(n_2074),
.B(n_2129),
.Y(n_3098)
);

OAI21xp33_ASAP7_75t_L g3099 ( 
.A1(n_2341),
.A2(n_2445),
.B(n_2412),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2803),
.A2(n_2895),
.B(n_2877),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_1964),
.B(n_1976),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_2431),
.Y(n_3102)
);

NAND2x1_ASAP7_75t_L g3103 ( 
.A(n_2073),
.B(n_2099),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_3009),
.A2(n_2084),
.B(n_2134),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2714),
.A2(n_2860),
.B(n_2721),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2860),
.A2(n_2876),
.B(n_2875),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_2804),
.B(n_2033),
.Y(n_3107)
);

OAI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2449),
.A2(n_2463),
.B1(n_2575),
.B2(n_2498),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_1976),
.B(n_2014),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2875),
.A2(n_2876),
.B(n_2904),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_2014),
.B(n_2029),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2950),
.A2(n_2123),
.B(n_2101),
.Y(n_3112)
);

A2O1A1Ixp33_ASAP7_75t_L g3113 ( 
.A1(n_2530),
.A2(n_2880),
.B(n_3059),
.C(n_2850),
.Y(n_3113)
);

OAI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2368),
.A2(n_2871),
.B(n_2395),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2123),
.A2(n_2113),
.B(n_2137),
.Y(n_3115)
);

INVx1_ASAP7_75t_SL g3116 ( 
.A(n_2109),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_2029),
.B(n_2044),
.Y(n_3117)
);

OAI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2878),
.A2(n_2926),
.B(n_1983),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2019),
.B(n_2061),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2113),
.A2(n_2057),
.B(n_2462),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2787),
.A2(n_2836),
.B1(n_3004),
.B2(n_2348),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2033),
.B(n_2112),
.Y(n_3122)
);

INVxp67_ASAP7_75t_SL g3123 ( 
.A(n_2122),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2112),
.B(n_2117),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2117),
.B(n_2126),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2471),
.A2(n_2474),
.B(n_2473),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2126),
.B(n_2019),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2300),
.Y(n_3128)
);

BUFx6f_ASAP7_75t_L g3129 ( 
.A(n_2035),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2564),
.A2(n_2703),
.B(n_2638),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2158),
.A2(n_2127),
.B(n_2124),
.Y(n_3131)
);

AOI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_2131),
.A2(n_2202),
.B(n_2152),
.Y(n_3132)
);

OAI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_1983),
.A2(n_2099),
.B(n_2073),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2080),
.B(n_2106),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2044),
.B(n_2348),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2106),
.B(n_2118),
.Y(n_3136)
);

NOR2xp67_ASAP7_75t_L g3137 ( 
.A(n_2095),
.B(n_2035),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2551),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2262),
.A2(n_2313),
.B(n_2118),
.Y(n_3139)
);

A2O1A1Ixp33_ASAP7_75t_L g3140 ( 
.A1(n_2374),
.A2(n_2376),
.B(n_2586),
.C(n_1980),
.Y(n_3140)
);

AOI21x1_ASAP7_75t_L g3141 ( 
.A1(n_2203),
.A2(n_2318),
.B(n_2140),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2358),
.B(n_2426),
.Y(n_3142)
);

OAI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_1959),
.A2(n_2352),
.B(n_1982),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2460),
.B(n_2640),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2706),
.B(n_2848),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2599),
.A2(n_2688),
.B1(n_2733),
.B2(n_2724),
.Y(n_3146)
);

AOI21x1_ASAP7_75t_L g3147 ( 
.A1(n_2015),
.A2(n_2148),
.B(n_2162),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2349),
.B(n_2353),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2128),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2153),
.A2(n_2167),
.B(n_2156),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2551),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2349),
.B(n_2353),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2804),
.B(n_2818),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2922),
.B(n_2935),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2487),
.B(n_2922),
.Y(n_3155)
);

OAI321xp33_ASAP7_75t_L g3156 ( 
.A1(n_2764),
.A2(n_2884),
.A3(n_2992),
.B1(n_2793),
.B2(n_2915),
.C(n_2866),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2171),
.A2(n_2175),
.B(n_2174),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2815),
.A2(n_2953),
.B(n_2818),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2815),
.A2(n_3023),
.B(n_2953),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2935),
.B(n_1979),
.Y(n_3160)
);

CKINVDCx10_ASAP7_75t_R g3161 ( 
.A(n_1965),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_1984),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2360),
.B(n_2369),
.Y(n_3163)
);

NOR3xp33_ASAP7_75t_L g3164 ( 
.A(n_2885),
.B(n_3030),
.C(n_1995),
.Y(n_3164)
);

NOR3xp33_ASAP7_75t_L g3165 ( 
.A(n_2039),
.B(n_2369),
.C(n_2360),
.Y(n_3165)
);

OR2x2_ASAP7_75t_L g3166 ( 
.A(n_1959),
.B(n_1982),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2111),
.B(n_2079),
.Y(n_3167)
);

BUFx8_ASAP7_75t_SL g3168 ( 
.A(n_2345),
.Y(n_3168)
);

NOR3xp33_ASAP7_75t_L g3169 ( 
.A(n_2383),
.B(n_2396),
.C(n_2394),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2352),
.B(n_2361),
.Y(n_3170)
);

HB1xp67_ASAP7_75t_L g3171 ( 
.A(n_2431),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2361),
.B(n_2388),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_1985),
.B(n_2083),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3174)
);

INVx2_ASAP7_75t_SL g3175 ( 
.A(n_1984),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3023),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2390),
.B(n_2439),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2122),
.A2(n_2458),
.B(n_2439),
.Y(n_3178)
);

NAND2x1p5_ASAP7_75t_L g3179 ( 
.A(n_2035),
.B(n_2419),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2383),
.B(n_2394),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_2458),
.A2(n_2507),
.B(n_2459),
.Y(n_3181)
);

AOI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_2459),
.A2(n_2538),
.B(n_2507),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2538),
.A2(n_2579),
.B(n_2576),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_SL g3184 ( 
.A(n_2561),
.B(n_2626),
.Y(n_3184)
);

NOR2xp67_ASAP7_75t_L g3185 ( 
.A(n_2035),
.B(n_2419),
.Y(n_3185)
);

OAI22xp5_ASAP7_75t_L g3186 ( 
.A1(n_2774),
.A2(n_2996),
.B1(n_3043),
.B2(n_2941),
.Y(n_3186)
);

OAI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2576),
.A2(n_2612),
.B(n_2579),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2612),
.B(n_2641),
.Y(n_3188)
);

OAI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2641),
.A2(n_2729),
.B(n_2645),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_2419),
.Y(n_3190)
);

INVx4_ASAP7_75t_L g3191 ( 
.A(n_2419),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2645),
.A2(n_2747),
.B(n_2729),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_1954),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_L g3194 ( 
.A(n_2396),
.B(n_2398),
.Y(n_3194)
);

AO21x2_ASAP7_75t_L g3195 ( 
.A1(n_2103),
.A2(n_2246),
.B(n_2270),
.Y(n_3195)
);

OAI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_3058),
.A2(n_2398),
.B1(n_2409),
.B2(n_2400),
.Y(n_3196)
);

AOI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_2747),
.A2(n_2767),
.B(n_2752),
.Y(n_3197)
);

OAI21xp33_ASAP7_75t_L g3198 ( 
.A1(n_2400),
.A2(n_2433),
.B(n_2409),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2752),
.B(n_2767),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_2433),
.A2(n_2451),
.B(n_2455),
.C(n_2443),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2780),
.A2(n_2799),
.B(n_2784),
.Y(n_3201)
);

AND2x2_ASAP7_75t_SL g3202 ( 
.A(n_2780),
.B(n_2784),
.Y(n_3202)
);

AND2x2_ASAP7_75t_SL g3203 ( 
.A(n_2799),
.B(n_2814),
.Y(n_3203)
);

HB1xp67_ASAP7_75t_L g3204 ( 
.A(n_2569),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_L g3205 ( 
.A(n_2443),
.B(n_2451),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2814),
.B(n_2851),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_2569),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_1960),
.Y(n_3208)
);

A2O1A1Ixp33_ASAP7_75t_L g3209 ( 
.A1(n_2455),
.A2(n_2480),
.B(n_2489),
.C(n_2481),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2480),
.A2(n_2481),
.B(n_2491),
.C(n_2489),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2851),
.B(n_2891),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_2891),
.A2(n_2961),
.B(n_2921),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2921),
.B(n_2961),
.Y(n_3213)
);

OAI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_2969),
.A2(n_3013),
.B(n_2998),
.Y(n_3214)
);

BUFx12f_ASAP7_75t_L g3215 ( 
.A(n_2040),
.Y(n_3215)
);

OAI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_2969),
.A2(n_3013),
.B(n_2998),
.Y(n_3216)
);

OAI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3042),
.A2(n_3045),
.B(n_3044),
.Y(n_3217)
);

AOI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_3042),
.A2(n_3045),
.B(n_3044),
.Y(n_3218)
);

OAI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3067),
.A2(n_2051),
.B(n_2677),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2051),
.B(n_2677),
.Y(n_3220)
);

OAI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_2457),
.A2(n_2491),
.B1(n_2519),
.B2(n_2517),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2457),
.B(n_2517),
.Y(n_3222)
);

AOI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3067),
.A2(n_2176),
.B(n_2151),
.Y(n_3223)
);

AND2x2_ASAP7_75t_SL g3224 ( 
.A(n_2072),
.B(n_2719),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_1953),
.B(n_1955),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_1961),
.B(n_1962),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2519),
.B(n_2520),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_1969),
.B(n_1972),
.Y(n_3228)
);

OAI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2974),
.A2(n_2070),
.B(n_2053),
.Y(n_3229)
);

O2A1O1Ixp33_ASAP7_75t_SL g3230 ( 
.A1(n_2042),
.A2(n_2071),
.B(n_2047),
.C(n_2110),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_1975),
.B(n_1978),
.Y(n_3231)
);

NOR2xp67_ASAP7_75t_L g3232 ( 
.A(n_2739),
.B(n_2237),
.Y(n_3232)
);

BUFx4_ASAP7_75t_SL g3233 ( 
.A(n_2252),
.Y(n_3233)
);

BUFx24_ASAP7_75t_L g3234 ( 
.A(n_2359),
.Y(n_3234)
);

AND2x2_ASAP7_75t_SL g3235 ( 
.A(n_2072),
.B(n_2520),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2145),
.A2(n_2176),
.B(n_2143),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_2192),
.A2(n_2308),
.B(n_2108),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_1981),
.B(n_1988),
.Y(n_3238)
);

A2O1A1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_2537),
.A2(n_2545),
.B(n_2565),
.C(n_2555),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_1952),
.B(n_2654),
.Y(n_3240)
);

CKINVDCx5p33_ASAP7_75t_R g3241 ( 
.A(n_2654),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_1989),
.B(n_1990),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2308),
.A2(n_2974),
.B(n_3070),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_1991),
.B(n_1992),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_1999),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_2759),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_1994),
.B(n_1996),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_1946),
.A2(n_2350),
.B(n_2347),
.Y(n_3248)
);

O2A1O1Ixp33_ASAP7_75t_L g3249 ( 
.A1(n_2537),
.A2(n_2555),
.B(n_2565),
.C(n_2545),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_1997),
.B(n_1998),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2010),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2806),
.B(n_2856),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2408),
.A2(n_2427),
.B(n_2413),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2440),
.A2(n_2493),
.B(n_2450),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2002),
.B(n_2005),
.Y(n_3255)
);

AOI21x1_ASAP7_75t_L g3256 ( 
.A1(n_2326),
.A2(n_2328),
.B(n_2022),
.Y(n_3256)
);

NOR3xp33_ASAP7_75t_L g3257 ( 
.A(n_2570),
.B(n_2593),
.C(n_2584),
.Y(n_3257)
);

AOI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_2503),
.A2(n_2528),
.B(n_2504),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_2529),
.A2(n_2542),
.B(n_2540),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2007),
.B(n_2009),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_2806),
.B(n_2856),
.Y(n_3261)
);

NOR2x1p5_ASAP7_75t_L g3262 ( 
.A(n_2096),
.B(n_2583),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_2141),
.A2(n_2142),
.B(n_2546),
.Y(n_3263)
);

O2A1O1Ixp33_ASAP7_75t_L g3264 ( 
.A1(n_2570),
.A2(n_2593),
.B(n_2605),
.C(n_2584),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2605),
.B(n_2609),
.Y(n_3265)
);

OAI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_2222),
.A2(n_2271),
.B(n_2013),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_2550),
.A2(n_2567),
.B(n_2558),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2012),
.B(n_2018),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_1984),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2024),
.B(n_2025),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_2130),
.B(n_2161),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2026),
.B(n_2027),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2028),
.B(n_2031),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2037),
.B(n_2041),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_2609),
.B(n_2628),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2572),
.A2(n_2639),
.B(n_2602),
.Y(n_3276)
);

NOR3xp33_ASAP7_75t_L g3277 ( 
.A(n_2628),
.B(n_2635),
.C(n_2629),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2034),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2050),
.B(n_2058),
.Y(n_3279)
);

OR2x6_ASAP7_75t_L g3280 ( 
.A(n_2209),
.B(n_2121),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_2739),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_2629),
.B(n_2635),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2651),
.A2(n_2664),
.B(n_2655),
.Y(n_3283)
);

BUFx12f_ASAP7_75t_L g3284 ( 
.A(n_2120),
.Y(n_3284)
);

NAND2x1_ASAP7_75t_L g3285 ( 
.A(n_2206),
.B(n_2322),
.Y(n_3285)
);

CKINVDCx5p33_ASAP7_75t_R g3286 ( 
.A(n_2937),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2063),
.B(n_2066),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2346),
.B(n_2364),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2673),
.A2(n_2686),
.B(n_2679),
.Y(n_3289)
);

A2O1A1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_2653),
.A2(n_2658),
.B(n_2704),
.C(n_2683),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2367),
.B(n_2370),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2687),
.A2(n_2694),
.B(n_2690),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2377),
.B(n_2378),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2386),
.B(n_2387),
.Y(n_3294)
);

AOI22xp33_ASAP7_75t_L g3295 ( 
.A1(n_2653),
.A2(n_2683),
.B1(n_2704),
.B2(n_2658),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_2128),
.Y(n_3296)
);

BUFx6f_ASAP7_75t_L g3297 ( 
.A(n_2739),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2399),
.B(n_2402),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_2094),
.B(n_2239),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2404),
.B(n_2407),
.Y(n_3300)
);

CKINVDCx5p33_ASAP7_75t_R g3301 ( 
.A(n_2937),
.Y(n_3301)
);

BUFx12f_ASAP7_75t_L g3302 ( 
.A(n_2120),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2695),
.A2(n_2710),
.B(n_2699),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_2045),
.B(n_2188),
.Y(n_3304)
);

BUFx4f_ASAP7_75t_L g3305 ( 
.A(n_1947),
.Y(n_3305)
);

NOR2x1_ASAP7_75t_R g3306 ( 
.A(n_2068),
.B(n_2177),
.Y(n_3306)
);

OAI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_2410),
.A2(n_2417),
.B(n_2415),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_2730),
.A2(n_2746),
.B(n_2743),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2751),
.B(n_2781),
.Y(n_3309)
);

BUFx12f_ASAP7_75t_L g3310 ( 
.A(n_2163),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_2751),
.B(n_2781),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_2821),
.B(n_2823),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2821),
.B(n_2823),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2765),
.A2(n_2789),
.B(n_2766),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_2045),
.B(n_2188),
.Y(n_3315)
);

AND2x2_ASAP7_75t_SL g3316 ( 
.A(n_2825),
.B(n_2826),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_2795),
.A2(n_2801),
.B(n_2796),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_2985),
.B(n_2422),
.Y(n_3318)
);

A2O1A1Ixp33_ASAP7_75t_L g3319 ( 
.A1(n_2825),
.A2(n_2897),
.B(n_2898),
.C(n_2826),
.Y(n_3319)
);

O2A1O1Ixp33_ASAP7_75t_L g3320 ( 
.A1(n_2838),
.A2(n_2897),
.B(n_2898),
.C(n_2858),
.Y(n_3320)
);

NOR3xp33_ASAP7_75t_L g3321 ( 
.A(n_2838),
.B(n_2906),
.C(n_2858),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_SL g3322 ( 
.A(n_2985),
.B(n_2423),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2430),
.B(n_2432),
.Y(n_3323)
);

BUFx12f_ASAP7_75t_L g3324 ( 
.A(n_2163),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2434),
.B(n_2436),
.Y(n_3325)
);

OAI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2465),
.A2(n_2469),
.B(n_2468),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2807),
.A2(n_2837),
.B(n_2833),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2889),
.A2(n_2903),
.B(n_2900),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_2906),
.B(n_2910),
.Y(n_3329)
);

NOR2xp67_ASAP7_75t_L g3330 ( 
.A(n_2739),
.B(n_2242),
.Y(n_3330)
);

O2A1O1Ixp33_ASAP7_75t_SL g3331 ( 
.A1(n_3062),
.A2(n_3064),
.B(n_3068),
.C(n_3063),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_2912),
.A2(n_2938),
.B(n_2917),
.Y(n_3332)
);

AOI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_2939),
.A2(n_2949),
.B(n_2947),
.Y(n_3333)
);

OAI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2472),
.A2(n_2482),
.B(n_2477),
.Y(n_3334)
);

BUFx3_ASAP7_75t_L g3335 ( 
.A(n_2128),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2483),
.B(n_2485),
.Y(n_3336)
);

AOI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_2956),
.A2(n_2973),
.B(n_2971),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_2978),
.A2(n_3001),
.B(n_2988),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_2910),
.A2(n_2928),
.B1(n_2932),
.B2(n_2919),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_R g3340 ( 
.A(n_2011),
.B(n_2557),
.Y(n_3340)
);

OR2x2_ASAP7_75t_L g3341 ( 
.A(n_2702),
.B(n_2840),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2494),
.B(n_2495),
.Y(n_3342)
);

AO21x1_ASAP7_75t_L g3343 ( 
.A1(n_2246),
.A2(n_2270),
.B(n_2919),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2928),
.B(n_2932),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_2497),
.B(n_2501),
.Y(n_3345)
);

AND2x6_ASAP7_75t_L g3346 ( 
.A(n_2322),
.B(n_2324),
.Y(n_3346)
);

AOI21x1_ASAP7_75t_L g3347 ( 
.A1(n_2896),
.A2(n_2914),
.B(n_2215),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2049),
.Y(n_3348)
);

O2A1O1Ixp33_ASAP7_75t_L g3349 ( 
.A1(n_2940),
.A2(n_2966),
.B(n_2977),
.C(n_2942),
.Y(n_3349)
);

A2O1A1Ixp33_ASAP7_75t_L g3350 ( 
.A1(n_2940),
.A2(n_2966),
.B(n_2977),
.C(n_2942),
.Y(n_3350)
);

A2O1A1Ixp33_ASAP7_75t_L g3351 ( 
.A1(n_2981),
.A2(n_2986),
.B(n_3019),
.C(n_2982),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2506),
.B(n_2508),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3007),
.A2(n_3025),
.B(n_3024),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2510),
.B(n_2518),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_2981),
.B(n_2982),
.Y(n_3355)
);

AO21x1_ASAP7_75t_L g3356 ( 
.A1(n_2986),
.A2(n_3020),
.B(n_3019),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3032),
.A2(n_3033),
.B(n_2282),
.Y(n_3357)
);

NAND3xp33_ASAP7_75t_L g3358 ( 
.A(n_3020),
.B(n_3054),
.C(n_3038),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_2055),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_2525),
.B(n_2533),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3072),
.A2(n_2535),
.B(n_2534),
.Y(n_3361)
);

NOR3xp33_ASAP7_75t_L g3362 ( 
.A(n_3038),
.B(n_3055),
.C(n_3054),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_1956),
.B(n_2023),
.Y(n_3363)
);

O2A1O1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3055),
.A2(n_2541),
.B(n_2559),
.C(n_2549),
.Y(n_3364)
);

O2A1O1Ixp33_ASAP7_75t_L g3365 ( 
.A1(n_2568),
.A2(n_2581),
.B(n_2590),
.C(n_2588),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_2085),
.B(n_2362),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2081),
.Y(n_3367)
);

AOI21xp33_ASAP7_75t_L g3368 ( 
.A1(n_2155),
.A2(n_2726),
.B(n_2595),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_2754),
.A2(n_2770),
.B(n_2755),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_2067),
.B(n_2077),
.Y(n_3370)
);

INVx4_ASAP7_75t_L g3371 ( 
.A(n_1945),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2596),
.B(n_2616),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_2425),
.B(n_2448),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2622),
.B(n_2623),
.Y(n_3374)
);

OAI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_2627),
.A2(n_2642),
.B(n_2633),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2646),
.B(n_2650),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2656),
.B(n_2659),
.Y(n_3377)
);

O2A1O1Ixp33_ASAP7_75t_L g3378 ( 
.A1(n_2660),
.A2(n_2663),
.B(n_2670),
.C(n_2668),
.Y(n_3378)
);

CKINVDCx20_ASAP7_75t_R g3379 ( 
.A(n_2267),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_2299),
.B(n_2306),
.Y(n_3380)
);

BUFx4f_ASAP7_75t_L g3381 ( 
.A(n_1947),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2698),
.A2(n_2798),
.B(n_2772),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2082),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2674),
.B(n_2685),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2691),
.B(n_2693),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2088),
.Y(n_3386)
);

BUFx3_ASAP7_75t_L g3387 ( 
.A(n_2725),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2089),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_2500),
.B(n_2661),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2775),
.A2(n_2790),
.B(n_2776),
.Y(n_3390)
);

A2O1A1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_2696),
.A2(n_2705),
.B(n_2709),
.C(n_2708),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_L g3392 ( 
.A(n_2711),
.B(n_2718),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_2805),
.A2(n_2899),
.B(n_2846),
.Y(n_3393)
);

AND2x4_ASAP7_75t_L g3394 ( 
.A(n_2315),
.B(n_2317),
.Y(n_3394)
);

AOI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_3060),
.A2(n_2732),
.B(n_2720),
.Y(n_3395)
);

INVx3_ASAP7_75t_L g3396 ( 
.A(n_2321),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2735),
.A2(n_2750),
.B(n_2736),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_2762),
.B(n_2763),
.Y(n_3398)
);

OAI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_2768),
.A2(n_2791),
.B(n_2783),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2792),
.B(n_2810),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_2811),
.B(n_2817),
.Y(n_3401)
);

OR2x2_ASAP7_75t_SL g3402 ( 
.A(n_2822),
.B(n_2835),
.Y(n_3402)
);

AOI21x1_ASAP7_75t_L g3403 ( 
.A1(n_2276),
.A2(n_1949),
.B(n_2338),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_SL g3404 ( 
.A(n_2843),
.B(n_2845),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_2853),
.A2(n_2863),
.B(n_2861),
.Y(n_3405)
);

AOI21xp5_ASAP7_75t_L g3406 ( 
.A1(n_2865),
.A2(n_2870),
.B(n_2868),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2879),
.B(n_2882),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_2886),
.B(n_2888),
.Y(n_3408)
);

NAND2x1p5_ASAP7_75t_L g3409 ( 
.A(n_2475),
.B(n_2496),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2890),
.A2(n_2924),
.B(n_2892),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_2894),
.A2(n_2913),
.B(n_2911),
.Y(n_3411)
);

INVx2_ASAP7_75t_SL g3412 ( 
.A(n_2725),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2923),
.B(n_2927),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_2930),
.A2(n_2945),
.B(n_2944),
.Y(n_3414)
);

AO21x1_ASAP7_75t_L g3415 ( 
.A1(n_2191),
.A2(n_2209),
.B(n_2136),
.Y(n_3415)
);

OAI21x1_ASAP7_75t_L g3416 ( 
.A1(n_2238),
.A2(n_2496),
.B(n_2475),
.Y(n_3416)
);

AOI21x1_ASAP7_75t_L g3417 ( 
.A1(n_2100),
.A2(n_2114),
.B(n_2105),
.Y(n_3417)
);

BUFx12f_ASAP7_75t_L g3418 ( 
.A(n_2539),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2115),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_2759),
.Y(n_3420)
);

A2O1A1Ixp33_ASAP7_75t_L g3421 ( 
.A1(n_2948),
.A2(n_2954),
.B(n_2955),
.C(n_2952),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_2957),
.A2(n_2962),
.B(n_2958),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_2681),
.B(n_2844),
.Y(n_3423)
);

OAI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_2964),
.A2(n_2975),
.B1(n_2980),
.B2(n_2970),
.Y(n_3424)
);

AOI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_2984),
.A2(n_2993),
.B(n_2990),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_SL g3426 ( 
.A(n_2994),
.B(n_2995),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_2997),
.B(n_3002),
.Y(n_3427)
);

AOI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_2155),
.A2(n_3005),
.B1(n_3015),
.B2(n_3003),
.Y(n_3428)
);

AOI21x1_ASAP7_75t_L g3429 ( 
.A1(n_2149),
.A2(n_2166),
.B(n_2159),
.Y(n_3429)
);

OAI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3016),
.A2(n_3026),
.B1(n_3027),
.B2(n_3017),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3034),
.B(n_3036),
.Y(n_3431)
);

BUFx6f_ASAP7_75t_L g3432 ( 
.A(n_1947),
.Y(n_3432)
);

INVxp67_ASAP7_75t_L g3433 ( 
.A(n_2157),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3037),
.B(n_3039),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_2869),
.B(n_2908),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3041),
.B(n_3050),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_2030),
.B(n_2102),
.Y(n_3437)
);

AOI22xp5_ASAP7_75t_L g3438 ( 
.A1(n_2201),
.A2(n_2183),
.B1(n_2169),
.B2(n_2197),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_2030),
.B(n_2909),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_L g3440 ( 
.A1(n_2872),
.A2(n_2893),
.B1(n_2178),
.B2(n_2365),
.Y(n_3440)
);

INVx4_ASAP7_75t_L g3441 ( 
.A(n_1945),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_2243),
.A2(n_2191),
.B(n_2286),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2287),
.B(n_2197),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2268),
.B(n_2170),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_2342),
.A2(n_2379),
.B1(n_2384),
.B2(n_2381),
.Y(n_3445)
);

O2A1O1Ixp33_ASAP7_75t_SL g3446 ( 
.A1(n_2332),
.A2(n_2165),
.B(n_2232),
.C(n_2198),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2268),
.B(n_2187),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_SL g3448 ( 
.A(n_2236),
.B(n_1957),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2182),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2136),
.B(n_1950),
.Y(n_3450)
);

NOR2x1_ASAP7_75t_L g3451 ( 
.A(n_2438),
.B(n_2717),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_2968),
.B(n_3040),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2354),
.B(n_2391),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_2392),
.A2(n_2393),
.B1(n_2401),
.B2(n_2397),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_3061),
.B(n_2086),
.Y(n_3455)
);

OR2x2_ASAP7_75t_L g3456 ( 
.A(n_2087),
.B(n_2091),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2411),
.B(n_2414),
.Y(n_3457)
);

AND2x2_ASAP7_75t_SL g3458 ( 
.A(n_3069),
.B(n_2223),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_2418),
.B(n_2437),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_2416),
.A2(n_2453),
.B1(n_2466),
.B2(n_2435),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_1957),
.B(n_2344),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2441),
.B(n_2446),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2447),
.B(n_2454),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2484),
.B(n_2486),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_2505),
.B(n_2547),
.Y(n_3465)
);

OAI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2223),
.A2(n_2121),
.B(n_2275),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_2093),
.B(n_2344),
.Y(n_3467)
);

AND2x4_ASAP7_75t_L g3468 ( 
.A(n_2594),
.B(n_2600),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_2442),
.B(n_2456),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_2442),
.B(n_2456),
.Y(n_3470)
);

A2O1A1Ixp33_ASAP7_75t_L g3471 ( 
.A1(n_2824),
.A2(n_2278),
.B(n_2205),
.C(n_2244),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_2184),
.A2(n_2186),
.B(n_2185),
.Y(n_3472)
);

AOI21x1_ASAP7_75t_L g3473 ( 
.A1(n_2189),
.A2(n_2199),
.B(n_2195),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2200),
.A2(n_2211),
.B(n_2210),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2553),
.B(n_2562),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2563),
.B(n_2566),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2580),
.B(n_2591),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_2601),
.B(n_2620),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_1947),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2636),
.B(n_2643),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_1966),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_2600),
.A2(n_2741),
.B(n_2607),
.Y(n_3482)
);

AO21x1_ASAP7_75t_L g3483 ( 
.A1(n_2238),
.A2(n_2233),
.B(n_2205),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_1970),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_2470),
.A2(n_2499),
.B1(n_2512),
.B2(n_2490),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_2059),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_1974),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_2059),
.Y(n_3488)
);

OAI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_2280),
.A2(n_2244),
.B(n_2233),
.Y(n_3489)
);

O2A1O1Ixp33_ASAP7_75t_SL g3490 ( 
.A1(n_2340),
.A2(n_2160),
.B(n_2307),
.C(n_2304),
.Y(n_3490)
);

OAI321xp33_ASAP7_75t_L g3491 ( 
.A1(n_2502),
.A2(n_2715),
.A3(n_2573),
.B1(n_2808),
.B2(n_2779),
.C(n_2621),
.Y(n_3491)
);

OAI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_2097),
.A2(n_2573),
.B(n_2502),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_2515),
.A2(n_2526),
.B1(n_2527),
.B2(n_2516),
.Y(n_3493)
);

A2O1A1Ixp33_ASAP7_75t_L g3494 ( 
.A1(n_2260),
.A2(n_2290),
.B(n_2285),
.C(n_2294),
.Y(n_3494)
);

AOI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_2607),
.A2(n_2782),
.B(n_2741),
.Y(n_3495)
);

OAI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_2532),
.A2(n_2544),
.B1(n_2548),
.B2(n_2536),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_2967),
.A2(n_2260),
.B(n_2285),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_1977),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_2000),
.Y(n_3499)
);

A2O1A1Ixp33_ASAP7_75t_L g3500 ( 
.A1(n_2290),
.A2(n_2241),
.B(n_2003),
.C(n_2644),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_2667),
.B(n_2675),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2676),
.B(n_2678),
.Y(n_3502)
);

A2O1A1Ixp33_ASAP7_75t_L g3503 ( 
.A1(n_2680),
.A2(n_2689),
.B(n_2734),
.C(n_2728),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_2004),
.A2(n_2036),
.B(n_2032),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_2043),
.A2(n_2060),
.B(n_2054),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_2062),
.A2(n_2075),
.B(n_2069),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_2076),
.A2(n_2107),
.B(n_2078),
.Y(n_3507)
);

AOI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_2132),
.A2(n_2181),
.B(n_2168),
.Y(n_3508)
);

INVx1_ASAP7_75t_SL g3509 ( 
.A(n_3047),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_2343),
.B(n_2356),
.Y(n_3510)
);

BUFx6f_ASAP7_75t_L g3511 ( 
.A(n_2343),
.Y(n_3511)
);

OAI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_2280),
.A2(n_2258),
.B(n_2255),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_2194),
.A2(n_2212),
.B(n_2207),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_2214),
.A2(n_2219),
.B(n_2218),
.Y(n_3514)
);

OAI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_2582),
.A2(n_2614),
.B1(n_2632),
.B2(n_2598),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2742),
.B(n_2744),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_2745),
.B(n_2749),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_2621),
.B(n_2715),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_2829),
.B(n_2852),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_2059),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_2221),
.A2(n_2229),
.B(n_2225),
.Y(n_3521)
);

OR2x6_ASAP7_75t_L g3522 ( 
.A(n_1971),
.B(n_2006),
.Y(n_3522)
);

BUFx2_ASAP7_75t_L g3523 ( 
.A(n_3053),
.Y(n_3523)
);

OAI21xp33_ASAP7_75t_L g3524 ( 
.A1(n_2097),
.A2(n_2808),
.B(n_2779),
.Y(n_3524)
);

AND2x4_ASAP7_75t_L g3525 ( 
.A(n_2343),
.B(n_2356),
.Y(n_3525)
);

AO21x1_ASAP7_75t_L g3526 ( 
.A1(n_2263),
.A2(n_2288),
.B(n_2234),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_2230),
.A2(n_2247),
.B(n_2235),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_2854),
.B(n_2855),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_2249),
.A2(n_2256),
.B(n_2253),
.Y(n_3529)
);

HB1xp67_ASAP7_75t_L g3530 ( 
.A(n_3053),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2059),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_2867),
.B(n_2918),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2933),
.Y(n_3533)
);

OAI21xp33_ASAP7_75t_L g3534 ( 
.A1(n_2859),
.A2(n_2154),
.B(n_2008),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_2859),
.B(n_2157),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_2259),
.A2(n_2269),
.B(n_2264),
.Y(n_3536)
);

INVxp67_ASAP7_75t_L g3537 ( 
.A(n_3066),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_2169),
.A2(n_2154),
.B1(n_2092),
.B2(n_2359),
.Y(n_3538)
);

HB1xp67_ASAP7_75t_L g3539 ( 
.A(n_3066),
.Y(n_3539)
);

AOI21x1_ASAP7_75t_L g3540 ( 
.A1(n_2273),
.A2(n_2284),
.B(n_2281),
.Y(n_3540)
);

AO21x1_ASAP7_75t_L g3541 ( 
.A1(n_2291),
.A2(n_2293),
.B(n_2647),
.Y(n_3541)
);

CKINVDCx8_ASAP7_75t_R g3542 ( 
.A(n_2177),
.Y(n_3542)
);

AOI21xp5_ASAP7_75t_L g3543 ( 
.A1(n_2946),
.A2(n_3011),
.B(n_2983),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3021),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3031),
.A2(n_3046),
.B(n_3035),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3052),
.B(n_3065),
.Y(n_3546)
);

O2A1O1Ixp33_ASAP7_75t_L g3547 ( 
.A1(n_2193),
.A2(n_1971),
.B(n_2173),
.C(n_2213),
.Y(n_3547)
);

BUFx4f_ASAP7_75t_L g3548 ( 
.A(n_2343),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_2135),
.B(n_2119),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_1945),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_2356),
.A2(n_2464),
.B(n_2373),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_2356),
.A2(n_2464),
.B(n_2373),
.Y(n_3552)
);

NAND2x1p5_ASAP7_75t_L g3553 ( 
.A(n_2373),
.B(n_2464),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_1945),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_2298),
.A2(n_2682),
.B(n_2737),
.C(n_2697),
.Y(n_3555)
);

INVx2_ASAP7_75t_SL g3556 ( 
.A(n_2725),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_SL g3557 ( 
.A(n_2382),
.B(n_2421),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_2172),
.B(n_2193),
.Y(n_3558)
);

O2A1O1Ixp33_ASAP7_75t_SL g3559 ( 
.A1(n_2738),
.A2(n_2740),
.B(n_2778),
.C(n_2753),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_2373),
.A2(n_2492),
.B(n_2464),
.Y(n_3560)
);

O2A1O1Ixp33_ASAP7_75t_SL g3561 ( 
.A1(n_2785),
.A2(n_2800),
.B(n_2813),
.C(n_2802),
.Y(n_3561)
);

O2A1O1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_2173),
.A2(n_2046),
.B(n_2138),
.C(n_2104),
.Y(n_3562)
);

BUFx6f_ASAP7_75t_L g3563 ( 
.A(n_2492),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_2492),
.A2(n_2637),
.B(n_2523),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2492),
.A2(n_2637),
.B(n_2523),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_2523),
.A2(n_2657),
.B(n_2637),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_1993),
.B(n_1987),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_2523),
.A2(n_2657),
.B(n_2637),
.Y(n_3568)
);

AOI21x1_ASAP7_75t_L g3569 ( 
.A1(n_2217),
.A2(n_2227),
.B(n_2224),
.Y(n_3569)
);

O2A1O1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_2046),
.A2(n_2104),
.B(n_2138),
.C(n_1987),
.Y(n_3570)
);

BUFx6f_ASAP7_75t_L g3571 ( 
.A(n_2657),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_1945),
.Y(n_3572)
);

AND2x4_ASAP7_75t_L g3573 ( 
.A(n_2657),
.B(n_2713),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_2713),
.A2(n_2883),
.B(n_2296),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2713),
.A2(n_2883),
.B(n_2819),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_2713),
.A2(n_2883),
.B(n_2820),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2816),
.B(n_2828),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_2830),
.B(n_2839),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_2571),
.B(n_2577),
.Y(n_3579)
);

OR2x2_ASAP7_75t_L g3580 ( 
.A(n_2841),
.B(n_2842),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_2883),
.A2(n_2849),
.B(n_2847),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_2298),
.A2(n_2887),
.B(n_2905),
.C(n_2874),
.Y(n_3582)
);

NOR3xp33_ASAP7_75t_L g3583 ( 
.A(n_2240),
.B(n_2250),
.C(n_2248),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_2920),
.B(n_2925),
.Y(n_3584)
);

AOI33xp33_ASAP7_75t_L g3585 ( 
.A1(n_2929),
.A2(n_3073),
.A3(n_2931),
.B1(n_2934),
.B2(n_2936),
.B3(n_2943),
.Y(n_3585)
);

BUFx6f_ASAP7_75t_L g3586 ( 
.A(n_2424),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_2951),
.B(n_2959),
.Y(n_3587)
);

OR2x2_ASAP7_75t_SL g3588 ( 
.A(n_2266),
.B(n_2228),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_2960),
.B(n_2963),
.Y(n_3589)
);

NAND2x1p5_ASAP7_75t_L g3590 ( 
.A(n_2571),
.B(n_2577),
.Y(n_3590)
);

NOR2xp33_ASAP7_75t_L g3591 ( 
.A(n_2295),
.B(n_2289),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2424),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_2965),
.A2(n_2987),
.B(n_2979),
.Y(n_3593)
);

NAND2xp33_ASAP7_75t_L g3594 ( 
.A(n_2476),
.B(n_2521),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_2989),
.B(n_2991),
.Y(n_3595)
);

OR2x2_ASAP7_75t_L g3596 ( 
.A(n_3000),
.B(n_3006),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_2597),
.B(n_2603),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3010),
.B(n_3012),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3014),
.B(n_3022),
.Y(n_3599)
);

O2A1O1Ixp5_ASAP7_75t_L g3600 ( 
.A1(n_2336),
.A2(n_2339),
.B(n_3028),
.C(n_3029),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_2001),
.A2(n_2420),
.B(n_2403),
.Y(n_3601)
);

INVxp67_ASAP7_75t_L g3602 ( 
.A(n_2216),
.Y(n_3602)
);

AOI22xp5_ASAP7_75t_L g3603 ( 
.A1(n_2597),
.A2(n_2672),
.B1(n_2603),
.B2(n_2707),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_2065),
.B(n_2757),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_2424),
.Y(n_3605)
);

OAI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_2001),
.A2(n_2190),
.B1(n_2618),
.B2(n_2420),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_2424),
.B(n_2611),
.Y(n_3607)
);

O2A1O1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_2272),
.A2(n_2309),
.B(n_2316),
.C(n_2312),
.Y(n_3608)
);

INVxp67_ASAP7_75t_SL g3609 ( 
.A(n_2279),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_2424),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_L g3611 ( 
.A(n_2065),
.B(n_2761),
.Y(n_3611)
);

NOR3xp33_ASAP7_75t_L g3612 ( 
.A(n_2297),
.B(n_2707),
.C(n_2672),
.Y(n_3612)
);

O2A1O1Ixp5_ASAP7_75t_L g3613 ( 
.A1(n_2314),
.A2(n_2329),
.B(n_2331),
.C(n_3018),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_2611),
.Y(n_3614)
);

OAI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_2611),
.A2(n_2831),
.B(n_2617),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_2611),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2403),
.A2(n_2618),
.B(n_2420),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2403),
.A2(n_2648),
.B(n_2618),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_2976),
.B(n_3018),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_2611),
.B(n_2831),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_2831),
.Y(n_3621)
);

BUFx12f_ASAP7_75t_L g3622 ( 
.A(n_2539),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2648),
.A2(n_2716),
.B(n_2649),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_2831),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_2831),
.B(n_2976),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_2587),
.B(n_2617),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_2587),
.A2(n_2665),
.B(n_2662),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_R g3628 ( 
.A(n_2786),
.B(n_2827),
.Y(n_3628)
);

HB1xp67_ASAP7_75t_L g3629 ( 
.A(n_2216),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_2907),
.B(n_2301),
.Y(n_3630)
);

AND2x6_ASAP7_75t_SL g3631 ( 
.A(n_2330),
.B(n_2006),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_2177),
.B(n_2292),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_2662),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_2665),
.B(n_2857),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_2857),
.B(n_2648),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_2245),
.B(n_2251),
.Y(n_3636)
);

AOI21x1_ASAP7_75t_L g3637 ( 
.A1(n_2302),
.A2(n_2251),
.B(n_2325),
.Y(n_3637)
);

INVx5_ASAP7_75t_L g3638 ( 
.A(n_2090),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_2303),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_2649),
.A2(n_2812),
.B(n_2723),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_2649),
.B(n_2716),
.Y(n_3641)
);

AND2x2_ASAP7_75t_SL g3642 ( 
.A(n_2064),
.B(n_2327),
.Y(n_3642)
);

NOR2xp33_ASAP7_75t_L g3643 ( 
.A(n_2323),
.B(n_2064),
.Y(n_3643)
);

HB1xp67_ASAP7_75t_L g3644 ( 
.A(n_2716),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_1948),
.Y(n_3645)
);

INVx3_ASAP7_75t_L g3646 ( 
.A(n_2098),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_2723),
.B(n_2812),
.Y(n_3647)
);

OAI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_2723),
.A2(n_2812),
.B1(n_2006),
.B2(n_1965),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_1948),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_2864),
.B(n_2881),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2864),
.B(n_2881),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_SL g3652 ( 
.A(n_2017),
.B(n_2125),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_1948),
.Y(n_3653)
);

AO21x2_ASAP7_75t_L g3654 ( 
.A1(n_2319),
.A2(n_2335),
.B(n_2333),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_2177),
.B(n_2133),
.Y(n_3655)
);

OR2x2_ASAP7_75t_L g3656 ( 
.A(n_1951),
.B(n_1986),
.Y(n_3656)
);

AOI21x1_ASAP7_75t_L g3657 ( 
.A1(n_2196),
.A2(n_2204),
.B(n_2330),
.Y(n_3657)
);

AOI21x1_ASAP7_75t_L g3658 ( 
.A1(n_2196),
.A2(n_2204),
.B(n_2330),
.Y(n_3658)
);

OAI21xp33_ASAP7_75t_L g3659 ( 
.A1(n_2329),
.A2(n_2331),
.B(n_2543),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_2864),
.B(n_2881),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_2901),
.B(n_1967),
.Y(n_3661)
);

OAI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_2320),
.A2(n_2196),
.B(n_2204),
.Y(n_3662)
);

AOI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_2901),
.A2(n_2452),
.B(n_3051),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_2901),
.B(n_1967),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2428),
.B(n_2479),
.Y(n_3665)
);

OAI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_2320),
.A2(n_2380),
.B(n_2700),
.Y(n_3666)
);

A2O1A1Ixp33_ASAP7_75t_L g3667 ( 
.A1(n_2524),
.A2(n_2671),
.B(n_2788),
.C(n_2556),
.Y(n_3667)
);

AOI22xp33_ASAP7_75t_L g3668 ( 
.A1(n_2017),
.A2(n_2334),
.B1(n_2220),
.B2(n_2488),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_2048),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_2428),
.B(n_2479),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_1948),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_2514),
.B(n_2585),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_2560),
.A2(n_2610),
.B(n_2652),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_2020),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_2020),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2514),
.B(n_2585),
.Y(n_3676)
);

INVx3_ASAP7_75t_L g3677 ( 
.A(n_2020),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_2429),
.B(n_2631),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_2589),
.B(n_3071),
.Y(n_3679)
);

OAI21xp33_ASAP7_75t_L g3680 ( 
.A1(n_2809),
.A2(n_2016),
.B(n_2021),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_2701),
.A2(n_2902),
.B(n_3008),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_2589),
.B(n_3071),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_2020),
.Y(n_3683)
);

CKINVDCx8_ASAP7_75t_R g3684 ( 
.A(n_2363),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_2274),
.Y(n_3685)
);

OAI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_2310),
.A2(n_3057),
.B(n_2619),
.Y(n_3686)
);

AND2x4_ASAP7_75t_SL g3687 ( 
.A(n_2619),
.B(n_3057),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_2666),
.A2(n_2873),
.B(n_2669),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_2666),
.A2(n_2873),
.B(n_2669),
.Y(n_3689)
);

NOR2xp67_ASAP7_75t_L g3690 ( 
.A(n_2277),
.B(n_2261),
.Y(n_3690)
);

INVx3_ASAP7_75t_L g3691 ( 
.A(n_2274),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_2017),
.A2(n_2429),
.B(n_2631),
.Y(n_3692)
);

OAI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_2257),
.A2(n_2038),
.B(n_2056),
.Y(n_3693)
);

CKINVDCx10_ASAP7_75t_R g3694 ( 
.A(n_2252),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_2274),
.B(n_2283),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_2274),
.A2(n_2283),
.B(n_3056),
.Y(n_3696)
);

AND2x4_ASAP7_75t_L g3697 ( 
.A(n_2150),
.B(n_2357),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_2722),
.B(n_2972),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_2283),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_2283),
.B(n_2773),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_2794),
.B(n_2797),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_2862),
.B(n_2999),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_2146),
.B(n_2254),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_2252),
.B(n_2265),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_2405),
.A2(n_3049),
.B(n_2771),
.Y(n_3705)
);

NAND2x1_ASAP7_75t_L g3706 ( 
.A(n_2265),
.B(n_2261),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_2267),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_2478),
.A2(n_2552),
.B(n_2769),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_2305),
.Y(n_3709)
);

BUFx2_ASAP7_75t_L g3710 ( 
.A(n_2592),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_2727),
.B(n_2265),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_2146),
.Y(n_3712)
);

AO21x2_ASAP7_75t_L g3713 ( 
.A1(n_2337),
.A2(n_2625),
.B(n_2406),
.Y(n_3713)
);

A2O1A1Ixp33_ASAP7_75t_L g3714 ( 
.A1(n_2144),
.A2(n_2226),
.B(n_2180),
.C(n_2147),
.Y(n_3714)
);

OAI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_2916),
.A2(n_2116),
.B1(n_2208),
.B2(n_2254),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_2144),
.A2(n_2226),
.B(n_2164),
.Y(n_3716)
);

OR2x6_ASAP7_75t_L g3717 ( 
.A(n_2144),
.B(n_2226),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_2231),
.B(n_2139),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_2179),
.B(n_1968),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3720)
);

AOI22xp5_ASAP7_75t_L g3721 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3722)
);

INVx4_ASAP7_75t_L g3723 ( 
.A(n_2035),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_2311),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3727)
);

A2O1A1Ixp33_ASAP7_75t_L g3728 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3728)
);

O2A1O1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_2311),
.Y(n_3731)
);

HB1xp67_ASAP7_75t_L g3732 ( 
.A(n_2431),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_2074),
.B(n_2052),
.Y(n_3733)
);

OR2x2_ASAP7_75t_L g3734 ( 
.A(n_1983),
.B(n_1959),
.Y(n_3734)
);

BUFx8_ASAP7_75t_SL g3735 ( 
.A(n_2345),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3736)
);

NOR2x2_ASAP7_75t_L g3737 ( 
.A(n_2252),
.B(n_2265),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_2311),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_2431),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_2311),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3745)
);

O2A1O1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3746)
);

A2O1A1Ixp33_ASAP7_75t_L g3747 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_2311),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_2311),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_L g3750 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3750)
);

NOR2xp33_ASAP7_75t_L g3751 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3751)
);

O2A1O1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3752)
);

BUFx3_ASAP7_75t_L g3753 ( 
.A(n_2128),
.Y(n_3753)
);

BUFx6f_ASAP7_75t_L g3754 ( 
.A(n_2300),
.Y(n_3754)
);

NAND3xp33_ASAP7_75t_L g3755 ( 
.A(n_2578),
.B(n_1051),
.C(n_1213),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3756)
);

NAND2xp33_ASAP7_75t_L g3757 ( 
.A(n_2578),
.B(n_2748),
.Y(n_3757)
);

AO21x1_ASAP7_75t_L g3758 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3759)
);

AOI21x1_ASAP7_75t_L g3760 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_2311),
.Y(n_3761)
);

AO21x1_ASAP7_75t_L g3762 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3764)
);

NOR2xp33_ASAP7_75t_R g3765 ( 
.A(n_2011),
.B(n_1030),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_2311),
.Y(n_3767)
);

NOR2xp33_ASAP7_75t_L g3768 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3770)
);

BUFx6f_ASAP7_75t_L g3771 ( 
.A(n_2300),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3772)
);

OR2x6_ASAP7_75t_L g3773 ( 
.A(n_2084),
.B(n_2158),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3780)
);

O2A1O1Ixp33_ASAP7_75t_SL g3781 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3782)
);

AO21x1_ASAP7_75t_L g3783 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3786)
);

OAI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3789)
);

INVx2_ASAP7_75t_SL g3790 ( 
.A(n_1984),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3791)
);

AOI22xp33_ASAP7_75t_L g3792 ( 
.A1(n_1968),
.A2(n_2371),
.B1(n_2375),
.B2(n_2366),
.Y(n_3792)
);

AOI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3795)
);

BUFx8_ASAP7_75t_L g3796 ( 
.A(n_1965),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_L g3797 ( 
.A(n_2300),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3798)
);

INVx2_ASAP7_75t_SL g3799 ( 
.A(n_1984),
.Y(n_3799)
);

CKINVDCx20_ASAP7_75t_R g3800 ( 
.A(n_2011),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3801)
);

AOI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3804)
);

O2A1O1Ixp33_ASAP7_75t_L g3805 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3805)
);

AOI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_2128),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3808)
);

AOI21x1_ASAP7_75t_L g3809 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3810)
);

AO21x1_ASAP7_75t_L g3811 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3811)
);

AOI21x1_ASAP7_75t_L g3812 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3812)
);

OAI22xp5_ASAP7_75t_L g3813 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_SL g3814 ( 
.A(n_2561),
.B(n_2626),
.Y(n_3814)
);

OAI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3815)
);

AO21x1_ASAP7_75t_L g3816 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_2311),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3820)
);

O2A1O1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_L g3823 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_2311),
.Y(n_3830)
);

INVxp67_ASAP7_75t_L g3831 ( 
.A(n_2157),
.Y(n_3831)
);

AOI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3832)
);

BUFx6f_ASAP7_75t_L g3833 ( 
.A(n_2300),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_2074),
.B(n_2052),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3837)
);

NOR2xp33_ASAP7_75t_SL g3838 ( 
.A(n_2561),
.B(n_2626),
.Y(n_3838)
);

AOI21xp5_ASAP7_75t_L g3839 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3842)
);

AOI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3846)
);

OAI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3849)
);

A2O1A1Ixp33_ASAP7_75t_L g3850 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3851)
);

AND2x4_ASAP7_75t_L g3852 ( 
.A(n_2074),
.B(n_2052),
.Y(n_3852)
);

NOR2xp67_ASAP7_75t_L g3853 ( 
.A(n_2095),
.B(n_2035),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3854)
);

AOI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3855)
);

A2O1A1Ixp33_ASAP7_75t_L g3856 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_L g3857 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3857)
);

O2A1O1Ixp33_ASAP7_75t_SL g3858 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3858)
);

OAI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3859)
);

AOI21xp5_ASAP7_75t_L g3860 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3863)
);

NOR2xp33_ASAP7_75t_L g3864 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3864)
);

INVx4_ASAP7_75t_L g3865 ( 
.A(n_2035),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_2311),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_2311),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3869)
);

A2O1A1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_2311),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3876)
);

OAI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_2311),
.Y(n_3881)
);

O2A1O1Ixp33_ASAP7_75t_L g3882 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_SL g3883 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3883)
);

CKINVDCx5p33_ASAP7_75t_R g3884 ( 
.A(n_2654),
.Y(n_3884)
);

O2A1O1Ixp5_ASAP7_75t_L g3885 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3887)
);

BUFx2_ASAP7_75t_L g3888 ( 
.A(n_2431),
.Y(n_3888)
);

O2A1O1Ixp33_ASAP7_75t_SL g3889 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_SL g3890 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_L g3893 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3893)
);

AOI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3897)
);

O2A1O1Ixp33_ASAP7_75t_L g3898 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3899)
);

INVx2_ASAP7_75t_SL g3900 ( 
.A(n_1984),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_2311),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3903)
);

CKINVDCx8_ASAP7_75t_R g3904 ( 
.A(n_2177),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_SL g3906 ( 
.A(n_2561),
.B(n_2626),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3909)
);

NOR2xp33_ASAP7_75t_L g3910 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3913)
);

OAI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3915)
);

BUFx6f_ASAP7_75t_L g3916 ( 
.A(n_2300),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_2311),
.Y(n_3919)
);

OAI21xp33_ASAP7_75t_L g3920 ( 
.A1(n_2341),
.A2(n_1109),
.B(n_1013),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_2311),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_2311),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3925)
);

BUFx12f_ASAP7_75t_L g3926 ( 
.A(n_2040),
.Y(n_3926)
);

O2A1O1Ixp33_ASAP7_75t_L g3927 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_3927)
);

NOR2xp33_ASAP7_75t_L g3928 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3928)
);

OAI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3929)
);

AOI21x1_ASAP7_75t_L g3930 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3931)
);

O2A1O1Ixp5_ASAP7_75t_L g3932 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3932)
);

OAI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_2311),
.Y(n_3938)
);

OAI21x1_ASAP7_75t_L g3939 ( 
.A1(n_2574),
.A2(n_2158),
.B(n_2203),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3941)
);

OAI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3943)
);

A2O1A1Ixp33_ASAP7_75t_L g3944 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3946)
);

AOI21x1_ASAP7_75t_L g3947 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3947)
);

NAND2x1_ASAP7_75t_L g3948 ( 
.A(n_2073),
.B(n_2099),
.Y(n_3948)
);

BUFx4f_ASAP7_75t_L g3949 ( 
.A(n_1947),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3952)
);

A2O1A1Ixp33_ASAP7_75t_L g3953 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3953)
);

AOI21xp33_ASAP7_75t_L g3954 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3955)
);

AOI21x1_ASAP7_75t_L g3956 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3957)
);

INVx4_ASAP7_75t_L g3958 ( 
.A(n_2035),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3959)
);

INVxp67_ASAP7_75t_L g3960 ( 
.A(n_2157),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_2311),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3965)
);

AO21x1_ASAP7_75t_L g3966 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_2804),
.B(n_2578),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3972)
);

HB1xp67_ASAP7_75t_L g3973 ( 
.A(n_2431),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3974)
);

INVx4_ASAP7_75t_L g3975 ( 
.A(n_2035),
.Y(n_3975)
);

AO21x2_ASAP7_75t_L g3976 ( 
.A1(n_2158),
.A2(n_2366),
.B(n_1968),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_2311),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3978)
);

INVx2_ASAP7_75t_SL g3979 ( 
.A(n_1984),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_2311),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_2311),
.Y(n_3981)
);

INVx5_ASAP7_75t_L g3982 ( 
.A(n_2035),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3983)
);

AOI21x1_ASAP7_75t_L g3984 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_3984)
);

O2A1O1Ixp5_ASAP7_75t_L g3985 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_2311),
.Y(n_3986)
);

O2A1O1Ixp5_ASAP7_75t_L g3987 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_2074),
.B(n_2052),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_1973),
.B(n_1958),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_2351),
.B(n_2624),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_3993)
);

A2O1A1Ixp33_ASAP7_75t_L g3994 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3995)
);

AO21x1_ASAP7_75t_L g3996 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3996)
);

OAI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_3997)
);

NOR3xp33_ASAP7_75t_L g3998 ( 
.A(n_2834),
.B(n_1119),
.C(n_1090),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_1968),
.B(n_2366),
.Y(n_3999)
);

HB1xp67_ASAP7_75t_L g4000 ( 
.A(n_2431),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_2311),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4003)
);

NAND2x1p5_ASAP7_75t_L g4004 ( 
.A(n_2035),
.B(n_2419),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4006)
);

OAI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4007)
);

O2A1O1Ixp33_ASAP7_75t_SL g4008 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_4008)
);

INVx4_ASAP7_75t_L g4009 ( 
.A(n_2035),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_2311),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_2311),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4016)
);

O2A1O1Ixp5_ASAP7_75t_L g4017 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4019)
);

INVxp67_ASAP7_75t_L g4020 ( 
.A(n_2157),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4026)
);

AO21x1_ASAP7_75t_L g4027 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_2311),
.Y(n_4028)
);

AOI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4030)
);

BUFx8_ASAP7_75t_SL g4031 ( 
.A(n_2345),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4034)
);

BUFx12f_ASAP7_75t_L g4035 ( 
.A(n_2040),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4036)
);

HB1xp67_ASAP7_75t_L g4037 ( 
.A(n_2431),
.Y(n_4037)
);

BUFx2_ASAP7_75t_SL g4038 ( 
.A(n_2035),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4039)
);

AOI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_SL g4043 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_2311),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4045)
);

INVx4_ASAP7_75t_L g4046 ( 
.A(n_2035),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_2311),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4050)
);

OAI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4051)
);

O2A1O1Ixp5_ASAP7_75t_L g4052 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_4052)
);

BUFx6f_ASAP7_75t_L g4053 ( 
.A(n_2300),
.Y(n_4053)
);

AOI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4054)
);

OAI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4055)
);

INVxp67_ASAP7_75t_L g4056 ( 
.A(n_2157),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4057)
);

INVx1_ASAP7_75t_SL g4058 ( 
.A(n_2109),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_2311),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_2311),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_2311),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4067)
);

O2A1O1Ixp5_ASAP7_75t_L g4068 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4069)
);

A2O1A1Ixp33_ASAP7_75t_L g4070 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4070)
);

AND2x4_ASAP7_75t_L g4071 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4071)
);

OAI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_2311),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4076)
);

O2A1O1Ixp33_ASAP7_75t_L g4077 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4079)
);

INVx1_ASAP7_75t_SL g4080 ( 
.A(n_2109),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_2311),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_2431),
.Y(n_4082)
);

OAI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4085)
);

OAI21xp5_ASAP7_75t_L g4086 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4087)
);

OAI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4089)
);

A2O1A1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4092)
);

OAI21x1_ASAP7_75t_L g4093 ( 
.A1(n_2574),
.A2(n_2158),
.B(n_2203),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_2431),
.Y(n_4094)
);

AOI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_L g4098 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4098)
);

BUFx2_ASAP7_75t_L g4099 ( 
.A(n_2431),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4100)
);

AOI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4101)
);

INVx4_ASAP7_75t_L g4102 ( 
.A(n_2035),
.Y(n_4102)
);

BUFx2_ASAP7_75t_L g4103 ( 
.A(n_2431),
.Y(n_4103)
);

INVx4_ASAP7_75t_L g4104 ( 
.A(n_2035),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_2311),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_SL g4106 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4107)
);

BUFx2_ASAP7_75t_SL g4108 ( 
.A(n_2035),
.Y(n_4108)
);

A2O1A1Ixp33_ASAP7_75t_L g4109 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4110)
);

AOI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_2311),
.Y(n_4112)
);

OAI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4113)
);

BUFx4f_ASAP7_75t_L g4114 ( 
.A(n_1947),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4115)
);

OAI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_L g4117 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4118)
);

INVx3_ASAP7_75t_L g4119 ( 
.A(n_2052),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4120)
);

INVx3_ASAP7_75t_L g4121 ( 
.A(n_2052),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4122)
);

AOI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4124)
);

AOI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4125)
);

INVx3_ASAP7_75t_L g4126 ( 
.A(n_2052),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4127)
);

OAI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_2311),
.Y(n_4129)
);

INVxp67_ASAP7_75t_L g4130 ( 
.A(n_2157),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4133)
);

AO21x1_ASAP7_75t_L g4134 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_2311),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4141)
);

AOI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4142)
);

NOR2x1_ASAP7_75t_L g4143 ( 
.A(n_2101),
.B(n_2123),
.Y(n_4143)
);

OAI21xp5_ASAP7_75t_L g4144 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4144)
);

NOR2xp67_ASAP7_75t_L g4145 ( 
.A(n_2095),
.B(n_2035),
.Y(n_4145)
);

AOI21xp33_ASAP7_75t_L g4146 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4148)
);

NOR2x1_ASAP7_75t_L g4149 ( 
.A(n_2101),
.B(n_2123),
.Y(n_4149)
);

OAI22xp5_ASAP7_75t_L g4150 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_L g4152 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_2311),
.Y(n_4153)
);

INVx4_ASAP7_75t_L g4154 ( 
.A(n_2035),
.Y(n_4154)
);

O2A1O1Ixp33_ASAP7_75t_L g4155 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4156)
);

OAI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4157)
);

OAI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4161)
);

INVx4_ASAP7_75t_L g4162 ( 
.A(n_2035),
.Y(n_4162)
);

NOR2xp33_ASAP7_75t_L g4163 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4163)
);

AOI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4166)
);

O2A1O1Ixp33_ASAP7_75t_L g4167 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4169)
);

AOI21xp5_ASAP7_75t_L g4170 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4170)
);

O2A1O1Ixp33_ASAP7_75t_L g4171 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4171)
);

OAI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4174)
);

INVx3_ASAP7_75t_L g4175 ( 
.A(n_2052),
.Y(n_4175)
);

CKINVDCx5p33_ASAP7_75t_R g4176 ( 
.A(n_2654),
.Y(n_4176)
);

OAI21x1_ASAP7_75t_L g4177 ( 
.A1(n_2574),
.A2(n_2158),
.B(n_2203),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_2311),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4179)
);

A2O1A1Ixp33_ASAP7_75t_L g4180 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4180)
);

BUFx6f_ASAP7_75t_L g4181 ( 
.A(n_2300),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4183)
);

NOR2xp33_ASAP7_75t_L g4184 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4184)
);

AOI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4187)
);

AOI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4188)
);

OAI21xp33_ASAP7_75t_L g4189 ( 
.A1(n_2341),
.A2(n_1109),
.B(n_1013),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4190)
);

NAND3xp33_ASAP7_75t_L g4191 ( 
.A(n_2578),
.B(n_1051),
.C(n_1213),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4192)
);

INVx4_ASAP7_75t_L g4193 ( 
.A(n_2035),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4194)
);

A2O1A1Ixp33_ASAP7_75t_L g4195 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4195)
);

OAI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4197)
);

AOI21xp5_ASAP7_75t_L g4198 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4198)
);

OAI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_SL g4202 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4203)
);

BUFx2_ASAP7_75t_L g4204 ( 
.A(n_2431),
.Y(n_4204)
);

NOR2xp33_ASAP7_75t_R g4205 ( 
.A(n_2011),
.B(n_1030),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4206)
);

NOR2xp33_ASAP7_75t_L g4207 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4207)
);

AOI21xp5_ASAP7_75t_L g4208 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4208)
);

INVx2_ASAP7_75t_SL g4209 ( 
.A(n_1984),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4210)
);

AOI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4211)
);

BUFx6f_ASAP7_75t_L g4212 ( 
.A(n_2300),
.Y(n_4212)
);

BUFx2_ASAP7_75t_L g4213 ( 
.A(n_2431),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4218)
);

AOI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_2311),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4223)
);

OAI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_1983),
.B(n_1959),
.Y(n_4227)
);

BUFx6f_ASAP7_75t_L g4228 ( 
.A(n_2300),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4229)
);

AOI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_2654),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4235)
);

HB1xp67_ASAP7_75t_L g4236 ( 
.A(n_2431),
.Y(n_4236)
);

O2A1O1Ixp33_ASAP7_75t_L g4237 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4239)
);

NOR3xp33_ASAP7_75t_L g4240 ( 
.A(n_2834),
.B(n_1119),
.C(n_1090),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_2311),
.Y(n_4241)
);

OR2x2_ASAP7_75t_L g4242 ( 
.A(n_1983),
.B(n_1959),
.Y(n_4242)
);

BUFx2_ASAP7_75t_L g4243 ( 
.A(n_2431),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4247)
);

INVx2_ASAP7_75t_SL g4248 ( 
.A(n_1984),
.Y(n_4248)
);

INVx3_ASAP7_75t_L g4249 ( 
.A(n_2052),
.Y(n_4249)
);

INVx3_ASAP7_75t_L g4250 ( 
.A(n_2052),
.Y(n_4250)
);

OAI321xp33_ASAP7_75t_L g4251 ( 
.A1(n_1968),
.A2(n_1090),
.A3(n_1119),
.B1(n_2366),
.B2(n_2375),
.C(n_2371),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4252)
);

AO21x1_ASAP7_75t_L g4253 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4253)
);

AOI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4255)
);

BUFx2_ASAP7_75t_L g4256 ( 
.A(n_2431),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4257)
);

OAI21xp33_ASAP7_75t_L g4258 ( 
.A1(n_2341),
.A2(n_1109),
.B(n_1013),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_2157),
.Y(n_4259)
);

OR2x6_ASAP7_75t_L g4260 ( 
.A(n_2084),
.B(n_2158),
.Y(n_4260)
);

AOI21xp5_ASAP7_75t_L g4261 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_2311),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4265)
);

AOI21x1_ASAP7_75t_L g4266 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_4266)
);

BUFx6f_ASAP7_75t_L g4267 ( 
.A(n_2300),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4268)
);

AOI21xp5_ASAP7_75t_L g4269 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4269)
);

OR2x6_ASAP7_75t_SL g4270 ( 
.A(n_2461),
.B(n_2531),
.Y(n_4270)
);

AND2x4_ASAP7_75t_L g4271 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_2300),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4274)
);

A2O1A1Ixp33_ASAP7_75t_L g4275 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4276)
);

CKINVDCx5p33_ASAP7_75t_R g4277 ( 
.A(n_2654),
.Y(n_4277)
);

AO22x1_ASAP7_75t_L g4278 ( 
.A1(n_2578),
.A2(n_1013),
.B1(n_1148),
.B2(n_1109),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_2311),
.Y(n_4279)
);

A2O1A1Ixp33_ASAP7_75t_L g4280 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_SL g4281 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4281)
);

BUFx4f_ASAP7_75t_L g4282 ( 
.A(n_1947),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4283)
);

AOI33xp33_ASAP7_75t_L g4284 ( 
.A1(n_2351),
.A2(n_1051),
.A3(n_1099),
.B1(n_1164),
.B2(n_1093),
.B3(n_1713),
.Y(n_4284)
);

BUFx6f_ASAP7_75t_L g4285 ( 
.A(n_2300),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_2311),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_SL g4287 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4287)
);

NOR2x1_ASAP7_75t_L g4288 ( 
.A(n_2101),
.B(n_2123),
.Y(n_4288)
);

OAI22xp5_ASAP7_75t_L g4289 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4289)
);

OAI21xp5_ASAP7_75t_L g4290 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4291)
);

AOI22xp33_ASAP7_75t_L g4292 ( 
.A1(n_1968),
.A2(n_2371),
.B1(n_2375),
.B2(n_2366),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4293)
);

HB1xp67_ASAP7_75t_L g4294 ( 
.A(n_2431),
.Y(n_4294)
);

INVx3_ASAP7_75t_L g4295 ( 
.A(n_2052),
.Y(n_4295)
);

OAI21xp33_ASAP7_75t_L g4296 ( 
.A1(n_2341),
.A2(n_1109),
.B(n_1013),
.Y(n_4296)
);

AOI22xp5_ASAP7_75t_L g4297 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_1983),
.B(n_1959),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_2311),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_L g4301 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4301)
);

HB1xp67_ASAP7_75t_L g4302 ( 
.A(n_2431),
.Y(n_4302)
);

A2O1A1Ixp33_ASAP7_75t_L g4303 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4303)
);

AOI22xp5_ASAP7_75t_L g4304 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4306)
);

AOI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4310)
);

AOI21xp5_ASAP7_75t_L g4311 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4312)
);

A2O1A1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4313)
);

NOR2xp33_ASAP7_75t_L g4314 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4314)
);

O2A1O1Ixp33_ASAP7_75t_SL g4315 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2375),
.C(n_2366),
.Y(n_4315)
);

INVx11_ASAP7_75t_L g4316 ( 
.A(n_2120),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4318)
);

NOR3xp33_ASAP7_75t_L g4319 ( 
.A(n_2834),
.B(n_1119),
.C(n_1090),
.Y(n_4319)
);

BUFx3_ASAP7_75t_L g4320 ( 
.A(n_2128),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4321)
);

AOI22xp33_ASAP7_75t_L g4322 ( 
.A1(n_1968),
.A2(n_2371),
.B1(n_2375),
.B2(n_2366),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4323)
);

OAI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_SL g4325 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_2804),
.B(n_2578),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4328)
);

OAI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4331)
);

OR2x6_ASAP7_75t_L g4332 ( 
.A(n_2084),
.B(n_2158),
.Y(n_4332)
);

NOR3xp33_ASAP7_75t_L g4333 ( 
.A(n_2834),
.B(n_1119),
.C(n_1090),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4334)
);

AOI21x1_ASAP7_75t_L g4335 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_4335)
);

AOI21xp5_ASAP7_75t_L g4336 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4336)
);

AND2x2_ASAP7_75t_SL g4337 ( 
.A(n_2551),
.B(n_2818),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_2311),
.Y(n_4339)
);

A2O1A1Ixp33_ASAP7_75t_L g4340 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4340)
);

A2O1A1Ixp33_ASAP7_75t_L g4341 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4342)
);

AOI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4344)
);

BUFx2_ASAP7_75t_L g4345 ( 
.A(n_2431),
.Y(n_4345)
);

CKINVDCx20_ASAP7_75t_R g4346 ( 
.A(n_2011),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_SL g4348 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4348)
);

NOR2x1_ASAP7_75t_L g4349 ( 
.A(n_2101),
.B(n_2123),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4351)
);

AOI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_SL g4353 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4353)
);

AOI21xp5_ASAP7_75t_L g4354 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4354)
);

OAI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4355)
);

AND2x4_ASAP7_75t_L g4356 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4356)
);

OAI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4358)
);

AOI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4359)
);

AOI21xp5_ASAP7_75t_L g4360 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4360)
);

AOI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4361)
);

INVx5_ASAP7_75t_L g4362 ( 
.A(n_2035),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4363)
);

OAI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4364)
);

A2O1A1Ixp33_ASAP7_75t_L g4365 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_2311),
.Y(n_4368)
);

AOI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_1968),
.A2(n_2371),
.B1(n_2375),
.B2(n_2366),
.Y(n_4369)
);

AO21x1_ASAP7_75t_L g4370 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4370)
);

AOI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4372)
);

O2A1O1Ixp33_ASAP7_75t_L g4373 ( 
.A1(n_2366),
.A2(n_1119),
.B(n_1090),
.C(n_1968),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_2074),
.B(n_2052),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_SL g4377 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4377)
);

AOI21xp33_ASAP7_75t_L g4378 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4379)
);

AO21x1_ASAP7_75t_L g4380 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4380)
);

OAI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4381)
);

AOI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4382)
);

OAI321xp33_ASAP7_75t_L g4383 ( 
.A1(n_1968),
.A2(n_1090),
.A3(n_1119),
.B1(n_2366),
.B2(n_2375),
.C(n_2371),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4384)
);

AOI21xp5_ASAP7_75t_L g4385 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4385)
);

NOR2xp33_ASAP7_75t_L g4386 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_2300),
.Y(n_4387)
);

AOI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4388)
);

AOI21x1_ASAP7_75t_L g4389 ( 
.A1(n_2123),
.A2(n_2084),
.B(n_2158),
.Y(n_4389)
);

BUFx12f_ASAP7_75t_L g4390 ( 
.A(n_2040),
.Y(n_4390)
);

INVxp67_ASAP7_75t_L g4391 ( 
.A(n_2157),
.Y(n_4391)
);

AOI21xp33_ASAP7_75t_L g4392 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_SL g4394 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4394)
);

NOR2x2_ASAP7_75t_L g4395 ( 
.A(n_2252),
.B(n_2265),
.Y(n_4395)
);

INVxp67_ASAP7_75t_SL g4396 ( 
.A(n_2122),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4397)
);

A2O1A1Ixp33_ASAP7_75t_L g4398 ( 
.A1(n_2444),
.A2(n_1013),
.B(n_1148),
.C(n_1109),
.Y(n_4398)
);

NAND2x1p5_ASAP7_75t_L g4399 ( 
.A(n_2035),
.B(n_2419),
.Y(n_4399)
);

OAI22xp5_ASAP7_75t_L g4400 ( 
.A1(n_2341),
.A2(n_1777),
.B1(n_1786),
.B2(n_1616),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4401)
);

BUFx8_ASAP7_75t_L g4402 ( 
.A(n_1965),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4403)
);

OAI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_1968),
.A2(n_2371),
.B(n_2366),
.Y(n_4404)
);

AOI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_2431),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_2311),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4408)
);

AOI21xp5_ASAP7_75t_L g4409 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4409)
);

AOI21xp5_ASAP7_75t_L g4410 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_1963),
.A2(n_2372),
.B(n_2355),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_1973),
.B(n_1958),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_2311),
.Y(n_4413)
);

AND2x6_ASAP7_75t_L g4414 ( 
.A(n_2052),
.B(n_2129),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_2787),
.A2(n_1255),
.B1(n_1533),
.B2(n_1251),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_SL g4416 ( 
.A(n_2351),
.B(n_2624),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_1968),
.B(n_2366),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_3084),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_SL g4419 ( 
.A(n_3202),
.B(n_3203),
.Y(n_4419)
);

AND2x6_ASAP7_75t_SL g4420 ( 
.A(n_3698),
.B(n_3701),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_3105),
.B(n_3106),
.Y(n_4421)
);

INVxp67_ASAP7_75t_L g4422 ( 
.A(n_3523),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_3084),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_3724),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3724),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_3223),
.B(n_3976),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_3976),
.B(n_3758),
.Y(n_4427)
);

AOI221xp5_ASAP7_75t_L g4428 ( 
.A1(n_3087),
.A2(n_3889),
.B1(n_4008),
.B2(n_3858),
.C(n_3781),
.Y(n_4428)
);

BUFx8_ASAP7_75t_SL g4429 ( 
.A(n_3168),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_3976),
.B(n_3758),
.Y(n_4430)
);

O2A1O1Ixp33_ASAP7_75t_L g4431 ( 
.A1(n_3728),
.A2(n_3747),
.B(n_3850),
.C(n_3820),
.Y(n_4431)
);

NAND2x1p5_ASAP7_75t_L g4432 ( 
.A(n_3939),
.B(n_4093),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_3762),
.B(n_3783),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_3128),
.B(n_3731),
.Y(n_4434)
);

BUFx4f_ASAP7_75t_L g4435 ( 
.A(n_3586),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_3202),
.B(n_3203),
.Y(n_4436)
);

OR2x2_ASAP7_75t_L g4437 ( 
.A(n_3138),
.B(n_3151),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_3762),
.B(n_3783),
.Y(n_4438)
);

NOR2xp33_ASAP7_75t_L g4439 ( 
.A(n_3202),
.B(n_3203),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_SL g4440 ( 
.A(n_3143),
.B(n_3187),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_3811),
.B(n_3816),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_3811),
.B(n_3816),
.Y(n_4442)
);

XNOR2xp5_ASAP7_75t_L g4443 ( 
.A(n_3121),
.B(n_3721),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_3743),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_L g4445 ( 
.A(n_4251),
.B(n_4383),
.Y(n_4445)
);

AOI22x1_ASAP7_75t_L g4446 ( 
.A1(n_3126),
.A2(n_3130),
.B1(n_3218),
.B2(n_3212),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_3966),
.B(n_3996),
.Y(n_4447)
);

INVx6_ASAP7_75t_L g4448 ( 
.A(n_3371),
.Y(n_4448)
);

NOR2x1p5_ASAP7_75t_L g4449 ( 
.A(n_3103),
.B(n_3948),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_3966),
.B(n_3996),
.Y(n_4450)
);

NAND3xp33_ASAP7_75t_L g4451 ( 
.A(n_3143),
.B(n_3189),
.C(n_3187),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_L g4452 ( 
.A1(n_3189),
.A2(n_3216),
.B1(n_3217),
.B2(n_3214),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4027),
.B(n_4134),
.Y(n_4453)
);

AOI22xp33_ASAP7_75t_L g4454 ( 
.A1(n_3214),
.A2(n_3217),
.B1(n_3216),
.B2(n_3099),
.Y(n_4454)
);

AOI22xp33_ASAP7_75t_L g4455 ( 
.A1(n_3099),
.A2(n_3165),
.B1(n_3160),
.B2(n_3181),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_3735),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_L g4457 ( 
.A(n_4251),
.B(n_4383),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4027),
.B(n_4134),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4253),
.B(n_4370),
.Y(n_4459)
);

BUFx2_ASAP7_75t_L g4460 ( 
.A(n_3773),
.Y(n_4460)
);

BUFx2_ASAP7_75t_L g4461 ( 
.A(n_3773),
.Y(n_4461)
);

INVx4_ASAP7_75t_L g4462 ( 
.A(n_3371),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_R g4463 ( 
.A(n_3542),
.B(n_3904),
.Y(n_4463)
);

AND2x4_ASAP7_75t_L g4464 ( 
.A(n_3773),
.B(n_4260),
.Y(n_4464)
);

AOI22xp33_ASAP7_75t_L g4465 ( 
.A1(n_3182),
.A2(n_3183),
.B1(n_3197),
.B2(n_3192),
.Y(n_4465)
);

AND2x2_ASAP7_75t_L g4466 ( 
.A(n_3748),
.B(n_4413),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4253),
.B(n_4370),
.Y(n_4467)
);

INVx3_ASAP7_75t_SL g4468 ( 
.A(n_3737),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4380),
.B(n_3091),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_3748),
.Y(n_4470)
);

BUFx4f_ASAP7_75t_L g4471 ( 
.A(n_3586),
.Y(n_4471)
);

AND2x4_ASAP7_75t_SL g4472 ( 
.A(n_3371),
.B(n_3441),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_SL g4473 ( 
.A(n_3201),
.B(n_3212),
.Y(n_4473)
);

INVx4_ASAP7_75t_L g4474 ( 
.A(n_3371),
.Y(n_4474)
);

INVx4_ASAP7_75t_L g4475 ( 
.A(n_3441),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_3767),
.Y(n_4476)
);

CKINVDCx5p33_ASAP7_75t_R g4477 ( 
.A(n_4031),
.Y(n_4477)
);

BUFx6f_ASAP7_75t_L g4478 ( 
.A(n_3773),
.Y(n_4478)
);

OR2x6_ASAP7_75t_L g4479 ( 
.A(n_3085),
.B(n_3726),
.Y(n_4479)
);

INVx1_ASAP7_75t_SL g4480 ( 
.A(n_3523),
.Y(n_4480)
);

NOR2xp67_ASAP7_75t_L g4481 ( 
.A(n_3357),
.B(n_3263),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4380),
.B(n_3095),
.Y(n_4482)
);

O2A1O1Ixp5_ASAP7_75t_L g4483 ( 
.A1(n_3218),
.A2(n_3119),
.B(n_3159),
.C(n_3158),
.Y(n_4483)
);

AOI22xp33_ASAP7_75t_L g4484 ( 
.A1(n_3083),
.A2(n_3751),
.B1(n_3768),
.B2(n_3750),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_3170),
.B(n_3172),
.Y(n_4485)
);

BUFx2_ASAP7_75t_SL g4486 ( 
.A(n_3982),
.Y(n_4486)
);

OR2x2_ASAP7_75t_L g4487 ( 
.A(n_3138),
.B(n_3151),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_3792),
.B(n_4292),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4322),
.B(n_4369),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_3076),
.B(n_3082),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_3076),
.B(n_3082),
.Y(n_4491)
);

AOI22xp5_ASAP7_75t_L g4492 ( 
.A1(n_3952),
.A2(n_4163),
.B1(n_3842),
.B2(n_3857),
.Y(n_4492)
);

AO22x1_ASAP7_75t_L g4493 ( 
.A1(n_3133),
.A2(n_3219),
.B1(n_3080),
.B2(n_3081),
.Y(n_4493)
);

BUFx12f_ASAP7_75t_L g4494 ( 
.A(n_3418),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_SL g4495 ( 
.A(n_3121),
.B(n_3178),
.Y(n_4495)
);

INVx1_ASAP7_75t_SL g4496 ( 
.A(n_3888),
.Y(n_4496)
);

INVx4_ASAP7_75t_L g4497 ( 
.A(n_3441),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_3086),
.B(n_3720),
.Y(n_4498)
);

NOR2xp33_ASAP7_75t_L g4499 ( 
.A(n_3170),
.B(n_3172),
.Y(n_4499)
);

AND2x4_ASAP7_75t_L g4500 ( 
.A(n_4260),
.B(n_4332),
.Y(n_4500)
);

CKINVDCx5p33_ASAP7_75t_R g4501 ( 
.A(n_3161),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_3156),
.B(n_3721),
.Y(n_4502)
);

BUFx4f_ASAP7_75t_L g4503 ( 
.A(n_3586),
.Y(n_4503)
);

BUFx6f_ASAP7_75t_L g4504 ( 
.A(n_4260),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_3793),
.A2(n_3843),
.B1(n_3894),
.B2(n_3806),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_3086),
.B(n_3720),
.Y(n_4506)
);

AOI22xp5_ASAP7_75t_L g4507 ( 
.A1(n_4358),
.A2(n_3864),
.B1(n_3893),
.B2(n_3823),
.Y(n_4507)
);

CKINVDCx5p33_ASAP7_75t_R g4508 ( 
.A(n_3161),
.Y(n_4508)
);

BUFx6f_ASAP7_75t_L g4509 ( 
.A(n_4260),
.Y(n_4509)
);

BUFx6f_ASAP7_75t_L g4510 ( 
.A(n_4332),
.Y(n_4510)
);

O2A1O1Ixp33_ASAP7_75t_L g4511 ( 
.A1(n_3856),
.A2(n_3944),
.B(n_3953),
.C(n_3870),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_3730),
.B(n_3736),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3730),
.B(n_3736),
.Y(n_4513)
);

OAI22xp5_ASAP7_75t_SL g4514 ( 
.A1(n_3235),
.A2(n_3295),
.B1(n_3316),
.B2(n_3152),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_3741),
.B(n_3759),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_3741),
.B(n_3759),
.Y(n_4516)
);

BUFx6f_ASAP7_75t_L g4517 ( 
.A(n_4332),
.Y(n_4517)
);

INVx4_ASAP7_75t_L g4518 ( 
.A(n_3441),
.Y(n_4518)
);

AND2x4_ASAP7_75t_L g4519 ( 
.A(n_4332),
.B(n_3486),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_SL g4520 ( 
.A(n_3156),
.B(n_3793),
.Y(n_4520)
);

AOI22xp33_ASAP7_75t_SL g4521 ( 
.A1(n_3133),
.A2(n_3177),
.B1(n_3188),
.B2(n_3174),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_3764),
.B(n_3772),
.Y(n_4522)
);

INVx4_ASAP7_75t_L g4523 ( 
.A(n_3982),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_3764),
.B(n_3772),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_3774),
.B(n_3775),
.Y(n_4525)
);

AO22x1_ASAP7_75t_L g4526 ( 
.A1(n_3219),
.A2(n_3080),
.B1(n_3081),
.B2(n_3075),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_3774),
.B(n_3775),
.Y(n_4527)
);

NOR2xp33_ASAP7_75t_L g4528 ( 
.A(n_3174),
.B(n_3177),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_4316),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3779),
.B(n_3780),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_3779),
.B(n_3780),
.Y(n_4531)
);

CKINVDCx5p33_ASAP7_75t_R g4532 ( 
.A(n_4316),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_3788),
.B(n_3789),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_3788),
.B(n_3789),
.Y(n_4534)
);

CKINVDCx5p33_ASAP7_75t_R g4535 ( 
.A(n_3765),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_3875),
.B(n_3902),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_3791),
.B(n_3798),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3791),
.B(n_3798),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3810),
.B(n_3819),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_3810),
.B(n_3819),
.Y(n_4540)
);

AND2x4_ASAP7_75t_L g4541 ( 
.A(n_4332),
.B(n_3488),
.Y(n_4541)
);

AO21x2_ASAP7_75t_L g4542 ( 
.A1(n_3090),
.A2(n_3096),
.B(n_3094),
.Y(n_4542)
);

AND3x1_ASAP7_75t_L g4543 ( 
.A(n_3910),
.B(n_3928),
.C(n_3917),
.Y(n_4543)
);

AND2x6_ASAP7_75t_L g4544 ( 
.A(n_3586),
.B(n_3605),
.Y(n_4544)
);

BUFx2_ASAP7_75t_L g4545 ( 
.A(n_3939),
.Y(n_4545)
);

NOR2xp33_ASAP7_75t_L g4546 ( 
.A(n_3188),
.B(n_3199),
.Y(n_4546)
);

BUFx6f_ASAP7_75t_L g4547 ( 
.A(n_4093),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3822),
.B(n_3826),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_3822),
.B(n_3826),
.Y(n_4549)
);

OR2x2_ASAP7_75t_L g4550 ( 
.A(n_3138),
.B(n_3151),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_SL g4551 ( 
.A(n_3806),
.B(n_3843),
.Y(n_4551)
);

AND2x6_ASAP7_75t_L g4552 ( 
.A(n_3586),
.B(n_3605),
.Y(n_4552)
);

INVxp33_ASAP7_75t_L g4553 ( 
.A(n_3455),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_4205),
.Y(n_4554)
);

AOI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_3957),
.A2(n_4148),
.B1(n_4117),
.B2(n_3990),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_3902),
.B(n_3919),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_SL g4557 ( 
.A(n_3542),
.B(n_3904),
.Y(n_4557)
);

INVxp67_ASAP7_75t_L g4558 ( 
.A(n_3888),
.Y(n_4558)
);

BUFx6f_ASAP7_75t_L g4559 ( 
.A(n_4177),
.Y(n_4559)
);

BUFx2_ASAP7_75t_L g4560 ( 
.A(n_4177),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_SL g4561 ( 
.A(n_3894),
.B(n_3912),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3827),
.B(n_3836),
.Y(n_4562)
);

OR2x6_ASAP7_75t_L g4563 ( 
.A(n_3085),
.B(n_3726),
.Y(n_4563)
);

NOR2xp33_ASAP7_75t_L g4564 ( 
.A(n_3199),
.B(n_3206),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_3827),
.B(n_3836),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_3837),
.B(n_3841),
.Y(n_4566)
);

BUFx2_ASAP7_75t_R g4567 ( 
.A(n_3684),
.Y(n_4567)
);

BUFx6f_ASAP7_75t_L g4568 ( 
.A(n_4335),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_3837),
.B(n_3841),
.Y(n_4569)
);

AOI22xp33_ASAP7_75t_L g4570 ( 
.A1(n_3936),
.A2(n_4084),
.B1(n_4127),
.B2(n_4098),
.Y(n_4570)
);

BUFx6f_ASAP7_75t_L g4571 ( 
.A(n_3760),
.Y(n_4571)
);

BUFx12f_ASAP7_75t_L g4572 ( 
.A(n_3418),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_SL g4573 ( 
.A(n_3912),
.B(n_4029),
.Y(n_4573)
);

OR2x2_ASAP7_75t_SL g4574 ( 
.A(n_3166),
.B(n_3755),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_3844),
.B(n_3845),
.Y(n_4575)
);

BUFx4f_ASAP7_75t_L g4576 ( 
.A(n_3586),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_3844),
.B(n_3845),
.Y(n_4577)
);

BUFx2_ASAP7_75t_L g4578 ( 
.A(n_3754),
.Y(n_4578)
);

AOI211xp5_ASAP7_75t_L g4579 ( 
.A1(n_3196),
.A2(n_3146),
.B(n_3186),
.C(n_3108),
.Y(n_4579)
);

NAND2xp33_ASAP7_75t_L g4580 ( 
.A(n_3998),
.B(n_4240),
.Y(n_4580)
);

BUFx2_ASAP7_75t_L g4581 ( 
.A(n_3754),
.Y(n_4581)
);

AOI22xp5_ASAP7_75t_L g4582 ( 
.A1(n_4207),
.A2(n_4184),
.B1(n_4214),
.B2(n_4152),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_3981),
.B(n_3986),
.Y(n_4583)
);

AND2x2_ASAP7_75t_SL g4584 ( 
.A(n_4337),
.B(n_3166),
.Y(n_4584)
);

AOI211xp5_ASAP7_75t_L g4585 ( 
.A1(n_3196),
.A2(n_3146),
.B(n_3186),
.C(n_3108),
.Y(n_4585)
);

NOR2xp33_ASAP7_75t_L g4586 ( 
.A(n_3206),
.B(n_3211),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_3848),
.B(n_3871),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_3740),
.A2(n_3744),
.B(n_3742),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_3848),
.B(n_3871),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_SL g4590 ( 
.A(n_4029),
.B(n_4054),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_3873),
.B(n_3876),
.Y(n_4591)
);

BUFx2_ASAP7_75t_L g4592 ( 
.A(n_3754),
.Y(n_4592)
);

AND2x4_ASAP7_75t_L g4593 ( 
.A(n_3520),
.B(n_3531),
.Y(n_4593)
);

CKINVDCx5p33_ASAP7_75t_R g4594 ( 
.A(n_3418),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_3873),
.B(n_3876),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_3878),
.B(n_3880),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4012),
.Y(n_4597)
);

INVx2_ASAP7_75t_SL g4598 ( 
.A(n_3982),
.Y(n_4598)
);

CKINVDCx8_ASAP7_75t_R g4599 ( 
.A(n_3631),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_L g4600 ( 
.A(n_3211),
.B(n_3213),
.Y(n_4600)
);

INVx2_ASAP7_75t_SL g4601 ( 
.A(n_3982),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_3878),
.B(n_3880),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_3895),
.B(n_3896),
.Y(n_4603)
);

BUFx2_ASAP7_75t_L g4604 ( 
.A(n_3754),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_3895),
.B(n_3896),
.Y(n_4605)
);

AOI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_3740),
.A2(n_3744),
.B(n_3742),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_3897),
.B(n_3899),
.Y(n_4607)
);

AND2x6_ASAP7_75t_L g4608 ( 
.A(n_3605),
.B(n_3129),
.Y(n_4608)
);

BUFx6f_ASAP7_75t_L g4609 ( 
.A(n_4266),
.Y(n_4609)
);

AOI22xp5_ASAP7_75t_L g4610 ( 
.A1(n_4386),
.A2(n_4314),
.B1(n_4412),
.B2(n_4301),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_3897),
.B(n_3899),
.Y(n_4611)
);

BUFx6f_ASAP7_75t_L g4612 ( 
.A(n_3930),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_SL g4613 ( 
.A(n_4054),
.B(n_4123),
.Y(n_4613)
);

INVx3_ASAP7_75t_L g4614 ( 
.A(n_3771),
.Y(n_4614)
);

AOI22x1_ASAP7_75t_L g4615 ( 
.A1(n_3110),
.A2(n_3112),
.B1(n_3093),
.B2(n_3075),
.Y(n_4615)
);

O2A1O1Ixp33_ASAP7_75t_L g4616 ( 
.A1(n_3994),
.A2(n_4090),
.B(n_4109),
.C(n_4070),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_3913),
.B(n_3915),
.Y(n_4617)
);

INVx2_ASAP7_75t_SL g4618 ( 
.A(n_4362),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_3913),
.B(n_3915),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_3918),
.B(n_3925),
.Y(n_4620)
);

AOI22xp33_ASAP7_75t_L g4621 ( 
.A1(n_3920),
.A2(n_4258),
.B1(n_4296),
.B2(n_4189),
.Y(n_4621)
);

BUFx2_ASAP7_75t_L g4622 ( 
.A(n_3771),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_3812),
.Y(n_4623)
);

BUFx8_ASAP7_75t_SL g4624 ( 
.A(n_3284),
.Y(n_4624)
);

BUFx2_ASAP7_75t_L g4625 ( 
.A(n_3771),
.Y(n_4625)
);

AOI22xp33_ASAP7_75t_L g4626 ( 
.A1(n_3920),
.A2(n_4258),
.B1(n_4296),
.B2(n_4189),
.Y(n_4626)
);

OAI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_4123),
.A2(n_4159),
.B1(n_4304),
.B2(n_4297),
.Y(n_4627)
);

NOR2xp33_ASAP7_75t_L g4628 ( 
.A(n_3213),
.B(n_4159),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4064),
.B(n_4075),
.Y(n_4629)
);

AOI22xp5_ASAP7_75t_L g4630 ( 
.A1(n_4415),
.A2(n_4304),
.B1(n_4307),
.B2(n_4297),
.Y(n_4630)
);

BUFx2_ASAP7_75t_L g4631 ( 
.A(n_3771),
.Y(n_4631)
);

INVx2_ASAP7_75t_SL g4632 ( 
.A(n_4362),
.Y(n_4632)
);

NOR2xp33_ASAP7_75t_L g4633 ( 
.A(n_4307),
.B(n_4405),
.Y(n_4633)
);

INVxp33_ASAP7_75t_L g4634 ( 
.A(n_3591),
.Y(n_4634)
);

NOR2xp67_ASAP7_75t_L g4635 ( 
.A(n_3263),
.B(n_3442),
.Y(n_4635)
);

CKINVDCx20_ASAP7_75t_R g4636 ( 
.A(n_3379),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4129),
.B(n_4140),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_3797),
.B(n_3833),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_3918),
.B(n_3925),
.Y(n_4639)
);

AND3x2_ASAP7_75t_SL g4640 ( 
.A(n_3176),
.B(n_4337),
.C(n_4270),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_3934),
.B(n_3935),
.Y(n_4641)
);

AOI221xp5_ASAP7_75t_L g4642 ( 
.A1(n_4315),
.A2(n_4378),
.B1(n_4392),
.B2(n_4146),
.C(n_3954),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_SL g4643 ( 
.A(n_4405),
.B(n_4415),
.Y(n_4643)
);

AND2x4_ASAP7_75t_L g4644 ( 
.A(n_3797),
.B(n_3833),
.Y(n_4644)
);

NOR2xp67_ASAP7_75t_L g4645 ( 
.A(n_3120),
.B(n_3236),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_3934),
.B(n_3935),
.Y(n_4646)
);

INVx2_ASAP7_75t_SL g4647 ( 
.A(n_4362),
.Y(n_4647)
);

NOR2xp33_ASAP7_75t_L g4648 ( 
.A(n_3734),
.B(n_4227),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_3937),
.B(n_3941),
.Y(n_4649)
);

INVx3_ASAP7_75t_L g4650 ( 
.A(n_3797),
.Y(n_4650)
);

BUFx6f_ASAP7_75t_L g4651 ( 
.A(n_3760),
.Y(n_4651)
);

CKINVDCx12_ASAP7_75t_R g4652 ( 
.A(n_3306),
.Y(n_4652)
);

NOR3xp33_ASAP7_75t_L g4653 ( 
.A(n_4278),
.B(n_4191),
.C(n_3755),
.Y(n_4653)
);

AND2x4_ASAP7_75t_L g4654 ( 
.A(n_3797),
.B(n_3833),
.Y(n_4654)
);

BUFx2_ASAP7_75t_L g4655 ( 
.A(n_3797),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_3937),
.B(n_3941),
.Y(n_4656)
);

OAI22xp33_ASAP7_75t_L g4657 ( 
.A1(n_3734),
.A2(n_4242),
.B1(n_4298),
.B2(n_4227),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_3950),
.B(n_3951),
.Y(n_4658)
);

AOI22xp33_ASAP7_75t_L g4659 ( 
.A1(n_3794),
.A2(n_3813),
.B1(n_3877),
.B2(n_3847),
.Y(n_4659)
);

AND2x4_ASAP7_75t_L g4660 ( 
.A(n_3833),
.B(n_3916),
.Y(n_4660)
);

O2A1O1Ixp33_ASAP7_75t_L g4661 ( 
.A1(n_4147),
.A2(n_4195),
.B(n_4275),
.C(n_4180),
.Y(n_4661)
);

BUFx6f_ASAP7_75t_L g4662 ( 
.A(n_4266),
.Y(n_4662)
);

INVxp67_ASAP7_75t_L g4663 ( 
.A(n_4099),
.Y(n_4663)
);

BUFx4f_ASAP7_75t_L g4664 ( 
.A(n_3179),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_4389),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_3950),
.B(n_3951),
.Y(n_4666)
);

NOR2xp33_ASAP7_75t_R g4667 ( 
.A(n_3184),
.B(n_3814),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_3916),
.B(n_4053),
.Y(n_4668)
);

AOI22xp5_ASAP7_75t_L g4669 ( 
.A1(n_3794),
.A2(n_3847),
.B1(n_3877),
.B2(n_3813),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_3961),
.B(n_3963),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_3961),
.B(n_3963),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4153),
.B(n_4178),
.Y(n_4672)
);

INVx1_ASAP7_75t_SL g4673 ( 
.A(n_4099),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_3916),
.B(n_4053),
.Y(n_4674)
);

BUFx6f_ASAP7_75t_L g4675 ( 
.A(n_3947),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_3965),
.B(n_3967),
.Y(n_4676)
);

INVxp67_ASAP7_75t_SL g4677 ( 
.A(n_4264),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_3965),
.B(n_3967),
.Y(n_4678)
);

BUFx6f_ASAP7_75t_L g4679 ( 
.A(n_3947),
.Y(n_4679)
);

INVx6_ASAP7_75t_L g4680 ( 
.A(n_4362),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_3970),
.B(n_3971),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_3970),
.B(n_3971),
.Y(n_4682)
);

INVx2_ASAP7_75t_SL g4683 ( 
.A(n_4362),
.Y(n_4683)
);

BUFx6f_ASAP7_75t_L g4684 ( 
.A(n_3984),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_3972),
.B(n_3978),
.Y(n_4685)
);

BUFx6f_ASAP7_75t_L g4686 ( 
.A(n_3984),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4286),
.B(n_4300),
.Y(n_4687)
);

NOR2xp33_ASAP7_75t_L g4688 ( 
.A(n_4242),
.B(n_4298),
.Y(n_4688)
);

INVxp67_ASAP7_75t_L g4689 ( 
.A(n_4103),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_3972),
.B(n_3978),
.Y(n_4690)
);

AND2x4_ASAP7_75t_L g4691 ( 
.A(n_3916),
.B(n_4053),
.Y(n_4691)
);

OR2x2_ASAP7_75t_L g4692 ( 
.A(n_3176),
.B(n_3142),
.Y(n_4692)
);

BUFx6f_ASAP7_75t_L g4693 ( 
.A(n_4389),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_3992),
.B(n_3995),
.Y(n_4694)
);

OAI22xp33_ASAP7_75t_L g4695 ( 
.A1(n_3942),
.A2(n_4003),
.B1(n_4055),
.B2(n_4024),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_3992),
.B(n_3995),
.Y(n_4696)
);

INVx5_ASAP7_75t_L g4697 ( 
.A(n_4362),
.Y(n_4697)
);

CKINVDCx8_ASAP7_75t_R g4698 ( 
.A(n_3631),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_SL g4699 ( 
.A(n_3235),
.B(n_4337),
.Y(n_4699)
);

INVxp67_ASAP7_75t_SL g4700 ( 
.A(n_4300),
.Y(n_4700)
);

AOI22xp33_ASAP7_75t_L g4701 ( 
.A1(n_3942),
.A2(n_4003),
.B1(n_4055),
.B2(n_4024),
.Y(n_4701)
);

AND2x4_ASAP7_75t_L g4702 ( 
.A(n_4053),
.B(n_4181),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_3622),
.Y(n_4703)
);

INVxp67_ASAP7_75t_L g4704 ( 
.A(n_4103),
.Y(n_4704)
);

CKINVDCx5p33_ASAP7_75t_R g4705 ( 
.A(n_3622),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_3999),
.B(n_4002),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_3999),
.B(n_4002),
.Y(n_4707)
);

CKINVDCx5p33_ASAP7_75t_R g4708 ( 
.A(n_3622),
.Y(n_4708)
);

INVx4_ASAP7_75t_L g4709 ( 
.A(n_4362),
.Y(n_4709)
);

INVx2_ASAP7_75t_SL g4710 ( 
.A(n_4053),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4006),
.B(n_4010),
.Y(n_4711)
);

OR2x6_ASAP7_75t_L g4712 ( 
.A(n_3745),
.B(n_3763),
.Y(n_4712)
);

OAI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4280),
.A2(n_4313),
.B(n_4303),
.Y(n_4713)
);

BUFx4f_ASAP7_75t_L g4714 ( 
.A(n_3179),
.Y(n_4714)
);

OR2x6_ASAP7_75t_L g4715 ( 
.A(n_3745),
.B(n_3763),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_4006),
.B(n_4010),
.Y(n_4716)
);

AOI22xp5_ASAP7_75t_L g4717 ( 
.A1(n_4116),
.A2(n_4157),
.B1(n_4158),
.B2(n_4150),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_SL g4718 ( 
.A(n_3235),
.B(n_3885),
.Y(n_4718)
);

HB1xp67_ASAP7_75t_L g4719 ( 
.A(n_3738),
.Y(n_4719)
);

OAI22xp5_ASAP7_75t_L g4720 ( 
.A1(n_3200),
.A2(n_3210),
.B1(n_3239),
.B2(n_3209),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4015),
.B(n_4019),
.Y(n_4721)
);

INVx3_ASAP7_75t_L g4722 ( 
.A(n_4053),
.Y(n_4722)
);

BUFx12f_ASAP7_75t_L g4723 ( 
.A(n_3796),
.Y(n_4723)
);

CKINVDCx14_ASAP7_75t_R g4724 ( 
.A(n_3340),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4015),
.B(n_4019),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4022),
.B(n_4025),
.Y(n_4726)
);

INVx1_ASAP7_75t_SL g4727 ( 
.A(n_4204),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4022),
.B(n_4025),
.Y(n_4728)
);

NAND2x1_ASAP7_75t_L g4729 ( 
.A(n_3191),
.B(n_3723),
.Y(n_4729)
);

INVxp67_ASAP7_75t_L g4730 ( 
.A(n_4204),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_3769),
.A2(n_3778),
.B(n_3777),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4048),
.Y(n_4732)
);

HB1xp67_ASAP7_75t_L g4733 ( 
.A(n_3738),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4034),
.B(n_4039),
.Y(n_4734)
);

AOI22xp33_ASAP7_75t_L g4735 ( 
.A1(n_4116),
.A2(n_4150),
.B1(n_4158),
.B2(n_4157),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_3725),
.B(n_3756),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_3867),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_3867),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4034),
.B(n_4039),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_SL g4740 ( 
.A(n_3932),
.B(n_3985),
.Y(n_4740)
);

BUFx6f_ASAP7_75t_L g4741 ( 
.A(n_3809),
.Y(n_4741)
);

AND3x1_ASAP7_75t_L g4742 ( 
.A(n_3169),
.B(n_3277),
.C(n_3257),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_3749),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_3924),
.Y(n_4744)
);

INVxp67_ASAP7_75t_L g4745 ( 
.A(n_4213),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_3924),
.Y(n_4746)
);

BUFx6f_ASAP7_75t_L g4747 ( 
.A(n_3956),
.Y(n_4747)
);

AND2x6_ASAP7_75t_L g4748 ( 
.A(n_3605),
.B(n_3129),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_3725),
.B(n_3756),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4065),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_SL g4751 ( 
.A(n_3987),
.B(n_4017),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4048),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_3962),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4047),
.B(n_4049),
.Y(n_4754)
);

NAND2xp33_ASAP7_75t_SL g4755 ( 
.A(n_3103),
.B(n_3948),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_3830),
.Y(n_4756)
);

AOI22xp5_ASAP7_75t_L g4757 ( 
.A1(n_4199),
.A2(n_4357),
.B1(n_4400),
.B2(n_4289),
.Y(n_4757)
);

AOI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4199),
.A2(n_4357),
.B1(n_4400),
.B2(n_4289),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_SL g4759 ( 
.A(n_4052),
.B(n_4068),
.Y(n_4759)
);

NOR2xp67_ASAP7_75t_L g4760 ( 
.A(n_3131),
.B(n_3150),
.Y(n_4760)
);

HB1xp67_ASAP7_75t_L g4761 ( 
.A(n_3761),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4047),
.B(n_4049),
.Y(n_4762)
);

NOR2xp67_ASAP7_75t_L g4763 ( 
.A(n_3157),
.B(n_3243),
.Y(n_4763)
);

INVx1_ASAP7_75t_SL g4764 ( 
.A(n_4213),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4050),
.B(n_4057),
.Y(n_4765)
);

AO221x2_ASAP7_75t_L g4766 ( 
.A1(n_3229),
.A2(n_4278),
.B1(n_4191),
.B2(n_3118),
.C(n_3815),
.Y(n_4766)
);

A2O1A1Ixp33_ASAP7_75t_L g4767 ( 
.A1(n_3729),
.A2(n_3752),
.B(n_3805),
.C(n_3746),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4050),
.B(n_4057),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4059),
.B(n_4063),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4059),
.B(n_4063),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_3818),
.Y(n_4771)
);

OAI22xp5_ASAP7_75t_L g4772 ( 
.A1(n_3290),
.A2(n_3350),
.B1(n_3351),
.B2(n_3319),
.Y(n_4772)
);

NAND2xp33_ASAP7_75t_L g4773 ( 
.A(n_4319),
.B(n_4333),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_3818),
.Y(n_4774)
);

BUFx6f_ASAP7_75t_SL g4775 ( 
.A(n_3191),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_3830),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_SL g4777 ( 
.A(n_3078),
.B(n_3140),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_3866),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4028),
.Y(n_4779)
);

INVx4_ASAP7_75t_L g4780 ( 
.A(n_3280),
.Y(n_4780)
);

AOI22xp33_ASAP7_75t_L g4781 ( 
.A1(n_3757),
.A2(n_4416),
.B1(n_3074),
.B2(n_3727),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4067),
.B(n_4073),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_3866),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_SL g4784 ( 
.A(n_3093),
.B(n_3787),
.Y(n_4784)
);

AND2x4_ASAP7_75t_L g4785 ( 
.A(n_4212),
.B(n_4228),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4067),
.B(n_4073),
.Y(n_4786)
);

AOI22xp5_ASAP7_75t_L g4787 ( 
.A1(n_3722),
.A2(n_3824),
.B1(n_3849),
.B2(n_3804),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4085),
.B(n_4097),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4085),
.B(n_4097),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_3881),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4115),
.B(n_4118),
.Y(n_4791)
);

HB1xp67_ASAP7_75t_L g4792 ( 
.A(n_3881),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_3921),
.Y(n_4793)
);

HB1xp67_ASAP7_75t_L g4794 ( 
.A(n_3921),
.Y(n_4794)
);

INVx2_ASAP7_75t_L g4795 ( 
.A(n_3938),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4115),
.B(n_4118),
.Y(n_4796)
);

OR2x4_ASAP7_75t_L g4797 ( 
.A(n_3134),
.B(n_3154),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4120),
.B(n_4132),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4120),
.B(n_4132),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_L g4800 ( 
.A(n_4133),
.B(n_4135),
.Y(n_4800)
);

INVx1_ASAP7_75t_SL g4801 ( 
.A(n_4243),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_3766),
.B(n_3770),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_3938),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4133),
.B(n_4135),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_3766),
.B(n_3770),
.Y(n_4805)
);

OAI21xp5_ASAP7_75t_L g4806 ( 
.A1(n_4340),
.A2(n_4365),
.B(n_4341),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_3198),
.B(n_3124),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_3776),
.B(n_3808),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_3962),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_L g4810 ( 
.A(n_3198),
.B(n_3124),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4136),
.B(n_4137),
.Y(n_4811)
);

NOR2xp33_ASAP7_75t_L g4812 ( 
.A(n_3125),
.B(n_3954),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_3977),
.Y(n_4813)
);

BUFx4f_ASAP7_75t_L g4814 ( 
.A(n_3179),
.Y(n_4814)
);

OR2x2_ASAP7_75t_L g4815 ( 
.A(n_3176),
.B(n_3142),
.Y(n_4815)
);

NOR2xp33_ASAP7_75t_L g4816 ( 
.A(n_3125),
.B(n_4146),
.Y(n_4816)
);

OR2x4_ASAP7_75t_L g4817 ( 
.A(n_3134),
.B(n_3154),
.Y(n_4817)
);

INVx3_ASAP7_75t_L g4818 ( 
.A(n_4228),
.Y(n_4818)
);

BUFx6f_ASAP7_75t_L g4819 ( 
.A(n_4228),
.Y(n_4819)
);

INVx4_ASAP7_75t_L g4820 ( 
.A(n_3280),
.Y(n_4820)
);

AOI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_3769),
.A2(n_3778),
.B(n_3777),
.Y(n_4821)
);

INVxp67_ASAP7_75t_SL g4822 ( 
.A(n_4407),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_3776),
.B(n_3808),
.Y(n_4823)
);

AOI22xp33_ASAP7_75t_L g4824 ( 
.A1(n_3863),
.A2(n_3890),
.B1(n_3892),
.B2(n_3883),
.Y(n_4824)
);

BUFx6f_ASAP7_75t_L g4825 ( 
.A(n_4267),
.Y(n_4825)
);

OAI221xp5_ASAP7_75t_L g4826 ( 
.A1(n_4398),
.A2(n_3113),
.B1(n_3092),
.B2(n_3089),
.C(n_3787),
.Y(n_4826)
);

HB1xp67_ASAP7_75t_L g4827 ( 
.A(n_3980),
.Y(n_4827)
);

AND2x4_ASAP7_75t_L g4828 ( 
.A(n_4267),
.B(n_4273),
.Y(n_4828)
);

AND2x4_ASAP7_75t_L g4829 ( 
.A(n_4267),
.B(n_4273),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_L g4830 ( 
.A(n_4136),
.B(n_4137),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_3980),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4001),
.Y(n_4832)
);

AOI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_3903),
.A2(n_3922),
.B1(n_3991),
.B2(n_3909),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4001),
.Y(n_4834)
);

CKINVDCx20_ASAP7_75t_R g4835 ( 
.A(n_3800),
.Y(n_4835)
);

AOI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4042),
.A2(n_4060),
.B1(n_4106),
.B2(n_4043),
.Y(n_4836)
);

AOI22xp5_ASAP7_75t_L g4837 ( 
.A1(n_4165),
.A2(n_4202),
.B1(n_4226),
.B2(n_4187),
.Y(n_4837)
);

INVxp67_ASAP7_75t_L g4838 ( 
.A(n_4243),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4139),
.B(n_4151),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_SL g4840 ( 
.A(n_3815),
.B(n_3859),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4139),
.B(n_4151),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4013),
.Y(n_4842)
);

CKINVDCx5p33_ASAP7_75t_R g4843 ( 
.A(n_3284),
.Y(n_4843)
);

BUFx6f_ASAP7_75t_L g4844 ( 
.A(n_4273),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4156),
.B(n_4161),
.Y(n_4845)
);

AO22x1_ASAP7_75t_L g4846 ( 
.A1(n_3859),
.A2(n_3874),
.B1(n_3914),
.B2(n_3905),
.Y(n_4846)
);

INVx1_ASAP7_75t_SL g4847 ( 
.A(n_4256),
.Y(n_4847)
);

A2O1A1Ixp33_ASAP7_75t_L g4848 ( 
.A1(n_3821),
.A2(n_3898),
.B(n_3927),
.C(n_3882),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4378),
.B(n_4392),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_3835),
.B(n_3846),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4028),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4044),
.Y(n_4852)
);

AOI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4274),
.A2(n_4287),
.B1(n_4317),
.B2(n_4281),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4156),
.B(n_4161),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_3835),
.B(n_3846),
.Y(n_4855)
);

NOR2xp67_ASAP7_75t_L g4856 ( 
.A(n_3115),
.B(n_3267),
.Y(n_4856)
);

OR2x6_ASAP7_75t_L g4857 ( 
.A(n_3782),
.B(n_3784),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4044),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4062),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4166),
.B(n_4169),
.Y(n_4860)
);

INVx3_ASAP7_75t_SL g4861 ( 
.A(n_4395),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4081),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4221),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4221),
.Y(n_4864)
);

AND2x6_ASAP7_75t_L g4865 ( 
.A(n_3129),
.B(n_3190),
.Y(n_4865)
);

INVx4_ASAP7_75t_L g4866 ( 
.A(n_3280),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4279),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4081),
.Y(n_4868)
);

NOR2xp33_ASAP7_75t_SL g4869 ( 
.A(n_3358),
.B(n_3316),
.Y(n_4869)
);

INVx1_ASAP7_75t_SL g4870 ( 
.A(n_4256),
.Y(n_4870)
);

INVx2_ASAP7_75t_SL g4871 ( 
.A(n_4285),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4166),
.B(n_4169),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4112),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_3886),
.B(n_3901),
.Y(n_4874)
);

INVx2_ASAP7_75t_L g4875 ( 
.A(n_4105),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4339),
.Y(n_4876)
);

INVxp67_ASAP7_75t_L g4877 ( 
.A(n_4345),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4174),
.B(n_4182),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4339),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4368),
.Y(n_4880)
);

AND3x1_ASAP7_75t_SL g4881 ( 
.A(n_3262),
.B(n_4348),
.C(n_4325),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_3886),
.B(n_3901),
.Y(n_4882)
);

OR2x6_ASAP7_75t_L g4883 ( 
.A(n_3782),
.B(n_3784),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_SL g4884 ( 
.A(n_3358),
.B(n_3316),
.Y(n_4884)
);

INVx5_ASAP7_75t_L g4885 ( 
.A(n_3129),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_4112),
.Y(n_4886)
);

CKINVDCx5p33_ASAP7_75t_R g4887 ( 
.A(n_3284),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_L g4888 ( 
.A(n_3167),
.B(n_4174),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4182),
.B(n_4192),
.Y(n_4889)
);

OR2x6_ASAP7_75t_L g4890 ( 
.A(n_3785),
.B(n_3786),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4192),
.B(n_4194),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_SL g4892 ( 
.A(n_3874),
.B(n_3905),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_SL g4893 ( 
.A(n_3914),
.B(n_3929),
.Y(n_4893)
);

OR2x6_ASAP7_75t_SL g4894 ( 
.A(n_3144),
.B(n_3145),
.Y(n_4894)
);

AOI21xp5_ASAP7_75t_L g4895 ( 
.A1(n_3785),
.A2(n_3795),
.B(n_3786),
.Y(n_4895)
);

NOR2xp67_ASAP7_75t_L g4896 ( 
.A(n_3267),
.B(n_3276),
.Y(n_4896)
);

AOI21xp5_ASAP7_75t_L g4897 ( 
.A1(n_3795),
.A2(n_3802),
.B(n_3801),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_L g4898 ( 
.A(n_4194),
.B(n_4200),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4200),
.B(n_4206),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_L g4900 ( 
.A(n_4206),
.B(n_4210),
.Y(n_4900)
);

NOR2xp67_ASAP7_75t_L g4901 ( 
.A(n_3276),
.B(n_3248),
.Y(n_4901)
);

HB1xp67_ASAP7_75t_L g4902 ( 
.A(n_4241),
.Y(n_4902)
);

INVx1_ASAP7_75t_SL g4903 ( 
.A(n_4345),
.Y(n_4903)
);

AOI221xp5_ASAP7_75t_L g4904 ( 
.A1(n_4077),
.A2(n_4171),
.B1(n_4237),
.B2(n_4167),
.C(n_4155),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_3417),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4210),
.B(n_4216),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_3417),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_3429),
.Y(n_4908)
);

CKINVDCx5p33_ASAP7_75t_R g4909 ( 
.A(n_3302),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_L g4910 ( 
.A1(n_4353),
.A2(n_4394),
.B1(n_4377),
.B2(n_4005),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4216),
.B(n_4217),
.Y(n_4911)
);

INVx4_ASAP7_75t_L g4912 ( 
.A(n_3280),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_L g4913 ( 
.A(n_3167),
.B(n_4217),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4218),
.B(n_4225),
.Y(n_4914)
);

O2A1O1Ixp33_ASAP7_75t_L g4915 ( 
.A1(n_4373),
.A2(n_3929),
.B(n_3940),
.C(n_3933),
.Y(n_4915)
);

INVx2_ASAP7_75t_L g4916 ( 
.A(n_3429),
.Y(n_4916)
);

HB1xp67_ASAP7_75t_L g4917 ( 
.A(n_3195),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4218),
.B(n_4225),
.Y(n_4918)
);

HB1xp67_ASAP7_75t_L g4919 ( 
.A(n_3195),
.Y(n_4919)
);

AND2x4_ASAP7_75t_L g4920 ( 
.A(n_4387),
.B(n_3098),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_3569),
.Y(n_4921)
);

NOR2xp33_ASAP7_75t_L g4922 ( 
.A(n_4229),
.B(n_4231),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4229),
.B(n_4231),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_3969),
.A2(n_4033),
.B1(n_4036),
.B2(n_4005),
.Y(n_4924)
);

INVx4_ASAP7_75t_L g4925 ( 
.A(n_3280),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4232),
.B(n_4235),
.Y(n_4926)
);

INVx2_ASAP7_75t_SL g4927 ( 
.A(n_4387),
.Y(n_4927)
);

AND2x4_ASAP7_75t_L g4928 ( 
.A(n_4387),
.B(n_3098),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_3569),
.Y(n_4929)
);

HB1xp67_ASAP7_75t_L g4930 ( 
.A(n_3195),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4232),
.B(n_4235),
.Y(n_4931)
);

INVx2_ASAP7_75t_SL g4932 ( 
.A(n_4387),
.Y(n_4932)
);

INVx4_ASAP7_75t_L g4933 ( 
.A(n_3129),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4238),
.B(n_4244),
.Y(n_4934)
);

NOR2xp33_ASAP7_75t_L g4935 ( 
.A(n_4238),
.B(n_4244),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4246),
.B(n_4247),
.Y(n_4936)
);

AOI22x1_ASAP7_75t_L g4937 ( 
.A1(n_4404),
.A2(n_3933),
.B1(n_3997),
.B2(n_3940),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4246),
.B(n_4247),
.Y(n_4938)
);

AOI21xp5_ASAP7_75t_L g4939 ( 
.A1(n_3801),
.A2(n_3803),
.B(n_3802),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_3969),
.B(n_4033),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_3141),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4252),
.B(n_4255),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_3141),
.Y(n_4943)
);

BUFx12f_ASAP7_75t_L g4944 ( 
.A(n_3796),
.Y(n_4944)
);

BUFx6f_ASAP7_75t_L g4945 ( 
.A(n_3098),
.Y(n_4945)
);

INVx2_ASAP7_75t_SL g4946 ( 
.A(n_3129),
.Y(n_4946)
);

OAI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_3097),
.A2(n_3101),
.B1(n_3111),
.B2(n_3109),
.Y(n_4947)
);

INVx5_ASAP7_75t_L g4948 ( 
.A(n_3190),
.Y(n_4948)
);

BUFx6f_ASAP7_75t_L g4949 ( 
.A(n_3098),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4252),
.B(n_4255),
.Y(n_4950)
);

AND2x4_ASAP7_75t_L g4951 ( 
.A(n_3733),
.B(n_3852),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_SL g4952 ( 
.A(n_3997),
.B(n_4007),
.Y(n_4952)
);

INVx2_ASAP7_75t_SL g4953 ( 
.A(n_3190),
.Y(n_4953)
);

AOI22x1_ASAP7_75t_L g4954 ( 
.A1(n_4404),
.A2(n_4007),
.B1(n_4072),
.B2(n_4051),
.Y(n_4954)
);

AOI211xp5_ASAP7_75t_L g4955 ( 
.A1(n_3221),
.A2(n_3339),
.B(n_3249),
.C(n_3320),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_4051),
.B(n_4072),
.Y(n_4956)
);

INVx2_ASAP7_75t_SL g4957 ( 
.A(n_3190),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_3302),
.Y(n_4958)
);

BUFx6f_ASAP7_75t_L g4959 ( 
.A(n_3733),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4036),
.B(n_4066),
.Y(n_4960)
);

BUFx3_ASAP7_75t_L g4961 ( 
.A(n_3588),
.Y(n_4961)
);

INVx6_ASAP7_75t_L g4962 ( 
.A(n_3191),
.Y(n_4962)
);

AND2x4_ASAP7_75t_L g4963 ( 
.A(n_3733),
.B(n_3834),
.Y(n_4963)
);

BUFx2_ASAP7_75t_L g4964 ( 
.A(n_4143),
.Y(n_4964)
);

BUFx6f_ASAP7_75t_L g4965 ( 
.A(n_3834),
.Y(n_4965)
);

BUFx4f_ASAP7_75t_L g4966 ( 
.A(n_4004),
.Y(n_4966)
);

INVx4_ASAP7_75t_L g4967 ( 
.A(n_3190),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4257),
.B(n_4263),
.Y(n_4968)
);

BUFx3_ASAP7_75t_L g4969 ( 
.A(n_3588),
.Y(n_4969)
);

NAND2xp5_ASAP7_75t_L g4970 ( 
.A(n_4257),
.B(n_4263),
.Y(n_4970)
);

INVx3_ASAP7_75t_L g4971 ( 
.A(n_3834),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4265),
.B(n_4293),
.Y(n_4972)
);

INVx3_ASAP7_75t_SL g4973 ( 
.A(n_3642),
.Y(n_4973)
);

AND2x4_ASAP7_75t_L g4974 ( 
.A(n_3852),
.B(n_4018),
.Y(n_4974)
);

AOI22xp5_ASAP7_75t_L g4975 ( 
.A1(n_3321),
.A2(n_3362),
.B1(n_3339),
.B2(n_3221),
.Y(n_4975)
);

BUFx3_ASAP7_75t_L g4976 ( 
.A(n_3522),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4265),
.B(n_4293),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4306),
.B(n_4309),
.Y(n_4978)
);

BUFx2_ASAP7_75t_L g4979 ( 
.A(n_4143),
.Y(n_4979)
);

BUFx6f_ASAP7_75t_L g4980 ( 
.A(n_3852),
.Y(n_4980)
);

OR2x2_ASAP7_75t_L g4981 ( 
.A(n_3144),
.B(n_3145),
.Y(n_4981)
);

BUFx4f_ASAP7_75t_SL g4982 ( 
.A(n_3302),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4066),
.B(n_4124),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4306),
.B(n_4309),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4310),
.B(n_4312),
.Y(n_4985)
);

INVx5_ASAP7_75t_L g4986 ( 
.A(n_3190),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_3310),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4310),
.B(n_4312),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4124),
.B(n_4131),
.Y(n_4989)
);

CKINVDCx20_ASAP7_75t_R g4990 ( 
.A(n_4346),
.Y(n_4990)
);

AOI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4131),
.A2(n_4190),
.B1(n_4203),
.B2(n_4160),
.Y(n_4991)
);

A2O1A1Ixp33_ASAP7_75t_L g4992 ( 
.A1(n_4284),
.A2(n_3118),
.B(n_4172),
.C(n_4083),
.Y(n_4992)
);

OAI22xp5_ASAP7_75t_L g4993 ( 
.A1(n_3117),
.A2(n_3135),
.B1(n_3163),
.B2(n_3148),
.Y(n_4993)
);

BUFx3_ASAP7_75t_L g4994 ( 
.A(n_3522),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4318),
.B(n_4321),
.Y(n_4995)
);

OAI22xp5_ASAP7_75t_L g4996 ( 
.A1(n_3180),
.A2(n_3194),
.B1(n_3222),
.B2(n_3205),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4318),
.B(n_4321),
.Y(n_4997)
);

BUFx2_ASAP7_75t_L g4998 ( 
.A(n_4149),
.Y(n_4998)
);

NOR2xp33_ASAP7_75t_L g4999 ( 
.A(n_4327),
.B(n_4328),
.Y(n_4999)
);

BUFx12f_ASAP7_75t_L g5000 ( 
.A(n_3796),
.Y(n_5000)
);

OR2x2_ASAP7_75t_L g5001 ( 
.A(n_3127),
.B(n_3155),
.Y(n_5001)
);

AOI21xp5_ASAP7_75t_L g5002 ( 
.A1(n_3803),
.A2(n_4087),
.B(n_4078),
.Y(n_5002)
);

A2O1A1Ixp33_ASAP7_75t_L g5003 ( 
.A1(n_4122),
.A2(n_4083),
.B(n_4086),
.C(n_4079),
.Y(n_5003)
);

BUFx6f_ASAP7_75t_L g5004 ( 
.A(n_3989),
.Y(n_5004)
);

BUFx6f_ASAP7_75t_L g5005 ( 
.A(n_4018),
.Y(n_5005)
);

NAND2xp5_ASAP7_75t_L g5006 ( 
.A(n_4327),
.B(n_4328),
.Y(n_5006)
);

AND2x4_ASAP7_75t_L g5007 ( 
.A(n_4018),
.B(n_4071),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_SL g5008 ( 
.A(n_4079),
.B(n_4086),
.Y(n_5008)
);

AOI22xp5_ASAP7_75t_L g5009 ( 
.A1(n_3227),
.A2(n_3265),
.B1(n_3282),
.B2(n_3275),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4330),
.B(n_4338),
.Y(n_5010)
);

INVx2_ASAP7_75t_SL g5011 ( 
.A(n_3281),
.Y(n_5011)
);

BUFx2_ASAP7_75t_L g5012 ( 
.A(n_4149),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4330),
.B(n_4338),
.Y(n_5013)
);

BUFx6f_ASAP7_75t_L g5014 ( 
.A(n_4071),
.Y(n_5014)
);

BUFx2_ASAP7_75t_L g5015 ( 
.A(n_4288),
.Y(n_5015)
);

AO22x1_ASAP7_75t_L g5016 ( 
.A1(n_4088),
.A2(n_4113),
.B1(n_4128),
.B2(n_4122),
.Y(n_5016)
);

BUFx2_ASAP7_75t_L g5017 ( 
.A(n_4288),
.Y(n_5017)
);

AND2x4_ASAP7_75t_L g5018 ( 
.A(n_4071),
.B(n_4271),
.Y(n_5018)
);

OAI22xp5_ASAP7_75t_L g5019 ( 
.A1(n_3309),
.A2(n_3311),
.B1(n_3313),
.B2(n_3312),
.Y(n_5019)
);

HB1xp67_ASAP7_75t_L g5020 ( 
.A(n_3195),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4342),
.B(n_4347),
.Y(n_5021)
);

NOR2xp33_ASAP7_75t_L g5022 ( 
.A(n_4342),
.B(n_4347),
.Y(n_5022)
);

BUFx3_ASAP7_75t_L g5023 ( 
.A(n_3522),
.Y(n_5023)
);

OR2x2_ASAP7_75t_L g5024 ( 
.A(n_3127),
.B(n_3356),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4350),
.B(n_4351),
.Y(n_5025)
);

BUFx3_ASAP7_75t_L g5026 ( 
.A(n_3522),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4350),
.B(n_4351),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4372),
.B(n_4379),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4372),
.B(n_4379),
.Y(n_5029)
);

A2O1A1Ixp33_ASAP7_75t_L g5030 ( 
.A1(n_4355),
.A2(n_4113),
.B(n_4128),
.C(n_4088),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4384),
.B(n_4397),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_3526),
.Y(n_5032)
);

INVx2_ASAP7_75t_SL g5033 ( 
.A(n_3281),
.Y(n_5033)
);

OR2x6_ASAP7_75t_L g5034 ( 
.A(n_4078),
.B(n_4087),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_3473),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_4384),
.B(n_4397),
.Y(n_5036)
);

OAI22xp5_ASAP7_75t_L g5037 ( 
.A1(n_3329),
.A2(n_3344),
.B1(n_3355),
.B2(n_3428),
.Y(n_5037)
);

NAND2xp33_ASAP7_75t_L g5038 ( 
.A(n_4144),
.B(n_4172),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_3526),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_3193),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_SL g5041 ( 
.A(n_4144),
.B(n_4196),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_3473),
.Y(n_5042)
);

INVx1_ASAP7_75t_SL g5043 ( 
.A(n_3116),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4401),
.B(n_4403),
.Y(n_5044)
);

INVx4_ASAP7_75t_L g5045 ( 
.A(n_3281),
.Y(n_5045)
);

AND3x1_ASAP7_75t_SL g5046 ( 
.A(n_3262),
.B(n_4270),
.C(n_3709),
.Y(n_5046)
);

NAND2x1p5_ASAP7_75t_L g5047 ( 
.A(n_4349),
.B(n_3104),
.Y(n_5047)
);

NOR2x1_ASAP7_75t_L g5048 ( 
.A(n_3137),
.B(n_3853),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_3193),
.Y(n_5049)
);

INVx2_ASAP7_75t_SL g5050 ( 
.A(n_3281),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4160),
.B(n_4190),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_3208),
.Y(n_5052)
);

INVxp67_ASAP7_75t_SL g5053 ( 
.A(n_3123),
.Y(n_5053)
);

HB1xp67_ASAP7_75t_L g5054 ( 
.A(n_3637),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4401),
.B(n_4403),
.Y(n_5055)
);

BUFx2_ASAP7_75t_L g5056 ( 
.A(n_4349),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4408),
.B(n_4417),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4408),
.B(n_4417),
.Y(n_5058)
);

BUFx6f_ASAP7_75t_L g5059 ( 
.A(n_4071),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_3245),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_SL g5061 ( 
.A(n_4196),
.B(n_4224),
.Y(n_5061)
);

OR2x2_ASAP7_75t_L g5062 ( 
.A(n_3356),
.B(n_3122),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4224),
.B(n_4290),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_SL g5064 ( 
.A(n_4290),
.B(n_4324),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_SL g5065 ( 
.A(n_4324),
.B(n_4329),
.Y(n_5065)
);

HB1xp67_ASAP7_75t_L g5066 ( 
.A(n_3637),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_4329),
.B(n_4355),
.Y(n_5067)
);

BUFx6f_ASAP7_75t_L g5068 ( 
.A(n_4271),
.Y(n_5068)
);

BUFx2_ASAP7_75t_L g5069 ( 
.A(n_3114),
.Y(n_5069)
);

INVx3_ASAP7_75t_L g5070 ( 
.A(n_4271),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_3245),
.Y(n_5071)
);

AND2x4_ASAP7_75t_L g5072 ( 
.A(n_4363),
.B(n_4375),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_SL g5073 ( 
.A(n_4364),
.B(n_4381),
.Y(n_5073)
);

AND3x1_ASAP7_75t_SL g5074 ( 
.A(n_3709),
.B(n_3712),
.C(n_3349),
.Y(n_5074)
);

O2A1O1Ixp33_ASAP7_75t_L g5075 ( 
.A1(n_4364),
.A2(n_4381),
.B(n_3077),
.C(n_3229),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_3251),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_3122),
.B(n_4203),
.Y(n_5077)
);

INVx4_ASAP7_75t_L g5078 ( 
.A(n_3281),
.Y(n_5078)
);

AOI22xp5_ASAP7_75t_SL g5079 ( 
.A1(n_3153),
.A2(n_4222),
.B1(n_4283),
.B2(n_4262),
.Y(n_5079)
);

BUFx6f_ASAP7_75t_L g5080 ( 
.A(n_4271),
.Y(n_5080)
);

NOR2xp33_ASAP7_75t_L g5081 ( 
.A(n_3173),
.B(n_3448),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4222),
.B(n_4262),
.Y(n_5082)
);

BUFx8_ASAP7_75t_L g5083 ( 
.A(n_3281),
.Y(n_5083)
);

BUFx12f_ASAP7_75t_L g5084 ( 
.A(n_3796),
.Y(n_5084)
);

HB1xp67_ASAP7_75t_L g5085 ( 
.A(n_3483),
.Y(n_5085)
);

A2O1A1Ixp33_ASAP7_75t_L g5086 ( 
.A1(n_3114),
.A2(n_3139),
.B(n_3264),
.C(n_3361),
.Y(n_5086)
);

AND3x2_ASAP7_75t_SL g5087 ( 
.A(n_3343),
.B(n_3147),
.C(n_3234),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_SL g5088 ( 
.A(n_3428),
.B(n_3438),
.Y(n_5088)
);

AND2x2_ASAP7_75t_L g5089 ( 
.A(n_4283),
.B(n_4305),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_3278),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_4305),
.B(n_4326),
.Y(n_5091)
);

NAND2x1p5_ASAP7_75t_L g5092 ( 
.A(n_3817),
.B(n_3825),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_4326),
.B(n_3369),
.Y(n_5093)
);

NOR3xp33_ASAP7_75t_L g5094 ( 
.A(n_3613),
.B(n_3368),
.C(n_3322),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_3348),
.Y(n_5095)
);

BUFx6f_ASAP7_75t_L g5096 ( 
.A(n_4356),
.Y(n_5096)
);

BUFx2_ASAP7_75t_L g5097 ( 
.A(n_3483),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_L g5098 ( 
.A(n_3369),
.B(n_3382),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_3359),
.Y(n_5099)
);

NOR2xp33_ASAP7_75t_L g5100 ( 
.A(n_3438),
.B(n_3318),
.Y(n_5100)
);

NAND2xp33_ASAP7_75t_L g5101 ( 
.A(n_3107),
.B(n_3164),
.Y(n_5101)
);

NOR2xp33_ASAP7_75t_L g5102 ( 
.A(n_3534),
.B(n_3136),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_3367),
.Y(n_5103)
);

BUFx6f_ASAP7_75t_L g5104 ( 
.A(n_4356),
.Y(n_5104)
);

AOI22xp33_ASAP7_75t_L g5105 ( 
.A1(n_3107),
.A2(n_3153),
.B1(n_3224),
.B2(n_3220),
.Y(n_5105)
);

NOR2xp33_ASAP7_75t_R g5106 ( 
.A(n_3184),
.B(n_3814),
.Y(n_5106)
);

NOR2xp33_ASAP7_75t_R g5107 ( 
.A(n_3838),
.B(n_3906),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_3382),
.B(n_3390),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_3102),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_3220),
.B(n_3304),
.Y(n_5110)
);

AOI22xp5_ASAP7_75t_L g5111 ( 
.A1(n_3224),
.A2(n_3458),
.B1(n_3534),
.B2(n_3376),
.Y(n_5111)
);

INVx2_ASAP7_75t_SL g5112 ( 
.A(n_3297),
.Y(n_5112)
);

BUFx6f_ASAP7_75t_L g5113 ( 
.A(n_4363),
.Y(n_5113)
);

AND2x4_ASAP7_75t_L g5114 ( 
.A(n_4363),
.B(n_4375),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_3383),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_3383),
.Y(n_5116)
);

BUFx2_ASAP7_75t_L g5117 ( 
.A(n_3415),
.Y(n_5117)
);

HB1xp67_ASAP7_75t_L g5118 ( 
.A(n_3171),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_3386),
.Y(n_5119)
);

AOI22xp33_ASAP7_75t_L g5120 ( 
.A1(n_3224),
.A2(n_3368),
.B1(n_3458),
.B2(n_3136),
.Y(n_5120)
);

BUFx2_ASAP7_75t_L g5121 ( 
.A(n_3415),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_SL g5122 ( 
.A(n_3458),
.B(n_3390),
.Y(n_5122)
);

OAI22xp5_ASAP7_75t_SL g5123 ( 
.A1(n_3684),
.A2(n_3402),
.B1(n_3642),
.B2(n_3701),
.Y(n_5123)
);

HB1xp67_ASAP7_75t_L g5124 ( 
.A(n_3204),
.Y(n_5124)
);

INVx4_ASAP7_75t_L g5125 ( 
.A(n_3297),
.Y(n_5125)
);

NOR2xp33_ASAP7_75t_L g5126 ( 
.A(n_3719),
.B(n_3304),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_3386),
.Y(n_5127)
);

NOR2xp33_ASAP7_75t_L g5128 ( 
.A(n_3719),
.B(n_3315),
.Y(n_5128)
);

BUFx3_ASAP7_75t_L g5129 ( 
.A(n_3522),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_SL g5130 ( 
.A(n_3393),
.B(n_3410),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_SL g5131 ( 
.A(n_3393),
.B(n_3410),
.Y(n_5131)
);

BUFx4f_ASAP7_75t_L g5132 ( 
.A(n_4004),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_3388),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_3372),
.B(n_3392),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_3388),
.Y(n_5135)
);

OR2x6_ASAP7_75t_L g5136 ( 
.A(n_4089),
.B(n_4091),
.Y(n_5136)
);

OAI22xp5_ASAP7_75t_L g5137 ( 
.A1(n_3401),
.A2(n_3421),
.B1(n_3391),
.B2(n_3226),
.Y(n_5137)
);

NOR2xp33_ASAP7_75t_L g5138 ( 
.A(n_3315),
.B(n_3424),
.Y(n_5138)
);

A2O1A1Ixp33_ASAP7_75t_L g5139 ( 
.A1(n_3395),
.A2(n_3405),
.B(n_3406),
.C(n_3397),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_4396),
.B(n_3424),
.Y(n_5140)
);

NOR2xp33_ASAP7_75t_L g5141 ( 
.A(n_3430),
.B(n_3364),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_3419),
.Y(n_5142)
);

INVxp67_ASAP7_75t_L g5143 ( 
.A(n_3207),
.Y(n_5143)
);

AO21x2_ASAP7_75t_L g5144 ( 
.A1(n_3090),
.A2(n_3096),
.B(n_3094),
.Y(n_5144)
);

INVx3_ASAP7_75t_L g5145 ( 
.A(n_4363),
.Y(n_5145)
);

AND2x6_ASAP7_75t_SL g5146 ( 
.A(n_3702),
.B(n_3636),
.Y(n_5146)
);

BUFx6f_ASAP7_75t_L g5147 ( 
.A(n_4375),
.Y(n_5147)
);

BUFx6f_ASAP7_75t_L g5148 ( 
.A(n_4375),
.Y(n_5148)
);

INVx3_ASAP7_75t_SL g5149 ( 
.A(n_3642),
.Y(n_5149)
);

AND2x4_ASAP7_75t_L g5150 ( 
.A(n_3271),
.B(n_3610),
.Y(n_5150)
);

AOI22x1_ASAP7_75t_L g5151 ( 
.A1(n_3828),
.A2(n_3832),
.B1(n_3839),
.B2(n_3829),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_3430),
.B(n_3443),
.Y(n_5152)
);

BUFx6f_ASAP7_75t_L g5153 ( 
.A(n_3147),
.Y(n_5153)
);

BUFx2_ASAP7_75t_L g5154 ( 
.A(n_3466),
.Y(n_5154)
);

BUFx2_ASAP7_75t_L g5155 ( 
.A(n_3466),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_3443),
.B(n_3411),
.Y(n_5156)
);

AOI22xp33_ASAP7_75t_L g5157 ( 
.A1(n_3414),
.A2(n_3425),
.B1(n_3422),
.B2(n_3343),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_3449),
.B(n_3307),
.Y(n_5158)
);

OR2x4_ASAP7_75t_L g5159 ( 
.A(n_3669),
.B(n_3297),
.Y(n_5159)
);

BUFx12f_ASAP7_75t_L g5160 ( 
.A(n_4402),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_3449),
.B(n_3307),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_3326),
.B(n_3334),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_3116),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_SL g5164 ( 
.A(n_3253),
.B(n_3254),
.Y(n_5164)
);

A2O1A1Ixp33_ASAP7_75t_L g5165 ( 
.A1(n_3365),
.A2(n_3378),
.B(n_3853),
.C(n_3137),
.Y(n_5165)
);

INVx5_ASAP7_75t_L g5166 ( 
.A(n_3297),
.Y(n_5166)
);

BUFx2_ASAP7_75t_L g5167 ( 
.A(n_3402),
.Y(n_5167)
);

NOR2xp33_ASAP7_75t_L g5168 ( 
.A(n_3492),
.B(n_3524),
.Y(n_5168)
);

NAND2xp5_ASAP7_75t_L g5169 ( 
.A(n_3326),
.B(n_3334),
.Y(n_5169)
);

BUFx4f_ASAP7_75t_L g5170 ( 
.A(n_4004),
.Y(n_5170)
);

BUFx6f_ASAP7_75t_L g5171 ( 
.A(n_3297),
.Y(n_5171)
);

BUFx2_ASAP7_75t_L g5172 ( 
.A(n_3266),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_3544),
.B(n_3481),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_SL g5174 ( 
.A(n_3258),
.B(n_3259),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_3375),
.B(n_3399),
.Y(n_5175)
);

CKINVDCx8_ASAP7_75t_R g5176 ( 
.A(n_4038),
.Y(n_5176)
);

NOR2xp33_ASAP7_75t_R g5177 ( 
.A(n_3838),
.B(n_3906),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_3225),
.B(n_3226),
.Y(n_5178)
);

BUFx3_ASAP7_75t_L g5179 ( 
.A(n_4399),
.Y(n_5179)
);

BUFx6f_ASAP7_75t_L g5180 ( 
.A(n_3297),
.Y(n_5180)
);

AOI22xp33_ASAP7_75t_L g5181 ( 
.A1(n_3325),
.A2(n_3345),
.B1(n_3404),
.B2(n_3360),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_3541),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_L g5183 ( 
.A(n_3225),
.B(n_3228),
.Y(n_5183)
);

INVx2_ASAP7_75t_SL g5184 ( 
.A(n_4399),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_3256),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_3228),
.B(n_3231),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_3256),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_3231),
.B(n_3238),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_3541),
.Y(n_5189)
);

OR2x2_ASAP7_75t_L g5190 ( 
.A(n_3444),
.B(n_3447),
.Y(n_5190)
);

A2O1A1Ixp33_ASAP7_75t_L g5191 ( 
.A1(n_4145),
.A2(n_3474),
.B(n_3472),
.C(n_4092),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_3540),
.Y(n_5192)
);

BUFx3_ASAP7_75t_L g5193 ( 
.A(n_4399),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_SL g5194 ( 
.A(n_3283),
.B(n_3289),
.Y(n_5194)
);

AOI21xp5_ASAP7_75t_L g5195 ( 
.A1(n_4089),
.A2(n_4092),
.B(n_4091),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_3238),
.B(n_3242),
.Y(n_5196)
);

INVx4_ASAP7_75t_L g5197 ( 
.A(n_3191),
.Y(n_5197)
);

BUFx3_ASAP7_75t_L g5198 ( 
.A(n_3638),
.Y(n_5198)
);

INVx2_ASAP7_75t_L g5199 ( 
.A(n_3540),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_3242),
.B(n_3244),
.Y(n_5200)
);

OR2x6_ASAP7_75t_L g5201 ( 
.A(n_4095),
.B(n_4096),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_3481),
.Y(n_5202)
);

INVx2_ASAP7_75t_SL g5203 ( 
.A(n_3723),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_SL g5204 ( 
.A(n_3292),
.B(n_3303),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_3484),
.Y(n_5205)
);

BUFx6f_ASAP7_75t_L g5206 ( 
.A(n_3346),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_SL g5207 ( 
.A(n_3308),
.B(n_3314),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_3244),
.B(n_3247),
.Y(n_5208)
);

AOI22xp33_ASAP7_75t_L g5209 ( 
.A1(n_3408),
.A2(n_3434),
.B1(n_3426),
.B2(n_3370),
.Y(n_5209)
);

NAND3xp33_ASAP7_75t_SL g5210 ( 
.A(n_3500),
.B(n_3471),
.C(n_3538),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_3544),
.B(n_3484),
.Y(n_5211)
);

AND2x2_ASAP7_75t_L g5212 ( 
.A(n_3544),
.B(n_3487),
.Y(n_5212)
);

AOI22xp33_ASAP7_75t_L g5213 ( 
.A1(n_3240),
.A2(n_3341),
.B1(n_3261),
.B2(n_3252),
.Y(n_5213)
);

AOI22xp5_ASAP7_75t_L g5214 ( 
.A1(n_3437),
.A2(n_3612),
.B1(n_3467),
.B2(n_3583),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_3403),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_3487),
.Y(n_5216)
);

NOR2x2_ASAP7_75t_L g5217 ( 
.A(n_3717),
.B(n_3674),
.Y(n_5217)
);

BUFx2_ASAP7_75t_L g5218 ( 
.A(n_3266),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_3498),
.Y(n_5219)
);

AOI22x1_ASAP7_75t_L g5220 ( 
.A1(n_3840),
.A2(n_3854),
.B1(n_3855),
.B2(n_3851),
.Y(n_5220)
);

AOI21xp5_ASAP7_75t_L g5221 ( 
.A1(n_4095),
.A2(n_4100),
.B(n_4096),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_3403),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_3498),
.Y(n_5223)
);

BUFx2_ASAP7_75t_L g5224 ( 
.A(n_3246),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_3247),
.B(n_3250),
.Y(n_5225)
);

HB1xp67_ASAP7_75t_L g5226 ( 
.A(n_3420),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_3250),
.B(n_3255),
.Y(n_5227)
);

INVx3_ASAP7_75t_L g5228 ( 
.A(n_3723),
.Y(n_5228)
);

BUFx6f_ASAP7_75t_L g5229 ( 
.A(n_3346),
.Y(n_5229)
);

BUFx6f_ASAP7_75t_L g5230 ( 
.A(n_3346),
.Y(n_5230)
);

AND2x2_ASAP7_75t_L g5231 ( 
.A(n_3499),
.B(n_3299),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_3255),
.B(n_3260),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_3299),
.B(n_3610),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_3260),
.B(n_3268),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_3268),
.B(n_3270),
.Y(n_5235)
);

CKINVDCx5p33_ASAP7_75t_R g5236 ( 
.A(n_3310),
.Y(n_5236)
);

AND2x2_ASAP7_75t_L g5237 ( 
.A(n_3610),
.B(n_3614),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_3550),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_3550),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_3270),
.B(n_3272),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_3530),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_3554),
.Y(n_5242)
);

NAND2xp33_ASAP7_75t_L g5243 ( 
.A(n_3272),
.B(n_3273),
.Y(n_5243)
);

INVx3_ASAP7_75t_L g5244 ( 
.A(n_3723),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_3273),
.B(n_3274),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_3274),
.B(n_3279),
.Y(n_5246)
);

NOR2xp33_ASAP7_75t_L g5247 ( 
.A(n_3492),
.B(n_3524),
.Y(n_5247)
);

INVxp33_ASAP7_75t_L g5248 ( 
.A(n_3549),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_3554),
.Y(n_5249)
);

AND2x4_ASAP7_75t_L g5250 ( 
.A(n_3271),
.B(n_3614),
.Y(n_5250)
);

INVx2_ASAP7_75t_SL g5251 ( 
.A(n_3865),
.Y(n_5251)
);

NOR2xp33_ASAP7_75t_L g5252 ( 
.A(n_3491),
.B(n_3279),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_3287),
.B(n_3288),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_3287),
.B(n_3288),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_3291),
.B(n_3293),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_3291),
.B(n_3293),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_3294),
.B(n_3298),
.Y(n_5257)
);

OAI22xp5_ASAP7_75t_SL g5258 ( 
.A1(n_3702),
.A2(n_3669),
.B1(n_3636),
.B2(n_3538),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_SL g5259 ( 
.A(n_3317),
.B(n_3327),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_3572),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_3294),
.B(n_3298),
.Y(n_5261)
);

AND2x4_ASAP7_75t_L g5262 ( 
.A(n_3271),
.B(n_3614),
.Y(n_5262)
);

HB1xp67_ASAP7_75t_L g5263 ( 
.A(n_3539),
.Y(n_5263)
);

BUFx3_ASAP7_75t_L g5264 ( 
.A(n_3638),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_3572),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_3592),
.Y(n_5266)
);

BUFx3_ASAP7_75t_L g5267 ( 
.A(n_3638),
.Y(n_5267)
);

BUFx6f_ASAP7_75t_L g5268 ( 
.A(n_3346),
.Y(n_5268)
);

NOR2xp33_ASAP7_75t_SL g5269 ( 
.A(n_3306),
.B(n_4145),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_3300),
.B(n_3323),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_3592),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_3300),
.B(n_3323),
.Y(n_5272)
);

AOI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_4100),
.A2(n_4107),
.B(n_4101),
.Y(n_5273)
);

AOI22xp5_ASAP7_75t_L g5274 ( 
.A1(n_3440),
.A2(n_3606),
.B1(n_3648),
.B2(n_3342),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_3621),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_3336),
.B(n_3342),
.Y(n_5276)
);

CKINVDCx16_ASAP7_75t_R g5277 ( 
.A(n_3648),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_3336),
.B(n_3352),
.Y(n_5278)
);

BUFx3_ASAP7_75t_L g5279 ( 
.A(n_3638),
.Y(n_5279)
);

NAND2xp33_ASAP7_75t_SL g5280 ( 
.A(n_3352),
.B(n_3354),
.Y(n_5280)
);

NOR2x1p5_ASAP7_75t_L g5281 ( 
.A(n_3657),
.B(n_3658),
.Y(n_5281)
);

INVx3_ASAP7_75t_L g5282 ( 
.A(n_3865),
.Y(n_5282)
);

OR2x2_ASAP7_75t_L g5283 ( 
.A(n_3341),
.B(n_3440),
.Y(n_5283)
);

NAND2xp5_ASAP7_75t_L g5284 ( 
.A(n_3354),
.B(n_3374),
.Y(n_5284)
);

HB1xp67_ASAP7_75t_L g5285 ( 
.A(n_3732),
.Y(n_5285)
);

OR2x6_ASAP7_75t_L g5286 ( 
.A(n_4101),
.B(n_4107),
.Y(n_5286)
);

INVx4_ASAP7_75t_L g5287 ( 
.A(n_3865),
.Y(n_5287)
);

INVx3_ASAP7_75t_L g5288 ( 
.A(n_3865),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_3621),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_4110),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_3616),
.B(n_3624),
.Y(n_5291)
);

AOI22xp33_ASAP7_75t_L g5292 ( 
.A1(n_3374),
.A2(n_3384),
.B1(n_3385),
.B2(n_3377),
.Y(n_5292)
);

BUFx3_ASAP7_75t_L g5293 ( 
.A(n_3638),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_4110),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4111),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4111),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_4197),
.Y(n_5297)
);

BUFx2_ASAP7_75t_L g5298 ( 
.A(n_3739),
.Y(n_5298)
);

BUFx3_ASAP7_75t_L g5299 ( 
.A(n_3638),
.Y(n_5299)
);

AND2x2_ASAP7_75t_L g5300 ( 
.A(n_3616),
.B(n_3624),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_3377),
.B(n_3384),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_3385),
.B(n_3398),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_4197),
.Y(n_5303)
);

AND2x2_ASAP7_75t_L g5304 ( 
.A(n_3616),
.B(n_3624),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4198),
.Y(n_5305)
);

CKINVDCx20_ASAP7_75t_R g5306 ( 
.A(n_3707),
.Y(n_5306)
);

AND2x4_ASAP7_75t_L g5307 ( 
.A(n_3079),
.B(n_3088),
.Y(n_5307)
);

OR2x6_ASAP7_75t_L g5308 ( 
.A(n_4198),
.B(n_4201),
.Y(n_5308)
);

OR2x2_ASAP7_75t_L g5309 ( 
.A(n_3456),
.B(n_4201),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_SL g5310 ( 
.A(n_3328),
.B(n_3332),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4208),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_3398),
.B(n_3400),
.Y(n_5312)
);

AOI21xp33_ASAP7_75t_L g5313 ( 
.A1(n_3489),
.A2(n_3491),
.B(n_3547),
.Y(n_5313)
);

BUFx6f_ASAP7_75t_L g5314 ( 
.A(n_3346),
.Y(n_5314)
);

BUFx2_ASAP7_75t_L g5315 ( 
.A(n_3973),
.Y(n_5315)
);

OR2x2_ASAP7_75t_SL g5316 ( 
.A(n_3669),
.B(n_3647),
.Y(n_5316)
);

OR2x6_ASAP7_75t_L g5317 ( 
.A(n_4208),
.B(n_4211),
.Y(n_5317)
);

OR2x6_ASAP7_75t_L g5318 ( 
.A(n_4211),
.B(n_4215),
.Y(n_5318)
);

NAND2xp5_ASAP7_75t_L g5319 ( 
.A(n_3400),
.B(n_3407),
.Y(n_5319)
);

NAND2xp5_ASAP7_75t_L g5320 ( 
.A(n_3407),
.B(n_3413),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4215),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_L g5322 ( 
.A(n_3413),
.B(n_3427),
.Y(n_5322)
);

INVx3_ASAP7_75t_L g5323 ( 
.A(n_3958),
.Y(n_5323)
);

AND3x2_ASAP7_75t_SL g5324 ( 
.A(n_3633),
.B(n_3685),
.C(n_3674),
.Y(n_5324)
);

AND2x2_ASAP7_75t_L g5325 ( 
.A(n_3533),
.B(n_3079),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_4219),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4219),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_3427),
.B(n_3431),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_3431),
.B(n_3436),
.Y(n_5329)
);

BUFx8_ASAP7_75t_L g5330 ( 
.A(n_3669),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_3436),
.B(n_3331),
.Y(n_5331)
);

HB1xp67_ASAP7_75t_L g5332 ( 
.A(n_4000),
.Y(n_5332)
);

INVx2_ASAP7_75t_SL g5333 ( 
.A(n_3958),
.Y(n_5333)
);

AOI22xp33_ASAP7_75t_L g5334 ( 
.A1(n_3439),
.A2(n_3456),
.B1(n_3366),
.B2(n_3373),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_3489),
.B(n_3494),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_3333),
.B(n_3337),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4220),
.Y(n_5337)
);

OR2x6_ASAP7_75t_L g5338 ( 
.A(n_4220),
.B(n_4261),
.Y(n_5338)
);

AOI22x1_ASAP7_75t_L g5339 ( 
.A1(n_3860),
.A2(n_3861),
.B1(n_3868),
.B2(n_3862),
.Y(n_5339)
);

NOR2x1_ASAP7_75t_L g5340 ( 
.A(n_3232),
.B(n_3330),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_4261),
.Y(n_5341)
);

INVxp67_ASAP7_75t_SL g5342 ( 
.A(n_4268),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_SL g5343 ( 
.A(n_3338),
.B(n_3353),
.Y(n_5343)
);

NOR2xp33_ASAP7_75t_L g5344 ( 
.A(n_3433),
.B(n_3831),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_3230),
.B(n_3237),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_L g5346 ( 
.A(n_3497),
.B(n_3450),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4268),
.Y(n_5347)
);

INVx6_ASAP7_75t_L g5348 ( 
.A(n_3958),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_L g5349 ( 
.A(n_3450),
.B(n_3585),
.Y(n_5349)
);

INVx2_ASAP7_75t_SL g5350 ( 
.A(n_3958),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_3555),
.B(n_3582),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_3609),
.B(n_3446),
.Y(n_5352)
);

INVx3_ASAP7_75t_L g5353 ( 
.A(n_3975),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4388),
.Y(n_5354)
);

OR2x2_ASAP7_75t_L g5355 ( 
.A(n_4388),
.B(n_4393),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_3512),
.B(n_3514),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_4393),
.Y(n_5357)
);

OAI21x1_ASAP7_75t_L g5358 ( 
.A1(n_3100),
.A2(n_4410),
.B(n_4409),
.Y(n_5358)
);

NAND2x1p5_ASAP7_75t_L g5359 ( 
.A(n_3869),
.B(n_3872),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_3512),
.B(n_3533),
.Y(n_5360)
);

BUFx2_ASAP7_75t_L g5361 ( 
.A(n_4037),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4409),
.Y(n_5362)
);

INVx4_ASAP7_75t_L g5363 ( 
.A(n_3975),
.Y(n_5363)
);

NOR2xp67_ASAP7_75t_L g5364 ( 
.A(n_3504),
.B(n_3505),
.Y(n_5364)
);

INVx3_ASAP7_75t_SL g5365 ( 
.A(n_3975),
.Y(n_5365)
);

AOI22xp33_ASAP7_75t_L g5366 ( 
.A1(n_3363),
.A2(n_3373),
.B1(n_3389),
.B2(n_3366),
.Y(n_5366)
);

OR2x4_ASAP7_75t_L g5367 ( 
.A(n_3669),
.B(n_3647),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_3459),
.B(n_3478),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_SL g5369 ( 
.A(n_3600),
.B(n_3132),
.Y(n_5369)
);

AOI22xp5_ASAP7_75t_L g5370 ( 
.A1(n_3606),
.A2(n_3535),
.B1(n_3659),
.B2(n_3603),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_4410),
.Y(n_5371)
);

BUFx3_ASAP7_75t_L g5372 ( 
.A(n_4402),
.Y(n_5372)
);

NOR2xp33_ASAP7_75t_L g5373 ( 
.A(n_3960),
.B(n_4020),
.Y(n_5373)
);

BUFx2_ASAP7_75t_L g5374 ( 
.A(n_4082),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_3459),
.B(n_3478),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_3532),
.B(n_3546),
.Y(n_5376)
);

CKINVDCx20_ASAP7_75t_R g5377 ( 
.A(n_4402),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_3532),
.B(n_3546),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_4411),
.Y(n_5379)
);

NOR2x1_ASAP7_75t_R g5380 ( 
.A(n_3310),
.B(n_3324),
.Y(n_5380)
);

HB1xp67_ASAP7_75t_L g5381 ( 
.A(n_4094),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_L g5382 ( 
.A(n_3521),
.B(n_3527),
.Y(n_5382)
);

NOR2xp33_ASAP7_75t_L g5383 ( 
.A(n_4056),
.B(n_4130),
.Y(n_5383)
);

AOI22xp33_ASAP7_75t_L g5384 ( 
.A1(n_3363),
.A2(n_3423),
.B1(n_3435),
.B2(n_3389),
.Y(n_5384)
);

INVx1_ASAP7_75t_SL g5385 ( 
.A(n_3509),
.Y(n_5385)
);

INVx6_ASAP7_75t_L g5386 ( 
.A(n_3975),
.Y(n_5386)
);

AND3x1_ASAP7_75t_L g5387 ( 
.A(n_3652),
.B(n_3646),
.C(n_3451),
.Y(n_5387)
);

NAND2xp33_ASAP7_75t_SL g5388 ( 
.A(n_3706),
.B(n_3669),
.Y(n_5388)
);

CKINVDCx11_ASAP7_75t_R g5389 ( 
.A(n_3324),
.Y(n_5389)
);

INVx3_ASAP7_75t_L g5390 ( 
.A(n_4009),
.Y(n_5390)
);

HB1xp67_ASAP7_75t_L g5391 ( 
.A(n_4236),
.Y(n_5391)
);

NAND2xp5_ASAP7_75t_L g5392 ( 
.A(n_3529),
.B(n_3536),
.Y(n_5392)
);

INVx5_ASAP7_75t_L g5393 ( 
.A(n_4414),
.Y(n_5393)
);

HB1xp67_ASAP7_75t_L g5394 ( 
.A(n_4294),
.Y(n_5394)
);

BUFx4f_ASAP7_75t_L g5395 ( 
.A(n_4414),
.Y(n_5395)
);

BUFx2_ASAP7_75t_L g5396 ( 
.A(n_4302),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_4411),
.Y(n_5397)
);

AND2x6_ASAP7_75t_L g5398 ( 
.A(n_3607),
.B(n_3620),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_3347),
.Y(n_5399)
);

INVx4_ASAP7_75t_L g5400 ( 
.A(n_4009),
.Y(n_5400)
);

OR2x6_ASAP7_75t_L g5401 ( 
.A(n_3100),
.B(n_3879),
.Y(n_5401)
);

OAI22xp5_ASAP7_75t_L g5402 ( 
.A1(n_4259),
.A2(n_4391),
.B1(n_3470),
.B2(n_3518),
.Y(n_5402)
);

INVx3_ASAP7_75t_L g5403 ( 
.A(n_4009),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_SL g5404 ( 
.A(n_3581),
.B(n_3659),
.Y(n_5404)
);

BUFx2_ASAP7_75t_L g5405 ( 
.A(n_4406),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_L g5406 ( 
.A(n_3506),
.B(n_3507),
.Y(n_5406)
);

HB1xp67_ASAP7_75t_L g5407 ( 
.A(n_3347),
.Y(n_5407)
);

AOI221x1_ASAP7_75t_L g5408 ( 
.A1(n_3887),
.A2(n_3908),
.B1(n_3911),
.B2(n_3907),
.C(n_3891),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_3923),
.Y(n_5409)
);

BUFx3_ASAP7_75t_L g5410 ( 
.A(n_4402),
.Y(n_5410)
);

INVx3_ASAP7_75t_L g5411 ( 
.A(n_4009),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_L g5412 ( 
.A(n_3508),
.B(n_3513),
.Y(n_5412)
);

BUFx4f_ASAP7_75t_L g5413 ( 
.A(n_4414),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_3453),
.B(n_3457),
.Y(n_5414)
);

CKINVDCx5p33_ASAP7_75t_R g5415 ( 
.A(n_3324),
.Y(n_5415)
);

NAND2xp5_ASAP7_75t_L g5416 ( 
.A(n_3453),
.B(n_3457),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_SL g5417 ( 
.A(n_3666),
.B(n_3232),
.Y(n_5417)
);

INVxp67_ASAP7_75t_L g5418 ( 
.A(n_3629),
.Y(n_5418)
);

NOR2xp67_ASAP7_75t_L g5419 ( 
.A(n_4046),
.B(n_4102),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_3462),
.B(n_3463),
.Y(n_5420)
);

BUFx3_ASAP7_75t_L g5421 ( 
.A(n_3654),
.Y(n_5421)
);

AO22x1_ASAP7_75t_L g5422 ( 
.A1(n_3615),
.A2(n_3451),
.B1(n_4102),
.B2(n_4046),
.Y(n_5422)
);

NOR2xp33_ASAP7_75t_L g5423 ( 
.A(n_3490),
.B(n_3461),
.Y(n_5423)
);

CKINVDCx11_ASAP7_75t_R g5424 ( 
.A(n_3215),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_3628),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_3931),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_3943),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_3462),
.B(n_3463),
.Y(n_5428)
);

INVx3_ASAP7_75t_L g5429 ( 
.A(n_4046),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_3945),
.Y(n_5430)
);

BUFx8_ASAP7_75t_L g5431 ( 
.A(n_3635),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_L g5432 ( 
.A(n_3509),
.B(n_4058),
.Y(n_5432)
);

HB1xp67_ASAP7_75t_L g5433 ( 
.A(n_3537),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_SL g5434 ( 
.A(n_3666),
.B(n_3330),
.Y(n_5434)
);

AOI22xp5_ASAP7_75t_L g5435 ( 
.A1(n_3603),
.A2(n_3567),
.B1(n_3435),
.B2(n_3452),
.Y(n_5435)
);

NOR2xp33_ASAP7_75t_L g5436 ( 
.A(n_4058),
.B(n_4080),
.Y(n_5436)
);

AOI22x1_ASAP7_75t_L g5437 ( 
.A1(n_3946),
.A2(n_3955),
.B1(n_3964),
.B2(n_3959),
.Y(n_5437)
);

NOR2xp67_ASAP7_75t_L g5438 ( 
.A(n_4046),
.B(n_4102),
.Y(n_5438)
);

NAND2xp5_ASAP7_75t_SL g5439 ( 
.A(n_3543),
.B(n_3545),
.Y(n_5439)
);

BUFx2_ASAP7_75t_L g5440 ( 
.A(n_3644),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_3464),
.B(n_3465),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_L g5442 ( 
.A(n_3464),
.B(n_3465),
.Y(n_5442)
);

INVx3_ASAP7_75t_L g5443 ( 
.A(n_4102),
.Y(n_5443)
);

AOI22xp33_ASAP7_75t_L g5444 ( 
.A1(n_3423),
.A2(n_3452),
.B1(n_3646),
.B2(n_3469),
.Y(n_5444)
);

NOR2xp33_ASAP7_75t_L g5445 ( 
.A(n_4080),
.B(n_3579),
.Y(n_5445)
);

BUFx4f_ASAP7_75t_L g5446 ( 
.A(n_3409),
.Y(n_5446)
);

OAI22xp5_ASAP7_75t_SL g5447 ( 
.A1(n_3241),
.A2(n_3301),
.B1(n_3884),
.B2(n_3286),
.Y(n_5447)
);

INVxp67_ASAP7_75t_L g5448 ( 
.A(n_3445),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_3475),
.B(n_3476),
.Y(n_5449)
);

CKINVDCx20_ASAP7_75t_R g5450 ( 
.A(n_3215),
.Y(n_5450)
);

AOI221xp5_ASAP7_75t_SL g5451 ( 
.A1(n_3593),
.A2(n_3562),
.B1(n_3503),
.B2(n_3445),
.C(n_3485),
.Y(n_5451)
);

INVx3_ASAP7_75t_L g5452 ( 
.A(n_4104),
.Y(n_5452)
);

BUFx6f_ASAP7_75t_L g5453 ( 
.A(n_4104),
.Y(n_5453)
);

NOR2xp33_ASAP7_75t_L g5454 ( 
.A(n_3619),
.B(n_3558),
.Y(n_5454)
);

A2O1A1Ixp33_ASAP7_75t_L g5455 ( 
.A1(n_3968),
.A2(n_3974),
.B(n_3988),
.C(n_3983),
.Y(n_5455)
);

BUFx3_ASAP7_75t_L g5456 ( 
.A(n_3654),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_L g5457 ( 
.A(n_3475),
.B(n_3476),
.Y(n_5457)
);

BUFx2_ASAP7_75t_L g5458 ( 
.A(n_3615),
.Y(n_5458)
);

BUFx6f_ASAP7_75t_L g5459 ( 
.A(n_4104),
.Y(n_5459)
);

NAND2xp5_ASAP7_75t_L g5460 ( 
.A(n_3477),
.B(n_3480),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_3993),
.Y(n_5461)
);

INVx3_ASAP7_75t_L g5462 ( 
.A(n_4104),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_3477),
.B(n_3480),
.Y(n_5463)
);

BUFx2_ASAP7_75t_L g5464 ( 
.A(n_3654),
.Y(n_5464)
);

INVx2_ASAP7_75t_SL g5465 ( 
.A(n_4154),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_4011),
.Y(n_5466)
);

CKINVDCx16_ASAP7_75t_R g5467 ( 
.A(n_4038),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_4014),
.Y(n_5468)
);

NOR2xp33_ASAP7_75t_L g5469 ( 
.A(n_3625),
.B(n_3639),
.Y(n_5469)
);

AND2x4_ASAP7_75t_SL g5470 ( 
.A(n_4154),
.B(n_4162),
.Y(n_5470)
);

BUFx2_ASAP7_75t_L g5471 ( 
.A(n_3654),
.Y(n_5471)
);

INVx3_ASAP7_75t_L g5472 ( 
.A(n_4154),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_3625),
.B(n_3632),
.Y(n_5473)
);

BUFx2_ASAP7_75t_L g5474 ( 
.A(n_4154),
.Y(n_5474)
);

BUFx2_ASAP7_75t_L g5475 ( 
.A(n_4162),
.Y(n_5475)
);

INVxp33_ASAP7_75t_SL g5476 ( 
.A(n_3233),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_3501),
.B(n_3502),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_SL g5478 ( 
.A(n_3601),
.B(n_3575),
.Y(n_5478)
);

AOI22xp5_ASAP7_75t_L g5479 ( 
.A1(n_3646),
.A2(n_3597),
.B1(n_3652),
.B2(n_3460),
.Y(n_5479)
);

NAND2xp5_ASAP7_75t_L g5480 ( 
.A(n_3501),
.B(n_3502),
.Y(n_5480)
);

INVx3_ASAP7_75t_L g5481 ( 
.A(n_4162),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_4016),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_3516),
.B(n_3517),
.Y(n_5483)
);

BUFx6f_ASAP7_75t_L g5484 ( 
.A(n_4162),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_SL g5485 ( 
.A(n_3576),
.B(n_3662),
.Y(n_5485)
);

CKINVDCx5p33_ASAP7_75t_R g5486 ( 
.A(n_3215),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_4021),
.Y(n_5487)
);

NOR2xp33_ASAP7_75t_R g5488 ( 
.A(n_3694),
.B(n_4176),
.Y(n_5488)
);

BUFx6f_ASAP7_75t_L g5489 ( 
.A(n_4193),
.Y(n_5489)
);

INVx2_ASAP7_75t_SL g5490 ( 
.A(n_4193),
.Y(n_5490)
);

NOR2xp33_ASAP7_75t_L g5491 ( 
.A(n_3608),
.B(n_3602),
.Y(n_5491)
);

BUFx2_ASAP7_75t_L g5492 ( 
.A(n_4193),
.Y(n_5492)
);

HB1xp67_ASAP7_75t_L g5493 ( 
.A(n_3454),
.Y(n_5493)
);

BUFx3_ASAP7_75t_L g5494 ( 
.A(n_3641),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_4023),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_3516),
.B(n_3517),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_3519),
.B(n_3528),
.Y(n_5497)
);

BUFx2_ASAP7_75t_SL g5498 ( 
.A(n_3185),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_3519),
.B(n_3528),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_3577),
.B(n_3578),
.Y(n_5500)
);

INVx3_ASAP7_75t_L g5501 ( 
.A(n_4193),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_3577),
.B(n_3578),
.Y(n_5502)
);

OR2x6_ASAP7_75t_L g5503 ( 
.A(n_4026),
.B(n_4030),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_3584),
.B(n_3587),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_3584),
.B(n_3587),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_4032),
.Y(n_5506)
);

AOI22xp33_ASAP7_75t_L g5507 ( 
.A1(n_3646),
.A2(n_3597),
.B1(n_3641),
.B2(n_3460),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_4040),
.Y(n_5508)
);

INVx1_ASAP7_75t_SL g5509 ( 
.A(n_3580),
.Y(n_5509)
);

HB1xp67_ASAP7_75t_L g5510 ( 
.A(n_3454),
.Y(n_5510)
);

AOI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_3597),
.A2(n_3493),
.B1(n_3496),
.B2(n_3485),
.Y(n_5511)
);

NOR2xp33_ASAP7_75t_L g5512 ( 
.A(n_3597),
.B(n_3590),
.Y(n_5512)
);

AND3x1_ASAP7_75t_SL g5513 ( 
.A(n_3712),
.B(n_3649),
.C(n_3645),
.Y(n_5513)
);

BUFx2_ASAP7_75t_L g5514 ( 
.A(n_3607),
.Y(n_5514)
);

NOR3xp33_ASAP7_75t_L g5515 ( 
.A(n_4041),
.B(n_4061),
.C(n_4045),
.Y(n_5515)
);

NOR2xp33_ASAP7_75t_L g5516 ( 
.A(n_3590),
.B(n_3700),
.Y(n_5516)
);

BUFx3_ASAP7_75t_L g5517 ( 
.A(n_3416),
.Y(n_5517)
);

OR2x6_ASAP7_75t_L g5518 ( 
.A(n_4069),
.B(n_4074),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_4076),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_L g5520 ( 
.A(n_3589),
.B(n_3595),
.Y(n_5520)
);

INVx1_ASAP7_75t_SL g5521 ( 
.A(n_3580),
.Y(n_5521)
);

NOR2xp33_ASAP7_75t_R g5522 ( 
.A(n_3694),
.B(n_4234),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_L g5523 ( 
.A(n_3589),
.B(n_3595),
.Y(n_5523)
);

XOR2xp5_ASAP7_75t_L g5524 ( 
.A(n_4277),
.B(n_3590),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_L g5525 ( 
.A(n_3598),
.B(n_3599),
.Y(n_5525)
);

NOR2xp33_ASAP7_75t_SL g5526 ( 
.A(n_3680),
.B(n_3692),
.Y(n_5526)
);

NOR2xp33_ASAP7_75t_R g5527 ( 
.A(n_3657),
.B(n_3658),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_SL g5528 ( 
.A(n_3662),
.B(n_3574),
.Y(n_5528)
);

BUFx3_ASAP7_75t_L g5529 ( 
.A(n_3416),
.Y(n_5529)
);

AOI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_3493),
.A2(n_3515),
.B1(n_3496),
.B2(n_3635),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_4732),
.Y(n_5531)
);

O2A1O1Ixp5_ASAP7_75t_L g5532 ( 
.A1(n_4502),
.A2(n_4366),
.B(n_4361),
.C(n_4360),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_4732),
.Y(n_5533)
);

O2A1O1Ixp33_ASAP7_75t_L g5534 ( 
.A1(n_4777),
.A2(n_3559),
.B(n_3561),
.C(n_3515),
.Y(n_5534)
);

BUFx3_ASAP7_75t_L g5535 ( 
.A(n_5159),
.Y(n_5535)
);

NOR2xp33_ASAP7_75t_L g5536 ( 
.A(n_4492),
.B(n_3617),
.Y(n_5536)
);

AOI22xp33_ASAP7_75t_L g5537 ( 
.A1(n_4484),
.A2(n_3618),
.B1(n_3640),
.B2(n_3623),
.Y(n_5537)
);

NOR2xp67_ASAP7_75t_L g5538 ( 
.A(n_5093),
.B(n_4125),
.Y(n_5538)
);

OAI22xp5_ASAP7_75t_L g5539 ( 
.A1(n_4452),
.A2(n_3596),
.B1(n_3598),
.B2(n_3599),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_4732),
.Y(n_5540)
);

INVx4_ASAP7_75t_L g5541 ( 
.A(n_4697),
.Y(n_5541)
);

OAI22xp5_ASAP7_75t_L g5542 ( 
.A1(n_4452),
.A2(n_4570),
.B1(n_4484),
.B2(n_4507),
.Y(n_5542)
);

NOR2xp33_ASAP7_75t_L g5543 ( 
.A(n_4492),
.B(n_3700),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_4737),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_SL g5545 ( 
.A(n_4507),
.B(n_4138),
.Y(n_5545)
);

INVx2_ASAP7_75t_L g5546 ( 
.A(n_4916),
.Y(n_5546)
);

AND2x6_ASAP7_75t_L g5547 ( 
.A(n_5206),
.B(n_3620),
.Y(n_5547)
);

INVx2_ASAP7_75t_SL g5548 ( 
.A(n_5517),
.Y(n_5548)
);

OAI22xp5_ASAP7_75t_SL g5549 ( 
.A1(n_4543),
.A2(n_3668),
.B1(n_3693),
.B2(n_3926),
.Y(n_5549)
);

AND2x4_ASAP7_75t_L g5550 ( 
.A(n_4519),
.B(n_4141),
.Y(n_5550)
);

INVx2_ASAP7_75t_L g5551 ( 
.A(n_4916),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_4737),
.Y(n_5552)
);

INVx4_ASAP7_75t_L g5553 ( 
.A(n_4697),
.Y(n_5553)
);

INVx2_ASAP7_75t_SL g5554 ( 
.A(n_5517),
.Y(n_5554)
);

AOI21x1_ASAP7_75t_L g5555 ( 
.A1(n_5369),
.A2(n_4164),
.B(n_4142),
.Y(n_5555)
);

BUFx3_ASAP7_75t_L g5556 ( 
.A(n_5159),
.Y(n_5556)
);

BUFx8_ASAP7_75t_L g5557 ( 
.A(n_4775),
.Y(n_5557)
);

NOR2xp33_ASAP7_75t_L g5558 ( 
.A(n_4555),
.B(n_3680),
.Y(n_5558)
);

AOI21xp5_ASAP7_75t_L g5559 ( 
.A1(n_5139),
.A2(n_4170),
.B(n_4168),
.Y(n_5559)
);

INVx2_ASAP7_75t_L g5560 ( 
.A(n_4916),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_4916),
.Y(n_5561)
);

AOI21xp5_ASAP7_75t_L g5562 ( 
.A1(n_5139),
.A2(n_4179),
.B(n_4173),
.Y(n_5562)
);

BUFx3_ASAP7_75t_L g5563 ( 
.A(n_5159),
.Y(n_5563)
);

INVx4_ASAP7_75t_L g5564 ( 
.A(n_4697),
.Y(n_5564)
);

AOI21xp5_ASAP7_75t_L g5565 ( 
.A1(n_5191),
.A2(n_4185),
.B(n_4183),
.Y(n_5565)
);

BUFx6f_ASAP7_75t_L g5566 ( 
.A(n_4478),
.Y(n_5566)
);

A2O1A1Ixp33_ASAP7_75t_L g5567 ( 
.A1(n_4436),
.A2(n_4311),
.B(n_4299),
.C(n_4291),
.Y(n_5567)
);

INVx1_ASAP7_75t_SL g5568 ( 
.A(n_5043),
.Y(n_5568)
);

O2A1O1Ixp33_ASAP7_75t_L g5569 ( 
.A1(n_4777),
.A2(n_3667),
.B(n_3655),
.C(n_3570),
.Y(n_5569)
);

AOI21xp5_ASAP7_75t_L g5570 ( 
.A1(n_5191),
.A2(n_4188),
.B(n_4186),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_4418),
.Y(n_5571)
);

AOI22xp33_ASAP7_75t_L g5572 ( 
.A1(n_4570),
.A2(n_3643),
.B1(n_3630),
.B2(n_3596),
.Y(n_5572)
);

NOR2xp33_ASAP7_75t_L g5573 ( 
.A(n_4555),
.B(n_3708),
.Y(n_5573)
);

CKINVDCx8_ASAP7_75t_R g5574 ( 
.A(n_5467),
.Y(n_5574)
);

INVxp67_ASAP7_75t_SL g5575 ( 
.A(n_5054),
.Y(n_5575)
);

BUFx6f_ASAP7_75t_L g5576 ( 
.A(n_4478),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_4737),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_4738),
.Y(n_5578)
);

NOR2x1_ASAP7_75t_L g5579 ( 
.A(n_5165),
.B(n_4108),
.Y(n_5579)
);

HB1xp67_ASAP7_75t_L g5580 ( 
.A(n_5054),
.Y(n_5580)
);

A2O1A1Ixp33_ASAP7_75t_L g5581 ( 
.A1(n_4436),
.A2(n_4272),
.B(n_4385),
.C(n_4382),
.Y(n_5581)
);

O2A1O1Ixp33_ASAP7_75t_L g5582 ( 
.A1(n_4502),
.A2(n_3715),
.B(n_3714),
.C(n_4308),
.Y(n_5582)
);

BUFx2_ASAP7_75t_SL g5583 ( 
.A(n_5176),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_4738),
.Y(n_5584)
);

NAND2xp5_ASAP7_75t_L g5585 ( 
.A(n_5190),
.B(n_4223),
.Y(n_5585)
);

BUFx4f_ASAP7_75t_L g5586 ( 
.A(n_4973),
.Y(n_5586)
);

AOI21xp5_ASAP7_75t_L g5587 ( 
.A1(n_5392),
.A2(n_4233),
.B(n_4230),
.Y(n_5587)
);

INVx2_ASAP7_75t_SL g5588 ( 
.A(n_5529),
.Y(n_5588)
);

BUFx3_ASAP7_75t_L g5589 ( 
.A(n_5159),
.Y(n_5589)
);

HB1xp67_ASAP7_75t_L g5590 ( 
.A(n_5066),
.Y(n_5590)
);

INVx1_ASAP7_75t_SL g5591 ( 
.A(n_5043),
.Y(n_5591)
);

INVxp67_ASAP7_75t_L g5592 ( 
.A(n_5167),
.Y(n_5592)
);

BUFx12f_ASAP7_75t_L g5593 ( 
.A(n_5389),
.Y(n_5593)
);

BUFx6f_ASAP7_75t_L g5594 ( 
.A(n_4478),
.Y(n_5594)
);

AND2x4_ASAP7_75t_L g5595 ( 
.A(n_4519),
.B(n_4239),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_4418),
.Y(n_5596)
);

HB1xp67_ASAP7_75t_L g5597 ( 
.A(n_5066),
.Y(n_5597)
);

NAND2xp5_ASAP7_75t_SL g5598 ( 
.A(n_4582),
.B(n_4245),
.Y(n_5598)
);

O2A1O1Ixp33_ASAP7_75t_L g5599 ( 
.A1(n_4520),
.A2(n_3715),
.B(n_4343),
.C(n_4336),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_4738),
.Y(n_5600)
);

BUFx3_ASAP7_75t_L g5601 ( 
.A(n_5159),
.Y(n_5601)
);

AOI22xp33_ASAP7_75t_SL g5602 ( 
.A1(n_4439),
.A2(n_4108),
.B1(n_4376),
.B2(n_4374),
.Y(n_5602)
);

CKINVDCx5p33_ASAP7_75t_R g5603 ( 
.A(n_4429),
.Y(n_5603)
);

INVx2_ASAP7_75t_L g5604 ( 
.A(n_4418),
.Y(n_5604)
);

NAND2xp5_ASAP7_75t_SL g5605 ( 
.A(n_4582),
.B(n_4254),
.Y(n_5605)
);

AND2x4_ASAP7_75t_L g5606 ( 
.A(n_4519),
.B(n_4269),
.Y(n_5606)
);

NAND2x1p5_ASAP7_75t_L g5607 ( 
.A(n_4697),
.B(n_4276),
.Y(n_5607)
);

AOI21xp5_ASAP7_75t_L g5608 ( 
.A1(n_5382),
.A2(n_4352),
.B(n_4371),
.Y(n_5608)
);

AOI22xp5_ASAP7_75t_L g5609 ( 
.A1(n_4543),
.A2(n_3704),
.B1(n_3713),
.B2(n_3697),
.Y(n_5609)
);

INVx2_ASAP7_75t_SL g5610 ( 
.A(n_5281),
.Y(n_5610)
);

O2A1O1Ixp33_ASAP7_75t_L g5611 ( 
.A1(n_4520),
.A2(n_4334),
.B(n_4331),
.C(n_4323),
.Y(n_5611)
);

AOI21xp33_ASAP7_75t_L g5612 ( 
.A1(n_4431),
.A2(n_4616),
.B(n_4511),
.Y(n_5612)
);

AOI22xp33_ASAP7_75t_L g5613 ( 
.A1(n_4610),
.A2(n_3704),
.B1(n_4367),
.B2(n_4359),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_4744),
.Y(n_5614)
);

OA21x2_ASAP7_75t_L g5615 ( 
.A1(n_5408),
.A2(n_5358),
.B(n_4606),
.Y(n_5615)
);

O2A1O1Ixp5_ASAP7_75t_L g5616 ( 
.A1(n_4713),
.A2(n_4806),
.B(n_5088),
.C(n_4561),
.Y(n_5616)
);

A2O1A1Ixp33_ASAP7_75t_SL g5617 ( 
.A1(n_4713),
.A2(n_3627),
.B(n_3686),
.C(n_3693),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_4541),
.B(n_4344),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_4744),
.Y(n_5619)
);

INVx1_ASAP7_75t_SL g5620 ( 
.A(n_5163),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_5382),
.A2(n_4354),
.B(n_3564),
.Y(n_5621)
);

O2A1O1Ixp33_ASAP7_75t_L g5622 ( 
.A1(n_4580),
.A2(n_3706),
.B(n_3686),
.C(n_3678),
.Y(n_5622)
);

BUFx6f_ASAP7_75t_L g5623 ( 
.A(n_4478),
.Y(n_5623)
);

AOI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_4610),
.A2(n_3713),
.B1(n_3697),
.B2(n_3557),
.Y(n_5624)
);

INVx2_ASAP7_75t_L g5625 ( 
.A(n_4418),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5093),
.B(n_4119),
.Y(n_5626)
);

AOI22xp33_ASAP7_75t_SL g5627 ( 
.A1(n_4439),
.A2(n_3149),
.B1(n_4320),
.B2(n_3807),
.Y(n_5627)
);

INVx2_ASAP7_75t_SL g5628 ( 
.A(n_5281),
.Y(n_5628)
);

AOI22xp5_ASAP7_75t_L g5629 ( 
.A1(n_4443),
.A2(n_3713),
.B1(n_3697),
.B2(n_3557),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5152),
.B(n_4119),
.Y(n_5630)
);

BUFx2_ASAP7_75t_SL g5631 ( 
.A(n_5176),
.Y(n_5631)
);

BUFx12f_ASAP7_75t_L g5632 ( 
.A(n_5389),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_4423),
.Y(n_5633)
);

OAI22xp5_ASAP7_75t_SL g5634 ( 
.A1(n_4742),
.A2(n_4390),
.B1(n_4035),
.B2(n_3926),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_4744),
.Y(n_5635)
);

INVxp67_ASAP7_75t_L g5636 ( 
.A(n_5167),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5152),
.B(n_4119),
.Y(n_5637)
);

INVx2_ASAP7_75t_L g5638 ( 
.A(n_4423),
.Y(n_5638)
);

AOI22xp33_ASAP7_75t_L g5639 ( 
.A1(n_4551),
.A2(n_3713),
.B1(n_3604),
.B2(n_3611),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_4888),
.B(n_4121),
.Y(n_5640)
);

INVx2_ASAP7_75t_L g5641 ( 
.A(n_4423),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_4888),
.B(n_4121),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_4746),
.Y(n_5643)
);

BUFx12f_ASAP7_75t_L g5644 ( 
.A(n_5424),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_SL g5645 ( 
.A(n_4695),
.B(n_3708),
.Y(n_5645)
);

A2O1A1Ixp33_ASAP7_75t_L g5646 ( 
.A1(n_5075),
.A2(n_3548),
.B(n_3381),
.C(n_4282),
.Y(n_5646)
);

OR2x6_ASAP7_75t_L g5647 ( 
.A(n_4478),
.B(n_3185),
.Y(n_5647)
);

CKINVDCx5p33_ASAP7_75t_R g5648 ( 
.A(n_4429),
.Y(n_5648)
);

INVx3_ASAP7_75t_SL g5649 ( 
.A(n_5217),
.Y(n_5649)
);

A2O1A1Ixp33_ASAP7_75t_L g5650 ( 
.A1(n_5075),
.A2(n_4826),
.B(n_4428),
.C(n_4451),
.Y(n_5650)
);

O2A1O1Ixp33_ASAP7_75t_L g5651 ( 
.A1(n_4580),
.A2(n_3626),
.B(n_3634),
.C(n_3703),
.Y(n_5651)
);

OR2x2_ASAP7_75t_L g5652 ( 
.A(n_4426),
.B(n_3685),
.Y(n_5652)
);

INVx2_ASAP7_75t_SL g5653 ( 
.A(n_5281),
.Y(n_5653)
);

OAI21xp5_ASAP7_75t_L g5654 ( 
.A1(n_4431),
.A2(n_3627),
.B(n_3495),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_L g5655 ( 
.A(n_4913),
.B(n_4121),
.Y(n_5655)
);

NAND2x1p5_ASAP7_75t_L g5656 ( 
.A(n_4697),
.B(n_3305),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4746),
.Y(n_5657)
);

OR2x2_ASAP7_75t_L g5658 ( 
.A(n_4426),
.B(n_3685),
.Y(n_5658)
);

O2A1O1Ixp33_ASAP7_75t_L g5659 ( 
.A1(n_4773),
.A2(n_3626),
.B(n_3634),
.C(n_3682),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_4746),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_5392),
.A2(n_3568),
.B(n_3566),
.Y(n_5661)
);

AOI22xp33_ASAP7_75t_L g5662 ( 
.A1(n_4551),
.A2(n_3710),
.B1(n_4320),
.B2(n_3807),
.Y(n_5662)
);

BUFx6f_ASAP7_75t_L g5663 ( 
.A(n_4478),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_4750),
.Y(n_5664)
);

CKINVDCx20_ASAP7_75t_R g5665 ( 
.A(n_4636),
.Y(n_5665)
);

NAND2xp5_ASAP7_75t_L g5666 ( 
.A(n_4913),
.B(n_5141),
.Y(n_5666)
);

NAND2xp5_ASAP7_75t_L g5667 ( 
.A(n_5141),
.B(n_4126),
.Y(n_5667)
);

AOI21xp5_ASAP7_75t_L g5668 ( 
.A1(n_4588),
.A2(n_3552),
.B(n_3565),
.Y(n_5668)
);

INVx1_ASAP7_75t_SL g5669 ( 
.A(n_5163),
.Y(n_5669)
);

BUFx8_ASAP7_75t_L g5670 ( 
.A(n_4775),
.Y(n_5670)
);

NOR2xp33_ASAP7_75t_L g5671 ( 
.A(n_5081),
.B(n_4826),
.Y(n_5671)
);

AOI21xp5_ASAP7_75t_L g5672 ( 
.A1(n_4588),
.A2(n_3560),
.B(n_3551),
.Y(n_5672)
);

INVxp67_ASAP7_75t_SL g5673 ( 
.A(n_5098),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_4750),
.Y(n_5674)
);

BUFx2_ASAP7_75t_L g5675 ( 
.A(n_4541),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_SL g5676 ( 
.A(n_4695),
.B(n_3633),
.Y(n_5676)
);

BUFx3_ASAP7_75t_L g5677 ( 
.A(n_5367),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_SL g5678 ( 
.A(n_4579),
.B(n_3633),
.Y(n_5678)
);

BUFx6f_ASAP7_75t_SL g5679 ( 
.A(n_4523),
.Y(n_5679)
);

INVx1_ASAP7_75t_SL g5680 ( 
.A(n_5385),
.Y(n_5680)
);

INVx4_ASAP7_75t_L g5681 ( 
.A(n_4697),
.Y(n_5681)
);

O2A1O1Ixp33_ASAP7_75t_L g5682 ( 
.A1(n_4773),
.A2(n_3672),
.B(n_3682),
.C(n_3679),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_4750),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_4752),
.Y(n_5684)
);

NAND2xp5_ASAP7_75t_SL g5685 ( 
.A(n_4579),
.B(n_3468),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_4812),
.B(n_4126),
.Y(n_5686)
);

INVx4_ASAP7_75t_L g5687 ( 
.A(n_4697),
.Y(n_5687)
);

BUFx6f_ASAP7_75t_L g5688 ( 
.A(n_4478),
.Y(n_5688)
);

NOR2xp33_ASAP7_75t_L g5689 ( 
.A(n_5081),
.B(n_3645),
.Y(n_5689)
);

NOR2xp33_ASAP7_75t_L g5690 ( 
.A(n_4495),
.B(n_3649),
.Y(n_5690)
);

O2A1O1Ixp33_ASAP7_75t_L g5691 ( 
.A1(n_4561),
.A2(n_3676),
.B(n_3665),
.C(n_3670),
.Y(n_5691)
);

A2O1A1Ixp33_ASAP7_75t_L g5692 ( 
.A1(n_4428),
.A2(n_3305),
.B(n_3381),
.C(n_4282),
.Y(n_5692)
);

AOI21xp5_ASAP7_75t_L g5693 ( 
.A1(n_4606),
.A2(n_3482),
.B(n_4114),
.Y(n_5693)
);

INVx4_ASAP7_75t_L g5694 ( 
.A(n_4697),
.Y(n_5694)
);

O2A1O1Ixp33_ASAP7_75t_L g5695 ( 
.A1(n_4573),
.A2(n_4590),
.B(n_4643),
.C(n_4613),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_4752),
.Y(n_5696)
);

INVx4_ASAP7_75t_L g5697 ( 
.A(n_4697),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_4752),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_L g5699 ( 
.A(n_4812),
.B(n_4126),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_L g5700 ( 
.A(n_4816),
.B(n_4922),
.Y(n_5700)
);

AOI21xp5_ASAP7_75t_L g5701 ( 
.A1(n_4731),
.A2(n_3305),
.B(n_3949),
.Y(n_5701)
);

BUFx6f_ASAP7_75t_L g5702 ( 
.A(n_4478),
.Y(n_5702)
);

A2O1A1Ixp33_ASAP7_75t_L g5703 ( 
.A1(n_4451),
.A2(n_3548),
.B(n_4114),
.C(n_3949),
.Y(n_5703)
);

INVx8_ASAP7_75t_L g5704 ( 
.A(n_4865),
.Y(n_5704)
);

OAI22xp5_ASAP7_75t_L g5705 ( 
.A1(n_4454),
.A2(n_3548),
.B1(n_3381),
.B2(n_4282),
.Y(n_5705)
);

HAxp5_ASAP7_75t_L g5706 ( 
.A(n_4449),
.B(n_3926),
.CON(n_5706),
.SN(n_5706)
);

AOI21xp5_ASAP7_75t_L g5707 ( 
.A1(n_4731),
.A2(n_3381),
.B(n_4114),
.Y(n_5707)
);

BUFx6f_ASAP7_75t_L g5708 ( 
.A(n_4478),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_4816),
.B(n_4126),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_4753),
.Y(n_5710)
);

AOI21xp5_ASAP7_75t_L g5711 ( 
.A1(n_4821),
.A2(n_3949),
.B(n_4282),
.Y(n_5711)
);

NOR2xp67_ASAP7_75t_L g5712 ( 
.A(n_5336),
.B(n_4175),
.Y(n_5712)
);

AOI21xp5_ASAP7_75t_L g5713 ( 
.A1(n_4821),
.A2(n_4114),
.B(n_3548),
.Y(n_5713)
);

O2A1O1Ixp33_ASAP7_75t_L g5714 ( 
.A1(n_4573),
.A2(n_3676),
.B(n_3679),
.C(n_3665),
.Y(n_5714)
);

OAI221xp5_ASAP7_75t_L g5715 ( 
.A1(n_4659),
.A2(n_3711),
.B1(n_3656),
.B2(n_3705),
.C(n_3673),
.Y(n_5715)
);

BUFx2_ASAP7_75t_L g5716 ( 
.A(n_4460),
.Y(n_5716)
);

AOI22xp33_ASAP7_75t_L g5717 ( 
.A1(n_4590),
.A2(n_3710),
.B1(n_4320),
.B2(n_3807),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_4753),
.Y(n_5718)
);

AND2x4_ASAP7_75t_L g5719 ( 
.A(n_4464),
.B(n_4175),
.Y(n_5719)
);

NAND2xp5_ASAP7_75t_SL g5720 ( 
.A(n_4585),
.B(n_3468),
.Y(n_5720)
);

INVx3_ASAP7_75t_L g5721 ( 
.A(n_4945),
.Y(n_5721)
);

AOI21xp5_ASAP7_75t_L g5722 ( 
.A1(n_4895),
.A2(n_3949),
.B(n_3305),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_4753),
.Y(n_5723)
);

NOR2xp67_ASAP7_75t_L g5724 ( 
.A(n_5336),
.B(n_5215),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_L g5725 ( 
.A(n_4922),
.B(n_4175),
.Y(n_5725)
);

NAND2xp5_ASAP7_75t_L g5726 ( 
.A(n_4935),
.B(n_4249),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_4756),
.Y(n_5727)
);

BUFx2_ASAP7_75t_L g5728 ( 
.A(n_4461),
.Y(n_5728)
);

BUFx2_ASAP7_75t_SL g5729 ( 
.A(n_5176),
.Y(n_5729)
);

INVx3_ASAP7_75t_L g5730 ( 
.A(n_4945),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_L g5731 ( 
.A(n_4935),
.B(n_4249),
.Y(n_5731)
);

NOR2xp33_ASAP7_75t_L g5732 ( 
.A(n_4495),
.B(n_3653),
.Y(n_5732)
);

AOI21x1_ASAP7_75t_L g5733 ( 
.A1(n_5369),
.A2(n_3285),
.B(n_3695),
.Y(n_5733)
);

AND2x2_ASAP7_75t_L g5734 ( 
.A(n_4464),
.B(n_4500),
.Y(n_5734)
);

INVx4_ASAP7_75t_L g5735 ( 
.A(n_5393),
.Y(n_5735)
);

NAND3xp33_ASAP7_75t_L g5736 ( 
.A(n_4585),
.B(n_3681),
.C(n_3663),
.Y(n_5736)
);

INVx1_ASAP7_75t_SL g5737 ( 
.A(n_5385),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_4756),
.Y(n_5738)
);

AND2x4_ASAP7_75t_L g5739 ( 
.A(n_4464),
.B(n_4295),
.Y(n_5739)
);

INVx1_ASAP7_75t_SL g5740 ( 
.A(n_4480),
.Y(n_5740)
);

OAI22xp5_ASAP7_75t_SL g5741 ( 
.A1(n_4742),
.A2(n_4390),
.B1(n_4035),
.B2(n_3149),
.Y(n_5741)
);

AND2x4_ASAP7_75t_L g5742 ( 
.A(n_4464),
.B(n_4295),
.Y(n_5742)
);

AOI222xp33_ASAP7_75t_L g5743 ( 
.A1(n_4443),
.A2(n_3594),
.B1(n_4035),
.B2(n_4390),
.C1(n_3697),
.C2(n_3718),
.Y(n_5743)
);

CKINVDCx5p33_ASAP7_75t_R g5744 ( 
.A(n_4456),
.Y(n_5744)
);

NAND2xp5_ASAP7_75t_SL g5745 ( 
.A(n_5137),
.B(n_3468),
.Y(n_5745)
);

AND2x4_ASAP7_75t_L g5746 ( 
.A(n_4500),
.B(n_4295),
.Y(n_5746)
);

OR2x6_ASAP7_75t_L g5747 ( 
.A(n_4504),
.B(n_3285),
.Y(n_5747)
);

AOI21xp5_ASAP7_75t_L g5748 ( 
.A1(n_4895),
.A2(n_3409),
.B(n_3468),
.Y(n_5748)
);

AOI222xp33_ASAP7_75t_L g5749 ( 
.A1(n_4443),
.A2(n_3718),
.B1(n_3753),
.B2(n_3149),
.C1(n_3296),
.C2(n_3335),
.Y(n_5749)
);

NAND2xp5_ASAP7_75t_L g5750 ( 
.A(n_4999),
.B(n_4295),
.Y(n_5750)
);

AOI21xp5_ASAP7_75t_L g5751 ( 
.A1(n_4897),
.A2(n_3409),
.B(n_3553),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_SL g5752 ( 
.A(n_5137),
.B(n_3563),
.Y(n_5752)
);

CKINVDCx5p33_ASAP7_75t_R g5753 ( 
.A(n_4456),
.Y(n_5753)
);

INVx5_ASAP7_75t_L g5754 ( 
.A(n_4568),
.Y(n_5754)
);

NOR2xp33_ASAP7_75t_L g5755 ( 
.A(n_5037),
.B(n_3699),
.Y(n_5755)
);

AOI21xp5_ASAP7_75t_L g5756 ( 
.A1(n_4897),
.A2(n_3553),
.B(n_3573),
.Y(n_5756)
);

NOR2xp33_ASAP7_75t_L g5757 ( 
.A(n_5037),
.B(n_3699),
.Y(n_5757)
);

NOR2xp33_ASAP7_75t_L g5758 ( 
.A(n_4633),
.B(n_3675),
.Y(n_5758)
);

NAND2xp5_ASAP7_75t_SL g5759 ( 
.A(n_4669),
.B(n_3563),
.Y(n_5759)
);

CKINVDCx6p67_ASAP7_75t_R g5760 ( 
.A(n_4723),
.Y(n_5760)
);

AND2x4_ASAP7_75t_L g5761 ( 
.A(n_4500),
.B(n_4250),
.Y(n_5761)
);

NAND2xp5_ASAP7_75t_L g5762 ( 
.A(n_4999),
.B(n_4250),
.Y(n_5762)
);

NAND2xp5_ASAP7_75t_L g5763 ( 
.A(n_5022),
.B(n_4250),
.Y(n_5763)
);

NAND2xp5_ASAP7_75t_L g5764 ( 
.A(n_5022),
.B(n_4250),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_SL g5765 ( 
.A(n_4669),
.B(n_3563),
.Y(n_5765)
);

AO21x2_ASAP7_75t_L g5766 ( 
.A1(n_4939),
.A2(n_3653),
.B(n_3675),
.Y(n_5766)
);

AOI22xp5_ASAP7_75t_L g5767 ( 
.A1(n_4633),
.A2(n_3335),
.B1(n_3753),
.B2(n_3296),
.Y(n_5767)
);

BUFx6f_ASAP7_75t_L g5768 ( 
.A(n_4504),
.Y(n_5768)
);

AOI21xp5_ASAP7_75t_L g5769 ( 
.A1(n_4939),
.A2(n_3553),
.B(n_3510),
.Y(n_5769)
);

INVx3_ASAP7_75t_L g5770 ( 
.A(n_4945),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_4756),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5156),
.B(n_4249),
.Y(n_5772)
);

AOI22xp33_ASAP7_75t_SL g5773 ( 
.A1(n_4505),
.A2(n_3335),
.B1(n_3296),
.B2(n_3753),
.Y(n_5773)
);

NAND2xp5_ASAP7_75t_L g5774 ( 
.A(n_5156),
.B(n_4249),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_4477),
.Y(n_5775)
);

A2O1A1Ixp33_ASAP7_75t_SL g5776 ( 
.A1(n_4806),
.A2(n_3696),
.B(n_3691),
.C(n_3677),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_4779),
.Y(n_5777)
);

OAI22xp5_ASAP7_75t_L g5778 ( 
.A1(n_4454),
.A2(n_3711),
.B1(n_3656),
.B2(n_3717),
.Y(n_5778)
);

BUFx6f_ASAP7_75t_L g5779 ( 
.A(n_4504),
.Y(n_5779)
);

BUFx8_ASAP7_75t_SL g5780 ( 
.A(n_4501),
.Y(n_5780)
);

INVx1_ASAP7_75t_SL g5781 ( 
.A(n_4480),
.Y(n_5781)
);

O2A1O1Ixp5_ASAP7_75t_L g5782 ( 
.A1(n_5088),
.A2(n_3394),
.B(n_3380),
.C(n_3396),
.Y(n_5782)
);

INVx2_ASAP7_75t_SL g5783 ( 
.A(n_4945),
.Y(n_5783)
);

INVx3_ASAP7_75t_L g5784 ( 
.A(n_4945),
.Y(n_5784)
);

OAI22x1_ASAP7_75t_L g5785 ( 
.A1(n_4717),
.A2(n_3683),
.B1(n_3671),
.B2(n_3677),
.Y(n_5785)
);

A2O1A1Ixp33_ASAP7_75t_L g5786 ( 
.A1(n_4915),
.A2(n_3387),
.B(n_3573),
.C(n_3525),
.Y(n_5786)
);

BUFx6f_ASAP7_75t_L g5787 ( 
.A(n_4504),
.Y(n_5787)
);

INVxp67_ASAP7_75t_SL g5788 ( 
.A(n_5098),
.Y(n_5788)
);

CKINVDCx8_ASAP7_75t_R g5789 ( 
.A(n_5467),
.Y(n_5789)
);

BUFx3_ASAP7_75t_L g5790 ( 
.A(n_5367),
.Y(n_5790)
);

OAI22xp5_ASAP7_75t_L g5791 ( 
.A1(n_4781),
.A2(n_3717),
.B1(n_3672),
.B2(n_3670),
.Y(n_5791)
);

OAI22xp5_ASAP7_75t_L g5792 ( 
.A1(n_4781),
.A2(n_3717),
.B1(n_3683),
.B2(n_3671),
.Y(n_5792)
);

INVx3_ASAP7_75t_L g5793 ( 
.A(n_4945),
.Y(n_5793)
);

NAND2xp5_ASAP7_75t_L g5794 ( 
.A(n_5077),
.B(n_3396),
.Y(n_5794)
);

AND2x2_ASAP7_75t_L g5795 ( 
.A(n_4500),
.B(n_4504),
.Y(n_5795)
);

O2A1O1Ixp33_ASAP7_75t_L g5796 ( 
.A1(n_4613),
.A2(n_3664),
.B(n_3661),
.C(n_3651),
.Y(n_5796)
);

OAI22xp5_ASAP7_75t_L g5797 ( 
.A1(n_4824),
.A2(n_3717),
.B1(n_3387),
.B2(n_3664),
.Y(n_5797)
);

BUFx12f_ASAP7_75t_L g5798 ( 
.A(n_5424),
.Y(n_5798)
);

OR2x6_ASAP7_75t_L g5799 ( 
.A(n_4504),
.B(n_3162),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_4779),
.Y(n_5800)
);

AND2x6_ASAP7_75t_L g5801 ( 
.A(n_5206),
.B(n_5229),
.Y(n_5801)
);

AOI21xp5_ASAP7_75t_L g5802 ( 
.A1(n_5002),
.A2(n_5221),
.B(n_5195),
.Y(n_5802)
);

BUFx4f_ASAP7_75t_L g5803 ( 
.A(n_4973),
.Y(n_5803)
);

A2O1A1Ixp33_ASAP7_75t_L g5804 ( 
.A1(n_4915),
.A2(n_3387),
.B(n_3573),
.C(n_3525),
.Y(n_5804)
);

CKINVDCx5p33_ASAP7_75t_R g5805 ( 
.A(n_4477),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_4779),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_4783),
.Y(n_5807)
);

AND2x4_ASAP7_75t_L g5808 ( 
.A(n_4500),
.B(n_3394),
.Y(n_5808)
);

AND2x4_ASAP7_75t_L g5809 ( 
.A(n_4500),
.B(n_3394),
.Y(n_5809)
);

BUFx6f_ASAP7_75t_L g5810 ( 
.A(n_4504),
.Y(n_5810)
);

INVx3_ASAP7_75t_SL g5811 ( 
.A(n_5217),
.Y(n_5811)
);

BUFx6f_ASAP7_75t_L g5812 ( 
.A(n_4504),
.Y(n_5812)
);

NAND2xp5_ASAP7_75t_L g5813 ( 
.A(n_5077),
.B(n_3396),
.Y(n_5813)
);

AOI22xp5_ASAP7_75t_L g5814 ( 
.A1(n_4787),
.A2(n_3661),
.B1(n_3175),
.B2(n_3269),
.Y(n_5814)
);

CKINVDCx20_ASAP7_75t_R g5815 ( 
.A(n_4636),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_4783),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_4783),
.Y(n_5817)
);

OAI221xp5_ASAP7_75t_L g5818 ( 
.A1(n_4659),
.A2(n_3650),
.B1(n_3660),
.B2(n_3651),
.C(n_3716),
.Y(n_5818)
);

NOR3xp33_ASAP7_75t_L g5819 ( 
.A(n_4720),
.B(n_3689),
.C(n_3688),
.Y(n_5819)
);

BUFx3_ASAP7_75t_L g5820 ( 
.A(n_5367),
.Y(n_5820)
);

NOR2xp33_ASAP7_75t_L g5821 ( 
.A(n_4643),
.B(n_3394),
.Y(n_5821)
);

INVx3_ASAP7_75t_L g5822 ( 
.A(n_4945),
.Y(n_5822)
);

BUFx3_ASAP7_75t_L g5823 ( 
.A(n_5367),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_4793),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_4793),
.Y(n_5825)
);

NAND2xp5_ASAP7_75t_SL g5826 ( 
.A(n_4717),
.B(n_3511),
.Y(n_5826)
);

INVx4_ASAP7_75t_L g5827 ( 
.A(n_5393),
.Y(n_5827)
);

AOI22xp33_ASAP7_75t_L g5828 ( 
.A1(n_4701),
.A2(n_3660),
.B1(n_3650),
.B2(n_3269),
.Y(n_5828)
);

INVx5_ASAP7_75t_L g5829 ( 
.A(n_4568),
.Y(n_5829)
);

INVx4_ASAP7_75t_L g5830 ( 
.A(n_5393),
.Y(n_5830)
);

INVx5_ASAP7_75t_L g5831 ( 
.A(n_4568),
.Y(n_5831)
);

AO21x1_ASAP7_75t_L g5832 ( 
.A1(n_4740),
.A2(n_3380),
.B(n_3573),
.Y(n_5832)
);

INVx3_ASAP7_75t_L g5833 ( 
.A(n_4945),
.Y(n_5833)
);

BUFx8_ASAP7_75t_L g5834 ( 
.A(n_4775),
.Y(n_5834)
);

AOI22xp33_ASAP7_75t_L g5835 ( 
.A1(n_4701),
.A2(n_3162),
.B1(n_3175),
.B2(n_4209),
.Y(n_5835)
);

NAND2xp5_ASAP7_75t_L g5836 ( 
.A(n_5140),
.B(n_3380),
.Y(n_5836)
);

AOI21xp5_ASAP7_75t_L g5837 ( 
.A1(n_5002),
.A2(n_3510),
.B(n_3525),
.Y(n_5837)
);

INVx1_ASAP7_75t_SL g5838 ( 
.A(n_4496),
.Y(n_5838)
);

OAI21xp33_ASAP7_75t_L g5839 ( 
.A1(n_4455),
.A2(n_3687),
.B(n_3716),
.Y(n_5839)
);

AOI21xp5_ASAP7_75t_L g5840 ( 
.A1(n_5195),
.A2(n_3510),
.B(n_3525),
.Y(n_5840)
);

AOI22xp5_ASAP7_75t_L g5841 ( 
.A1(n_4787),
.A2(n_4836),
.B1(n_4837),
.B2(n_4833),
.Y(n_5841)
);

AND2x6_ASAP7_75t_L g5842 ( 
.A(n_5206),
.B(n_3571),
.Y(n_5842)
);

INVxp67_ASAP7_75t_SL g5843 ( 
.A(n_5108),
.Y(n_5843)
);

NAND2x1_ASAP7_75t_L g5844 ( 
.A(n_4680),
.B(n_4448),
.Y(n_5844)
);

AO21x2_ASAP7_75t_L g5845 ( 
.A1(n_5221),
.A2(n_3380),
.B(n_3510),
.Y(n_5845)
);

A2O1A1Ixp33_ASAP7_75t_L g5846 ( 
.A1(n_4419),
.A2(n_3412),
.B(n_4209),
.C(n_3979),
.Y(n_5846)
);

O2A1O1Ixp33_ASAP7_75t_SL g5847 ( 
.A1(n_4419),
.A2(n_3412),
.B(n_3979),
.C(n_3900),
.Y(n_5847)
);

AOI21xp33_ASAP7_75t_L g5848 ( 
.A1(n_4511),
.A2(n_3432),
.B(n_3479),
.Y(n_5848)
);

OAI22xp5_ASAP7_75t_L g5849 ( 
.A1(n_4824),
.A2(n_3432),
.B1(n_3479),
.B2(n_3511),
.Y(n_5849)
);

BUFx6f_ASAP7_75t_L g5850 ( 
.A(n_4504),
.Y(n_5850)
);

AOI22xp5_ASAP7_75t_L g5851 ( 
.A1(n_4833),
.A2(n_4837),
.B1(n_4853),
.B2(n_4836),
.Y(n_5851)
);

NAND2xp5_ASAP7_75t_L g5852 ( 
.A(n_5140),
.B(n_3691),
.Y(n_5852)
);

AND2x2_ASAP7_75t_L g5853 ( 
.A(n_4509),
.B(n_3691),
.Y(n_5853)
);

A2O1A1Ixp33_ASAP7_75t_L g5854 ( 
.A1(n_4616),
.A2(n_4248),
.B(n_3900),
.C(n_3799),
.Y(n_5854)
);

AOI22xp33_ASAP7_75t_L g5855 ( 
.A1(n_4735),
.A2(n_4248),
.B1(n_3799),
.B2(n_3790),
.Y(n_5855)
);

INVxp67_ASAP7_75t_L g5856 ( 
.A(n_5167),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_4981),
.B(n_3691),
.Y(n_5857)
);

BUFx3_ASAP7_75t_L g5858 ( 
.A(n_5367),
.Y(n_5858)
);

BUFx6f_ASAP7_75t_L g5859 ( 
.A(n_4509),
.Y(n_5859)
);

NAND2x1p5_ASAP7_75t_L g5860 ( 
.A(n_5393),
.B(n_3432),
.Y(n_5860)
);

INVx4_ASAP7_75t_L g5861 ( 
.A(n_5393),
.Y(n_5861)
);

INVx4_ASAP7_75t_L g5862 ( 
.A(n_5393),
.Y(n_5862)
);

AOI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_4853),
.A2(n_3790),
.B1(n_3556),
.B2(n_3687),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_4509),
.B(n_3677),
.Y(n_5864)
);

NAND2xp5_ASAP7_75t_L g5865 ( 
.A(n_4981),
.B(n_3432),
.Y(n_5865)
);

AND2x2_ASAP7_75t_L g5866 ( 
.A(n_4509),
.B(n_3479),
.Y(n_5866)
);

OR2x2_ASAP7_75t_L g5867 ( 
.A(n_5309),
.B(n_3479),
.Y(n_5867)
);

AOI22xp33_ASAP7_75t_L g5868 ( 
.A1(n_4735),
.A2(n_3556),
.B1(n_3687),
.B2(n_3479),
.Y(n_5868)
);

BUFx6f_ASAP7_75t_L g5869 ( 
.A(n_4509),
.Y(n_5869)
);

INVxp67_ASAP7_75t_SL g5870 ( 
.A(n_5108),
.Y(n_5870)
);

INVx3_ASAP7_75t_SL g5871 ( 
.A(n_4680),
.Y(n_5871)
);

OAI22xp5_ASAP7_75t_L g5872 ( 
.A1(n_4910),
.A2(n_3479),
.B1(n_3511),
.B2(n_3563),
.Y(n_5872)
);

AND2x2_ASAP7_75t_L g5873 ( 
.A(n_4509),
.B(n_3511),
.Y(n_5873)
);

O2A1O1Ixp33_ASAP7_75t_L g5874 ( 
.A1(n_4661),
.A2(n_3690),
.B(n_3563),
.C(n_3571),
.Y(n_5874)
);

AOI21xp5_ASAP7_75t_L g5875 ( 
.A1(n_5273),
.A2(n_5131),
.B(n_5130),
.Y(n_5875)
);

BUFx3_ASAP7_75t_L g5876 ( 
.A(n_5198),
.Y(n_5876)
);

AOI22xp33_ASAP7_75t_L g5877 ( 
.A1(n_4505),
.A2(n_3511),
.B1(n_3563),
.B2(n_3571),
.Y(n_5877)
);

AOI22xp5_ASAP7_75t_L g5878 ( 
.A1(n_4627),
.A2(n_3690),
.B1(n_3511),
.B2(n_3571),
.Y(n_5878)
);

NOR2xp33_ASAP7_75t_L g5879 ( 
.A(n_5100),
.B(n_3571),
.Y(n_5879)
);

BUFx6f_ASAP7_75t_L g5880 ( 
.A(n_4509),
.Y(n_5880)
);

BUFx3_ASAP7_75t_L g5881 ( 
.A(n_5198),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_SL g5882 ( 
.A(n_4757),
.B(n_3571),
.Y(n_5882)
);

AOI21xp5_ASAP7_75t_L g5883 ( 
.A1(n_5273),
.A2(n_5131),
.B(n_5130),
.Y(n_5883)
);

OAI22xp5_ASAP7_75t_L g5884 ( 
.A1(n_4910),
.A2(n_5009),
.B1(n_4455),
.B2(n_4758),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_4509),
.B(n_4510),
.Y(n_5885)
);

INVx4_ASAP7_75t_L g5886 ( 
.A(n_5393),
.Y(n_5886)
);

NAND2x1_ASAP7_75t_L g5887 ( 
.A(n_4680),
.B(n_4448),
.Y(n_5887)
);

NAND2xp5_ASAP7_75t_L g5888 ( 
.A(n_4981),
.B(n_5158),
.Y(n_5888)
);

A2O1A1Ixp33_ASAP7_75t_L g5889 ( 
.A1(n_4661),
.A2(n_4630),
.B(n_4758),
.C(n_4757),
.Y(n_5889)
);

BUFx3_ASAP7_75t_L g5890 ( 
.A(n_5198),
.Y(n_5890)
);

BUFx6f_ASAP7_75t_SL g5891 ( 
.A(n_4523),
.Y(n_5891)
);

AND3x1_ASAP7_75t_SL g5892 ( 
.A(n_4449),
.B(n_4642),
.C(n_4904),
.Y(n_5892)
);

BUFx6f_ASAP7_75t_L g5893 ( 
.A(n_4509),
.Y(n_5893)
);

O2A1O1Ixp33_ASAP7_75t_SL g5894 ( 
.A1(n_5003),
.A2(n_5030),
.B(n_4992),
.C(n_4440),
.Y(n_5894)
);

BUFx2_ASAP7_75t_R g5895 ( 
.A(n_4624),
.Y(n_5895)
);

OR2x6_ASAP7_75t_L g5896 ( 
.A(n_4510),
.B(n_4517),
.Y(n_5896)
);

O2A1O1Ixp33_ASAP7_75t_L g5897 ( 
.A1(n_4720),
.A2(n_4772),
.B(n_4627),
.C(n_4767),
.Y(n_5897)
);

BUFx2_ASAP7_75t_SL g5898 ( 
.A(n_5372),
.Y(n_5898)
);

BUFx3_ASAP7_75t_L g5899 ( 
.A(n_5198),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_4444),
.Y(n_5900)
);

NAND2xp5_ASAP7_75t_L g5901 ( 
.A(n_5161),
.B(n_5138),
.Y(n_5901)
);

AOI22xp33_ASAP7_75t_L g5902 ( 
.A1(n_4440),
.A2(n_4772),
.B1(n_4653),
.B2(n_4630),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_4535),
.Y(n_5903)
);

OAI22xp5_ASAP7_75t_L g5904 ( 
.A1(n_5009),
.A2(n_4465),
.B1(n_4894),
.B2(n_4626),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_SL g5905 ( 
.A(n_4465),
.B(n_5165),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_L g5906 ( 
.A(n_5100),
.B(n_5214),
.Y(n_5906)
);

NAND2xp5_ASAP7_75t_L g5907 ( 
.A(n_5138),
.B(n_5162),
.Y(n_5907)
);

BUFx3_ASAP7_75t_L g5908 ( 
.A(n_5264),
.Y(n_5908)
);

INVx2_ASAP7_75t_SL g5909 ( 
.A(n_4949),
.Y(n_5909)
);

AOI22xp33_ASAP7_75t_L g5910 ( 
.A1(n_4653),
.A2(n_4628),
.B1(n_4445),
.B2(n_4457),
.Y(n_5910)
);

INVx3_ASAP7_75t_L g5911 ( 
.A(n_4949),
.Y(n_5911)
);

BUFx12f_ASAP7_75t_L g5912 ( 
.A(n_4501),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_L g5913 ( 
.A(n_5162),
.B(n_5169),
.Y(n_5913)
);

INVx4_ASAP7_75t_L g5914 ( 
.A(n_5393),
.Y(n_5914)
);

AOI22xp33_ASAP7_75t_L g5915 ( 
.A1(n_4628),
.A2(n_4445),
.B1(n_4457),
.B2(n_4766),
.Y(n_5915)
);

INVx3_ASAP7_75t_L g5916 ( 
.A(n_4949),
.Y(n_5916)
);

INVx3_ASAP7_75t_SL g5917 ( 
.A(n_4680),
.Y(n_5917)
);

O2A1O1Ixp33_ASAP7_75t_L g5918 ( 
.A1(n_4767),
.A2(n_4848),
.B(n_4992),
.C(n_5086),
.Y(n_5918)
);

OAI21x1_ASAP7_75t_SL g5919 ( 
.A1(n_5331),
.A2(n_5351),
.B(n_5345),
.Y(n_5919)
);

OR2x2_ASAP7_75t_L g5920 ( 
.A(n_5464),
.B(n_5471),
.Y(n_5920)
);

INVx2_ASAP7_75t_SL g5921 ( 
.A(n_4949),
.Y(n_5921)
);

BUFx6f_ASAP7_75t_L g5922 ( 
.A(n_4510),
.Y(n_5922)
);

INVxp67_ASAP7_75t_L g5923 ( 
.A(n_4964),
.Y(n_5923)
);

INVx3_ASAP7_75t_L g5924 ( 
.A(n_4949),
.Y(n_5924)
);

A2O1A1Ixp33_ASAP7_75t_L g5925 ( 
.A1(n_5111),
.A2(n_5003),
.B(n_5030),
.C(n_4955),
.Y(n_5925)
);

NAND2xp5_ASAP7_75t_SL g5926 ( 
.A(n_4446),
.B(n_4955),
.Y(n_5926)
);

OAI22xp33_ASAP7_75t_L g5927 ( 
.A1(n_5111),
.A2(n_4975),
.B1(n_4884),
.B2(n_4869),
.Y(n_5927)
);

INVx3_ASAP7_75t_L g5928 ( 
.A(n_4949),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_5175),
.B(n_5322),
.Y(n_5929)
);

BUFx6f_ASAP7_75t_L g5930 ( 
.A(n_4510),
.Y(n_5930)
);

OAI22xp5_ASAP7_75t_L g5931 ( 
.A1(n_4894),
.A2(n_4626),
.B1(n_4621),
.B2(n_4924),
.Y(n_5931)
);

BUFx2_ASAP7_75t_L g5932 ( 
.A(n_5421),
.Y(n_5932)
);

BUFx12f_ASAP7_75t_L g5933 ( 
.A(n_4508),
.Y(n_5933)
);

BUFx3_ASAP7_75t_L g5934 ( 
.A(n_5264),
.Y(n_5934)
);

INVx1_ASAP7_75t_SL g5935 ( 
.A(n_4496),
.Y(n_5935)
);

INVx3_ASAP7_75t_L g5936 ( 
.A(n_4949),
.Y(n_5936)
);

AND2x2_ASAP7_75t_L g5937 ( 
.A(n_4510),
.B(n_4517),
.Y(n_5937)
);

OAI21xp33_ASAP7_75t_L g5938 ( 
.A1(n_4975),
.A2(n_4621),
.B(n_4473),
.Y(n_5938)
);

O2A1O1Ixp5_ASAP7_75t_SL g5939 ( 
.A1(n_4740),
.A2(n_4751),
.B(n_4759),
.C(n_5032),
.Y(n_5939)
);

AOI21x1_ASAP7_75t_L g5940 ( 
.A1(n_4760),
.A2(n_4635),
.B(n_4645),
.Y(n_5940)
);

AOI22xp5_ASAP7_75t_L g5941 ( 
.A1(n_4514),
.A2(n_4766),
.B1(n_5101),
.B2(n_5210),
.Y(n_5941)
);

NAND2xp5_ASAP7_75t_SL g5942 ( 
.A(n_4446),
.B(n_4904),
.Y(n_5942)
);

AOI21xp5_ASAP7_75t_L g5943 ( 
.A1(n_5455),
.A2(n_4760),
.B(n_5342),
.Y(n_5943)
);

AOI21xp5_ASAP7_75t_SL g5944 ( 
.A1(n_4848),
.A2(n_5380),
.B(n_4759),
.Y(n_5944)
);

OR2x2_ASAP7_75t_L g5945 ( 
.A(n_5464),
.B(n_5471),
.Y(n_5945)
);

BUFx12f_ASAP7_75t_L g5946 ( 
.A(n_4508),
.Y(n_5946)
);

A2O1A1Ixp33_ASAP7_75t_L g5947 ( 
.A1(n_5122),
.A2(n_5210),
.B(n_4718),
.C(n_4483),
.Y(n_5947)
);

A2O1A1Ixp33_ASAP7_75t_L g5948 ( 
.A1(n_5122),
.A2(n_4718),
.B(n_4483),
.C(n_4751),
.Y(n_5948)
);

BUFx6f_ASAP7_75t_L g5949 ( 
.A(n_4510),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_4535),
.Y(n_5950)
);

NAND2xp5_ASAP7_75t_SL g5951 ( 
.A(n_4446),
.B(n_4584),
.Y(n_5951)
);

BUFx2_ASAP7_75t_L g5952 ( 
.A(n_5421),
.Y(n_5952)
);

AOI22xp5_ASAP7_75t_L g5953 ( 
.A1(n_4514),
.A2(n_4766),
.B1(n_5101),
.B2(n_5258),
.Y(n_5953)
);

INVx1_ASAP7_75t_SL g5954 ( 
.A(n_4673),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_4554),
.Y(n_5955)
);

NAND2xp5_ASAP7_75t_L g5956 ( 
.A(n_5322),
.B(n_5062),
.Y(n_5956)
);

NAND2xp5_ASAP7_75t_L g5957 ( 
.A(n_5062),
.B(n_5024),
.Y(n_5957)
);

AOI21xp5_ASAP7_75t_L g5958 ( 
.A1(n_5455),
.A2(n_5342),
.B(n_4563),
.Y(n_5958)
);

INVx4_ASAP7_75t_L g5959 ( 
.A(n_5393),
.Y(n_5959)
);

BUFx6f_ASAP7_75t_SL g5960 ( 
.A(n_4523),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_L g5961 ( 
.A(n_5062),
.B(n_5024),
.Y(n_5961)
);

BUFx2_ASAP7_75t_L g5962 ( 
.A(n_5421),
.Y(n_5962)
);

BUFx6f_ASAP7_75t_L g5963 ( 
.A(n_4510),
.Y(n_5963)
);

A2O1A1Ixp33_ASAP7_75t_L g5964 ( 
.A1(n_5038),
.A2(n_5157),
.B(n_5086),
.C(n_4473),
.Y(n_5964)
);

CKINVDCx5p33_ASAP7_75t_R g5965 ( 
.A(n_4554),
.Y(n_5965)
);

A2O1A1Ixp33_ASAP7_75t_L g5966 ( 
.A1(n_5038),
.A2(n_5157),
.B(n_4642),
.C(n_5079),
.Y(n_5966)
);

INVx1_ASAP7_75t_SL g5967 ( 
.A(n_4673),
.Y(n_5967)
);

OR2x2_ASAP7_75t_L g5968 ( 
.A(n_5464),
.B(n_5471),
.Y(n_5968)
);

NAND2x1_ASAP7_75t_SL g5969 ( 
.A(n_5048),
.B(n_5085),
.Y(n_5969)
);

AOI21xp5_ASAP7_75t_L g5970 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_5970)
);

NOR2xp33_ASAP7_75t_R g5971 ( 
.A(n_4724),
.B(n_4529),
.Y(n_5971)
);

BUFx2_ASAP7_75t_L g5972 ( 
.A(n_5421),
.Y(n_5972)
);

BUFx12f_ASAP7_75t_L g5973 ( 
.A(n_4529),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_SL g5974 ( 
.A(n_4584),
.B(n_5280),
.Y(n_5974)
);

OR2x4_ASAP7_75t_L g5975 ( 
.A(n_4849),
.B(n_5001),
.Y(n_5975)
);

AOI22xp5_ASAP7_75t_L g5976 ( 
.A1(n_4766),
.A2(n_5258),
.B1(n_4993),
.B2(n_5019),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_SL g5977 ( 
.A(n_4584),
.B(n_5280),
.Y(n_5977)
);

BUFx12f_ASAP7_75t_L g5978 ( 
.A(n_4532),
.Y(n_5978)
);

NOR2xp33_ASAP7_75t_L g5979 ( 
.A(n_5214),
.B(n_5082),
.Y(n_5979)
);

AOI21xp5_ASAP7_75t_L g5980 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_5980)
);

AOI22xp5_ASAP7_75t_L g5981 ( 
.A1(n_4766),
.A2(n_4993),
.B1(n_5019),
.B2(n_4947),
.Y(n_5981)
);

AOI22xp5_ASAP7_75t_L g5982 ( 
.A1(n_4766),
.A2(n_4996),
.B1(n_4947),
.B2(n_5102),
.Y(n_5982)
);

NOR2xp33_ASAP7_75t_L g5983 ( 
.A(n_5082),
.B(n_5091),
.Y(n_5983)
);

INVx4_ASAP7_75t_L g5984 ( 
.A(n_4885),
.Y(n_5984)
);

INVxp67_ASAP7_75t_SL g5985 ( 
.A(n_5035),
.Y(n_5985)
);

OR2x2_ASAP7_75t_SL g5986 ( 
.A(n_5277),
.B(n_5024),
.Y(n_5986)
);

CKINVDCx11_ASAP7_75t_R g5987 ( 
.A(n_5306),
.Y(n_5987)
);

A2O1A1Ixp33_ASAP7_75t_L g5988 ( 
.A1(n_5079),
.A2(n_4635),
.B(n_5313),
.C(n_4755),
.Y(n_5988)
);

A2O1A1Ixp33_ASAP7_75t_L g5989 ( 
.A1(n_5313),
.A2(n_4755),
.B(n_4584),
.C(n_5351),
.Y(n_5989)
);

CKINVDCx5p33_ASAP7_75t_R g5990 ( 
.A(n_5425),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_5425),
.Y(n_5991)
);

INVx3_ASAP7_75t_L g5992 ( 
.A(n_4959),
.Y(n_5992)
);

NAND2xp5_ASAP7_75t_SL g5993 ( 
.A(n_4869),
.B(n_4884),
.Y(n_5993)
);

NAND2xp5_ASAP7_75t_L g5994 ( 
.A(n_5053),
.B(n_4807),
.Y(n_5994)
);

INVx3_ASAP7_75t_SL g5995 ( 
.A(n_4680),
.Y(n_5995)
);

BUFx2_ASAP7_75t_L g5996 ( 
.A(n_5456),
.Y(n_5996)
);

INVx8_ASAP7_75t_L g5997 ( 
.A(n_4865),
.Y(n_5997)
);

BUFx2_ASAP7_75t_L g5998 ( 
.A(n_5456),
.Y(n_5998)
);

INVx3_ASAP7_75t_L g5999 ( 
.A(n_4959),
.Y(n_5999)
);

AND2x2_ASAP7_75t_SL g6000 ( 
.A(n_5154),
.B(n_5155),
.Y(n_6000)
);

AOI21xp5_ASAP7_75t_L g6001 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5053),
.B(n_4807),
.Y(n_6002)
);

NAND2xp5_ASAP7_75t_SL g6003 ( 
.A(n_5094),
.B(n_5048),
.Y(n_6003)
);

AOI21x1_ASAP7_75t_L g6004 ( 
.A1(n_4645),
.A2(n_5422),
.B(n_4481),
.Y(n_6004)
);

AOI21xp5_ASAP7_75t_L g6005 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_6005)
);

O2A1O1Ixp33_ASAP7_75t_L g6006 ( 
.A1(n_4996),
.A2(n_4840),
.B(n_4892),
.C(n_4784),
.Y(n_6006)
);

NOR2xp33_ASAP7_75t_L g6007 ( 
.A(n_5091),
.B(n_5102),
.Y(n_6007)
);

BUFx12f_ASAP7_75t_L g6008 ( 
.A(n_4532),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_4810),
.B(n_4849),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_4835),
.Y(n_6010)
);

NAND2xp5_ASAP7_75t_L g6011 ( 
.A(n_4810),
.B(n_4490),
.Y(n_6011)
);

NAND3xp33_ASAP7_75t_L g6012 ( 
.A(n_5094),
.B(n_4615),
.C(n_5120),
.Y(n_6012)
);

INVx1_ASAP7_75t_SL g6013 ( 
.A(n_4727),
.Y(n_6013)
);

BUFx6f_ASAP7_75t_L g6014 ( 
.A(n_4510),
.Y(n_6014)
);

AOI21xp5_ASAP7_75t_L g6015 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_6015)
);

BUFx2_ASAP7_75t_L g6016 ( 
.A(n_5456),
.Y(n_6016)
);

BUFx3_ASAP7_75t_L g6017 ( 
.A(n_5264),
.Y(n_6017)
);

OAI22xp5_ASAP7_75t_L g6018 ( 
.A1(n_4894),
.A2(n_4924),
.B1(n_4991),
.B2(n_5134),
.Y(n_6018)
);

NOR2xp33_ASAP7_75t_L g6019 ( 
.A(n_5252),
.B(n_4797),
.Y(n_6019)
);

AOI22xp33_ASAP7_75t_L g6020 ( 
.A1(n_4937),
.A2(n_4954),
.B1(n_4521),
.B2(n_5168),
.Y(n_6020)
);

BUFx6f_ASAP7_75t_L g6021 ( 
.A(n_4510),
.Y(n_6021)
);

INVx1_ASAP7_75t_SL g6022 ( 
.A(n_4727),
.Y(n_6022)
);

INVx3_ASAP7_75t_L g6023 ( 
.A(n_4959),
.Y(n_6023)
);

BUFx8_ASAP7_75t_L g6024 ( 
.A(n_4775),
.Y(n_6024)
);

BUFx6f_ASAP7_75t_L g6025 ( 
.A(n_4517),
.Y(n_6025)
);

INVx3_ASAP7_75t_L g6026 ( 
.A(n_4959),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_4517),
.B(n_5458),
.Y(n_6027)
);

OAI22xp5_ASAP7_75t_L g6028 ( 
.A1(n_4991),
.A2(n_5134),
.B1(n_4574),
.B2(n_5120),
.Y(n_6028)
);

OAI22xp5_ASAP7_75t_L g6029 ( 
.A1(n_4574),
.A2(n_5105),
.B1(n_4488),
.B2(n_4489),
.Y(n_6029)
);

O2A1O1Ixp33_ASAP7_75t_L g6030 ( 
.A1(n_4784),
.A2(n_4892),
.B(n_4893),
.C(n_4840),
.Y(n_6030)
);

BUFx2_ASAP7_75t_L g6031 ( 
.A(n_5456),
.Y(n_6031)
);

OAI22xp5_ASAP7_75t_L g6032 ( 
.A1(n_4574),
.A2(n_5105),
.B1(n_4488),
.B2(n_4489),
.Y(n_6032)
);

AOI22xp33_ASAP7_75t_L g6033 ( 
.A1(n_4937),
.A2(n_4954),
.B1(n_4521),
.B2(n_5168),
.Y(n_6033)
);

AOI21xp5_ASAP7_75t_L g6034 ( 
.A1(n_4479),
.A2(n_4712),
.B(n_4563),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_4490),
.B(n_4491),
.Y(n_6035)
);

OAI21xp33_ASAP7_75t_L g6036 ( 
.A1(n_5335),
.A2(n_5247),
.B(n_5106),
.Y(n_6036)
);

AOI22xp5_ASAP7_75t_L g6037 ( 
.A1(n_5247),
.A2(n_4881),
.B1(n_5123),
.B2(n_4499),
.Y(n_6037)
);

BUFx12f_ASAP7_75t_L g6038 ( 
.A(n_4594),
.Y(n_6038)
);

CKINVDCx5p33_ASAP7_75t_R g6039 ( 
.A(n_4835),
.Y(n_6039)
);

NAND2xp5_ASAP7_75t_SL g6040 ( 
.A(n_4615),
.B(n_5335),
.Y(n_6040)
);

CKINVDCx20_ASAP7_75t_R g6041 ( 
.A(n_4990),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_4470),
.Y(n_6042)
);

NOR2xp33_ASAP7_75t_L g6043 ( 
.A(n_5252),
.B(n_4797),
.Y(n_6043)
);

BUFx2_ASAP7_75t_L g6044 ( 
.A(n_5527),
.Y(n_6044)
);

OAI21xp5_ASAP7_75t_L g6045 ( 
.A1(n_4481),
.A2(n_4615),
.B(n_4763),
.Y(n_6045)
);

NOR2xp33_ASAP7_75t_L g6046 ( 
.A(n_4797),
.B(n_4817),
.Y(n_6046)
);

O2A1O1Ixp33_ASAP7_75t_L g6047 ( 
.A1(n_4893),
.A2(n_4956),
.B(n_5008),
.C(n_4952),
.Y(n_6047)
);

AOI22xp33_ASAP7_75t_L g6048 ( 
.A1(n_4937),
.A2(n_4954),
.B1(n_5106),
.B2(n_4667),
.Y(n_6048)
);

AOI21xp5_ASAP7_75t_L g6049 ( 
.A1(n_4479),
.A2(n_4715),
.B(n_4712),
.Y(n_6049)
);

INVx1_ASAP7_75t_SL g6050 ( 
.A(n_4764),
.Y(n_6050)
);

BUFx6f_ASAP7_75t_L g6051 ( 
.A(n_4517),
.Y(n_6051)
);

O2A1O1Ixp33_ASAP7_75t_L g6052 ( 
.A1(n_4952),
.A2(n_5008),
.B(n_5041),
.C(n_4956),
.Y(n_6052)
);

AOI21xp5_ASAP7_75t_L g6053 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6053)
);

AOI21xp5_ASAP7_75t_L g6054 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6054)
);

INVx3_ASAP7_75t_L g6055 ( 
.A(n_4959),
.Y(n_6055)
);

AOI22xp5_ASAP7_75t_L g6056 ( 
.A1(n_4881),
.A2(n_5123),
.B1(n_4499),
.B2(n_4528),
.Y(n_6056)
);

NAND2x2_ASAP7_75t_L g6057 ( 
.A(n_5372),
.B(n_5410),
.Y(n_6057)
);

INVx1_ASAP7_75t_SL g6058 ( 
.A(n_4764),
.Y(n_6058)
);

A2O1A1Ixp33_ASAP7_75t_L g6059 ( 
.A1(n_5154),
.A2(n_5155),
.B(n_4763),
.C(n_5061),
.Y(n_6059)
);

AOI21xp5_ASAP7_75t_L g6060 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_4470),
.Y(n_6061)
);

INVx2_ASAP7_75t_L g6062 ( 
.A(n_4470),
.Y(n_6062)
);

AOI22xp5_ASAP7_75t_L g6063 ( 
.A1(n_4485),
.A2(n_4528),
.B1(n_4564),
.B2(n_4546),
.Y(n_6063)
);

NAND3xp33_ASAP7_75t_L g6064 ( 
.A(n_5181),
.B(n_4493),
.C(n_5041),
.Y(n_6064)
);

BUFx6f_ASAP7_75t_L g6065 ( 
.A(n_4517),
.Y(n_6065)
);

NAND2xp5_ASAP7_75t_L g6066 ( 
.A(n_4491),
.B(n_4498),
.Y(n_6066)
);

OAI22xp5_ASAP7_75t_L g6067 ( 
.A1(n_5292),
.A2(n_4546),
.B1(n_4564),
.B2(n_4485),
.Y(n_6067)
);

INVx3_ASAP7_75t_L g6068 ( 
.A(n_4959),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_4517),
.B(n_5458),
.Y(n_6069)
);

NAND2x1p5_ASAP7_75t_L g6070 ( 
.A(n_4523),
.B(n_4709),
.Y(n_6070)
);

BUFx6f_ASAP7_75t_L g6071 ( 
.A(n_4517),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_4498),
.B(n_4506),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_4476),
.Y(n_6073)
);

NAND2xp33_ASAP7_75t_L g6074 ( 
.A(n_4667),
.B(n_5107),
.Y(n_6074)
);

INVx2_ASAP7_75t_L g6075 ( 
.A(n_4476),
.Y(n_6075)
);

O2A1O1Ixp5_ASAP7_75t_L g6076 ( 
.A1(n_4493),
.A2(n_4526),
.B(n_5016),
.C(n_4846),
.Y(n_6076)
);

NAND2xp5_ASAP7_75t_SL g6077 ( 
.A(n_5423),
.B(n_4973),
.Y(n_6077)
);

AOI21xp5_ASAP7_75t_L g6078 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6078)
);

AOI21x1_ASAP7_75t_L g6079 ( 
.A1(n_5422),
.A2(n_5039),
.B(n_5032),
.Y(n_6079)
);

INVx3_ASAP7_75t_L g6080 ( 
.A(n_4965),
.Y(n_6080)
);

NAND2xp5_ASAP7_75t_L g6081 ( 
.A(n_4506),
.B(n_4512),
.Y(n_6081)
);

BUFx4f_ASAP7_75t_L g6082 ( 
.A(n_4973),
.Y(n_6082)
);

AND2x6_ASAP7_75t_L g6083 ( 
.A(n_5206),
.B(n_5229),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_SL g6084 ( 
.A(n_5423),
.B(n_5149),
.Y(n_6084)
);

A2O1A1Ixp33_ASAP7_75t_L g6085 ( 
.A1(n_5154),
.A2(n_5155),
.B(n_5064),
.C(n_5065),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_4512),
.B(n_4513),
.Y(n_6086)
);

BUFx3_ASAP7_75t_L g6087 ( 
.A(n_5264),
.Y(n_6087)
);

INVx3_ASAP7_75t_L g6088 ( 
.A(n_4965),
.Y(n_6088)
);

INVx3_ASAP7_75t_L g6089 ( 
.A(n_4965),
.Y(n_6089)
);

OAI21xp5_ASAP7_75t_L g6090 ( 
.A1(n_5164),
.A2(n_5194),
.B(n_5174),
.Y(n_6090)
);

AOI21xp5_ASAP7_75t_L g6091 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6091)
);

INVx3_ASAP7_75t_L g6092 ( 
.A(n_4965),
.Y(n_6092)
);

INVx3_ASAP7_75t_L g6093 ( 
.A(n_4965),
.Y(n_6093)
);

AOI22xp5_ASAP7_75t_L g6094 ( 
.A1(n_4586),
.A2(n_4600),
.B1(n_4749),
.B2(n_4736),
.Y(n_6094)
);

OR2x6_ASAP7_75t_L g6095 ( 
.A(n_4517),
.B(n_5503),
.Y(n_6095)
);

CKINVDCx8_ASAP7_75t_R g6096 ( 
.A(n_5467),
.Y(n_6096)
);

BUFx6f_ASAP7_75t_L g6097 ( 
.A(n_4547),
.Y(n_6097)
);

NAND2xp5_ASAP7_75t_L g6098 ( 
.A(n_4513),
.B(n_4515),
.Y(n_6098)
);

AOI22xp33_ASAP7_75t_L g6099 ( 
.A1(n_5107),
.A2(n_5177),
.B1(n_4586),
.B2(n_4600),
.Y(n_6099)
);

O2A1O1Ixp33_ASAP7_75t_L g6100 ( 
.A1(n_5061),
.A2(n_5065),
.B(n_5073),
.C(n_5064),
.Y(n_6100)
);

BUFx6f_ASAP7_75t_L g6101 ( 
.A(n_4547),
.Y(n_6101)
);

CKINVDCx8_ASAP7_75t_R g6102 ( 
.A(n_4486),
.Y(n_6102)
);

BUFx2_ASAP7_75t_L g6103 ( 
.A(n_5527),
.Y(n_6103)
);

AOI21xp5_ASAP7_75t_L g6104 ( 
.A1(n_4715),
.A2(n_4883),
.B(n_4857),
.Y(n_6104)
);

NAND2xp5_ASAP7_75t_L g6105 ( 
.A(n_4515),
.B(n_4516),
.Y(n_6105)
);

AOI21xp5_ASAP7_75t_L g6106 ( 
.A1(n_4857),
.A2(n_4890),
.B(n_4883),
.Y(n_6106)
);

OAI21xp33_ASAP7_75t_L g6107 ( 
.A1(n_5177),
.A2(n_5073),
.B(n_4421),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_SL g6108 ( 
.A(n_5149),
.B(n_5352),
.Y(n_6108)
);

BUFx12f_ASAP7_75t_L g6109 ( 
.A(n_4594),
.Y(n_6109)
);

AOI21x1_ASAP7_75t_L g6110 ( 
.A1(n_5422),
.A2(n_5039),
.B(n_5032),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_4516),
.B(n_4522),
.Y(n_6111)
);

INVx3_ASAP7_75t_L g6112 ( 
.A(n_4965),
.Y(n_6112)
);

O2A1O1Ixp33_ASAP7_75t_L g6113 ( 
.A1(n_5243),
.A2(n_5174),
.B(n_5194),
.C(n_5164),
.Y(n_6113)
);

BUFx3_ASAP7_75t_L g6114 ( 
.A(n_5267),
.Y(n_6114)
);

A2O1A1Ixp33_ASAP7_75t_L g6115 ( 
.A1(n_4699),
.A2(n_4421),
.B(n_4482),
.C(n_4469),
.Y(n_6115)
);

BUFx6f_ASAP7_75t_L g6116 ( 
.A(n_4547),
.Y(n_6116)
);

BUFx3_ASAP7_75t_L g6117 ( 
.A(n_5267),
.Y(n_6117)
);

AOI21xp5_ASAP7_75t_L g6118 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6118)
);

BUFx6f_ASAP7_75t_L g6119 ( 
.A(n_4547),
.Y(n_6119)
);

CKINVDCx8_ASAP7_75t_R g6120 ( 
.A(n_4486),
.Y(n_6120)
);

NOR2xp33_ASAP7_75t_L g6121 ( 
.A(n_4797),
.B(n_4817),
.Y(n_6121)
);

AOI22xp33_ASAP7_75t_L g6122 ( 
.A1(n_5001),
.A2(n_4553),
.B1(n_4699),
.B2(n_4688),
.Y(n_6122)
);

OAI22xp5_ASAP7_75t_L g6123 ( 
.A1(n_5292),
.A2(n_5209),
.B1(n_4817),
.B2(n_4797),
.Y(n_6123)
);

INVx5_ASAP7_75t_L g6124 ( 
.A(n_4568),
.Y(n_6124)
);

NAND2x1_ASAP7_75t_SL g6125 ( 
.A(n_5085),
.B(n_5149),
.Y(n_6125)
);

BUFx12f_ASAP7_75t_L g6126 ( 
.A(n_4703),
.Y(n_6126)
);

NOR2x1_ASAP7_75t_L g6127 ( 
.A(n_5331),
.B(n_5345),
.Y(n_6127)
);

O2A1O1Ixp33_ASAP7_75t_L g6128 ( 
.A1(n_5243),
.A2(n_5207),
.B(n_5259),
.C(n_5204),
.Y(n_6128)
);

AO22x1_ASAP7_75t_L g6129 ( 
.A1(n_5330),
.A2(n_5149),
.B1(n_4861),
.B2(n_4468),
.Y(n_6129)
);

BUFx12f_ASAP7_75t_L g6130 ( 
.A(n_4703),
.Y(n_6130)
);

AOI21xp5_ASAP7_75t_L g6131 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_4851),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_4851),
.Y(n_6133)
);

BUFx6f_ASAP7_75t_L g6134 ( 
.A(n_4547),
.Y(n_6134)
);

INVx1_ASAP7_75t_L g6135 ( 
.A(n_4851),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_4522),
.B(n_4524),
.Y(n_6136)
);

BUFx6f_ASAP7_75t_L g6137 ( 
.A(n_4547),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_4990),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_4524),
.B(n_4525),
.Y(n_6139)
);

OAI22xp5_ASAP7_75t_SL g6140 ( 
.A1(n_5387),
.A2(n_4599),
.B1(n_4698),
.B2(n_5377),
.Y(n_6140)
);

BUFx2_ASAP7_75t_L g6141 ( 
.A(n_5503),
.Y(n_6141)
);

NAND2xp5_ASAP7_75t_L g6142 ( 
.A(n_4525),
.B(n_4527),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_4858),
.Y(n_6143)
);

NAND2xp5_ASAP7_75t_L g6144 ( 
.A(n_4527),
.B(n_4530),
.Y(n_6144)
);

AOI22xp33_ASAP7_75t_L g6145 ( 
.A1(n_5001),
.A2(n_4553),
.B1(n_4688),
.B2(n_4648),
.Y(n_6145)
);

AOI21xp33_ASAP7_75t_L g6146 ( 
.A1(n_4469),
.A2(n_4482),
.B(n_4441),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_4858),
.Y(n_6147)
);

OR2x2_ASAP7_75t_L g6148 ( 
.A(n_5097),
.B(n_5355),
.Y(n_6148)
);

AOI22xp33_ASAP7_75t_L g6149 ( 
.A1(n_4648),
.A2(n_4736),
.B1(n_4802),
.B2(n_4749),
.Y(n_6149)
);

NOR2xp33_ASAP7_75t_L g6150 ( 
.A(n_4817),
.B(n_4736),
.Y(n_6150)
);

AOI22xp33_ASAP7_75t_SL g6151 ( 
.A1(n_5063),
.A2(n_5067),
.B1(n_4749),
.B2(n_4805),
.Y(n_6151)
);

CKINVDCx5p33_ASAP7_75t_R g6152 ( 
.A(n_4624),
.Y(n_6152)
);

NOR2xp67_ASAP7_75t_L g6153 ( 
.A(n_5215),
.B(n_5222),
.Y(n_6153)
);

INVx3_ASAP7_75t_L g6154 ( 
.A(n_4965),
.Y(n_6154)
);

NAND2xp5_ASAP7_75t_L g6155 ( 
.A(n_4530),
.B(n_4531),
.Y(n_6155)
);

O2A1O1Ixp5_ASAP7_75t_SL g6156 ( 
.A1(n_5182),
.A2(n_5189),
.B(n_4905),
.C(n_4908),
.Y(n_6156)
);

BUFx10_ASAP7_75t_L g6157 ( 
.A(n_4775),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_4858),
.Y(n_6158)
);

NOR2xp33_ASAP7_75t_L g6159 ( 
.A(n_4817),
.B(n_4802),
.Y(n_6159)
);

OAI22xp5_ASAP7_75t_L g6160 ( 
.A1(n_5209),
.A2(n_5181),
.B1(n_4634),
.B2(n_5334),
.Y(n_6160)
);

INVx4_ASAP7_75t_L g6161 ( 
.A(n_4885),
.Y(n_6161)
);

OAI22xp5_ASAP7_75t_L g6162 ( 
.A1(n_4634),
.A2(n_5334),
.B1(n_5067),
.B2(n_5063),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_L g6163 ( 
.A(n_4531),
.B(n_4533),
.Y(n_6163)
);

INVx3_ASAP7_75t_L g6164 ( 
.A(n_4965),
.Y(n_6164)
);

AOI21xp5_ASAP7_75t_L g6165 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6165)
);

AOI21xp5_ASAP7_75t_L g6166 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6166)
);

INVx4_ASAP7_75t_L g6167 ( 
.A(n_4948),
.Y(n_6167)
);

NOR2xp33_ASAP7_75t_L g6168 ( 
.A(n_4802),
.B(n_4805),
.Y(n_6168)
);

AOI22xp33_ASAP7_75t_SL g6169 ( 
.A1(n_4805),
.A2(n_4808),
.B1(n_4850),
.B2(n_4823),
.Y(n_6169)
);

OAI22xp5_ASAP7_75t_SL g6170 ( 
.A1(n_5387),
.A2(n_4599),
.B1(n_4698),
.B2(n_5377),
.Y(n_6170)
);

BUFx6f_ASAP7_75t_L g6171 ( 
.A(n_4547),
.Y(n_6171)
);

BUFx2_ASAP7_75t_SL g6172 ( 
.A(n_5372),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_4863),
.Y(n_6173)
);

BUFx2_ASAP7_75t_L g6174 ( 
.A(n_5503),
.Y(n_6174)
);

O2A1O1Ixp33_ASAP7_75t_L g6175 ( 
.A1(n_5204),
.A2(n_5207),
.B(n_5310),
.C(n_5259),
.Y(n_6175)
);

AOI21xp5_ASAP7_75t_L g6176 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_4863),
.Y(n_6177)
);

BUFx3_ASAP7_75t_L g6178 ( 
.A(n_5267),
.Y(n_6178)
);

NAND2xp5_ASAP7_75t_L g6179 ( 
.A(n_4533),
.B(n_4534),
.Y(n_6179)
);

AOI21xp5_ASAP7_75t_L g6180 ( 
.A1(n_4890),
.A2(n_5136),
.B(n_5034),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_L g6181 ( 
.A(n_4534),
.B(n_4537),
.Y(n_6181)
);

AOI22xp33_ASAP7_75t_L g6182 ( 
.A1(n_4808),
.A2(n_4850),
.B1(n_4855),
.B2(n_4823),
.Y(n_6182)
);

AOI22xp33_ASAP7_75t_L g6183 ( 
.A1(n_4808),
.A2(n_4850),
.B1(n_4855),
.B2(n_4823),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_4863),
.Y(n_6184)
);

OAI22xp5_ASAP7_75t_L g6185 ( 
.A1(n_5366),
.A2(n_5384),
.B1(n_5274),
.B2(n_4874),
.Y(n_6185)
);

BUFx12f_ASAP7_75t_L g6186 ( 
.A(n_4705),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_SL g6187 ( 
.A(n_5352),
.B(n_5370),
.Y(n_6187)
);

BUFx2_ASAP7_75t_SL g6188 ( 
.A(n_5372),
.Y(n_6188)
);

NOR2xp33_ASAP7_75t_L g6189 ( 
.A(n_4855),
.B(n_4874),
.Y(n_6189)
);

OR2x2_ASAP7_75t_L g6190 ( 
.A(n_5097),
.B(n_5355),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_4864),
.Y(n_6191)
);

BUFx6f_ASAP7_75t_L g6192 ( 
.A(n_4547),
.Y(n_6192)
);

INVxp67_ASAP7_75t_L g6193 ( 
.A(n_4964),
.Y(n_6193)
);

BUFx2_ASAP7_75t_L g6194 ( 
.A(n_5503),
.Y(n_6194)
);

NAND2xp5_ASAP7_75t_L g6195 ( 
.A(n_4537),
.B(n_4538),
.Y(n_6195)
);

BUFx6f_ASAP7_75t_L g6196 ( 
.A(n_4547),
.Y(n_6196)
);

BUFx6f_ASAP7_75t_L g6197 ( 
.A(n_4559),
.Y(n_6197)
);

NOR2xp33_ASAP7_75t_L g6198 ( 
.A(n_4874),
.B(n_4882),
.Y(n_6198)
);

AOI21xp5_ASAP7_75t_L g6199 ( 
.A1(n_5034),
.A2(n_5201),
.B(n_5136),
.Y(n_6199)
);

OAI21xp33_ASAP7_75t_L g6200 ( 
.A1(n_4433),
.A2(n_4441),
.B(n_4438),
.Y(n_6200)
);

OAI22xp5_ASAP7_75t_L g6201 ( 
.A1(n_5366),
.A2(n_5384),
.B1(n_5274),
.B2(n_4940),
.Y(n_6201)
);

NOR2xp33_ASAP7_75t_L g6202 ( 
.A(n_4882),
.B(n_4940),
.Y(n_6202)
);

AOI21xp5_ASAP7_75t_L g6203 ( 
.A1(n_5201),
.A2(n_5308),
.B(n_5286),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_4864),
.Y(n_6204)
);

OAI22xp5_ASAP7_75t_L g6205 ( 
.A1(n_4882),
.A2(n_4960),
.B1(n_4983),
.B2(n_4940),
.Y(n_6205)
);

NOR2xp33_ASAP7_75t_L g6206 ( 
.A(n_4960),
.B(n_4983),
.Y(n_6206)
);

CKINVDCx8_ASAP7_75t_R g6207 ( 
.A(n_4486),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_4864),
.Y(n_6208)
);

NAND2xp5_ASAP7_75t_SL g6209 ( 
.A(n_5370),
.B(n_4657),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_4867),
.Y(n_6210)
);

O2A1O1Ixp5_ASAP7_75t_L g6211 ( 
.A1(n_4493),
.A2(n_4526),
.B(n_5016),
.C(n_4846),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_4867),
.Y(n_6212)
);

BUFx2_ASAP7_75t_L g6213 ( 
.A(n_5503),
.Y(n_6213)
);

BUFx2_ASAP7_75t_L g6214 ( 
.A(n_5503),
.Y(n_6214)
);

INVx1_ASAP7_75t_SL g6215 ( 
.A(n_4801),
.Y(n_6215)
);

BUFx6f_ASAP7_75t_L g6216 ( 
.A(n_4559),
.Y(n_6216)
);

BUFx2_ASAP7_75t_L g6217 ( 
.A(n_5503),
.Y(n_6217)
);

OAI22xp33_ASAP7_75t_L g6218 ( 
.A1(n_5435),
.A2(n_5248),
.B1(n_5269),
.B2(n_5526),
.Y(n_6218)
);

HAxp5_ASAP7_75t_L g6219 ( 
.A(n_4449),
.B(n_4526),
.CON(n_6219),
.SN(n_6219)
);

NAND2xp5_ASAP7_75t_SL g6220 ( 
.A(n_4657),
.B(n_5451),
.Y(n_6220)
);

NOR2xp33_ASAP7_75t_L g6221 ( 
.A(n_4960),
.B(n_4983),
.Y(n_6221)
);

BUFx2_ASAP7_75t_L g6222 ( 
.A(n_5518),
.Y(n_6222)
);

BUFx2_ASAP7_75t_L g6223 ( 
.A(n_5518),
.Y(n_6223)
);

O2A1O1Ixp33_ASAP7_75t_L g6224 ( 
.A1(n_5310),
.A2(n_5343),
.B(n_5491),
.C(n_5404),
.Y(n_6224)
);

AOI21xp5_ASAP7_75t_L g6225 ( 
.A1(n_5201),
.A2(n_5308),
.B(n_5286),
.Y(n_6225)
);

AOI22xp33_ASAP7_75t_SL g6226 ( 
.A1(n_4989),
.A2(n_5051),
.B1(n_5089),
.B2(n_5277),
.Y(n_6226)
);

AOI22xp5_ASAP7_75t_L g6227 ( 
.A1(n_4989),
.A2(n_5089),
.B1(n_5051),
.B2(n_5454),
.Y(n_6227)
);

INVx3_ASAP7_75t_L g6228 ( 
.A(n_4980),
.Y(n_6228)
);

OAI22x1_ASAP7_75t_L g6229 ( 
.A1(n_5069),
.A2(n_5097),
.B1(n_4964),
.B2(n_4998),
.Y(n_6229)
);

NOR2xp33_ASAP7_75t_L g6230 ( 
.A(n_4989),
.B(n_5051),
.Y(n_6230)
);

NOR2xp33_ASAP7_75t_L g6231 ( 
.A(n_5089),
.B(n_5526),
.Y(n_6231)
);

BUFx2_ASAP7_75t_L g6232 ( 
.A(n_5518),
.Y(n_6232)
);

BUFx3_ASAP7_75t_L g6233 ( 
.A(n_5267),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_4867),
.Y(n_6234)
);

CKINVDCx20_ASAP7_75t_R g6235 ( 
.A(n_5306),
.Y(n_6235)
);

BUFx6f_ASAP7_75t_L g6236 ( 
.A(n_4559),
.Y(n_6236)
);

AOI21x1_ASAP7_75t_L g6237 ( 
.A1(n_4941),
.A2(n_4943),
.B(n_5182),
.Y(n_6237)
);

AOI21xp5_ASAP7_75t_L g6238 ( 
.A1(n_5201),
.A2(n_5308),
.B(n_5286),
.Y(n_6238)
);

NAND2x1p5_ASAP7_75t_L g6239 ( 
.A(n_4523),
.B(n_4709),
.Y(n_6239)
);

BUFx2_ASAP7_75t_L g6240 ( 
.A(n_5518),
.Y(n_6240)
);

BUFx4f_ASAP7_75t_L g6241 ( 
.A(n_5206),
.Y(n_6241)
);

OR2x6_ASAP7_75t_L g6242 ( 
.A(n_5518),
.B(n_5401),
.Y(n_6242)
);

NAND2xp5_ASAP7_75t_L g6243 ( 
.A(n_4538),
.B(n_4539),
.Y(n_6243)
);

NAND2xp5_ASAP7_75t_SL g6244 ( 
.A(n_5451),
.B(n_4979),
.Y(n_6244)
);

NOR2xp33_ASAP7_75t_L g6245 ( 
.A(n_5491),
.B(n_4539),
.Y(n_6245)
);

BUFx12f_ASAP7_75t_L g6246 ( 
.A(n_4705),
.Y(n_6246)
);

NOR2xp33_ASAP7_75t_L g6247 ( 
.A(n_4540),
.B(n_4548),
.Y(n_6247)
);

INVx4_ASAP7_75t_L g6248 ( 
.A(n_4885),
.Y(n_6248)
);

BUFx4f_ASAP7_75t_L g6249 ( 
.A(n_5206),
.Y(n_6249)
);

AOI21xp5_ASAP7_75t_L g6250 ( 
.A1(n_5201),
.A2(n_5308),
.B(n_5286),
.Y(n_6250)
);

O2A1O1Ixp33_ASAP7_75t_L g6251 ( 
.A1(n_5343),
.A2(n_5404),
.B(n_5402),
.C(n_5528),
.Y(n_6251)
);

BUFx6f_ASAP7_75t_L g6252 ( 
.A(n_4559),
.Y(n_6252)
);

OAI22xp5_ASAP7_75t_L g6253 ( 
.A1(n_5178),
.A2(n_5186),
.B1(n_5188),
.B2(n_5183),
.Y(n_6253)
);

OAI22xp5_ASAP7_75t_L g6254 ( 
.A1(n_5178),
.A2(n_5186),
.B1(n_5188),
.B2(n_5183),
.Y(n_6254)
);

NOR2xp33_ASAP7_75t_L g6255 ( 
.A(n_4540),
.B(n_4548),
.Y(n_6255)
);

BUFx2_ASAP7_75t_L g6256 ( 
.A(n_5518),
.Y(n_6256)
);

INVx5_ASAP7_75t_L g6257 ( 
.A(n_4568),
.Y(n_6257)
);

O2A1O1Ixp33_ASAP7_75t_L g6258 ( 
.A1(n_5402),
.A2(n_5528),
.B(n_5349),
.C(n_5485),
.Y(n_6258)
);

INVx3_ASAP7_75t_L g6259 ( 
.A(n_4980),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_4873),
.Y(n_6260)
);

CKINVDCx5p33_ASAP7_75t_R g6261 ( 
.A(n_4724),
.Y(n_6261)
);

AOI22xp33_ASAP7_75t_SL g6262 ( 
.A1(n_5277),
.A2(n_5069),
.B1(n_4640),
.B2(n_4979),
.Y(n_6262)
);

CKINVDCx11_ASAP7_75t_R g6263 ( 
.A(n_4494),
.Y(n_6263)
);

NOR2xp33_ASAP7_75t_L g6264 ( 
.A(n_4549),
.B(n_4562),
.Y(n_6264)
);

BUFx2_ASAP7_75t_L g6265 ( 
.A(n_5518),
.Y(n_6265)
);

OAI22xp5_ASAP7_75t_L g6266 ( 
.A1(n_5196),
.A2(n_5208),
.B1(n_5225),
.B2(n_5200),
.Y(n_6266)
);

OR2x6_ASAP7_75t_L g6267 ( 
.A(n_5401),
.B(n_5201),
.Y(n_6267)
);

BUFx6f_ASAP7_75t_L g6268 ( 
.A(n_4559),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_4873),
.Y(n_6269)
);

BUFx2_ASAP7_75t_L g6270 ( 
.A(n_5069),
.Y(n_6270)
);

AOI22xp33_ASAP7_75t_L g6271 ( 
.A1(n_5248),
.A2(n_5454),
.B1(n_5128),
.B2(n_5126),
.Y(n_6271)
);

CKINVDCx20_ASAP7_75t_R g6272 ( 
.A(n_5450),
.Y(n_6272)
);

INVx5_ASAP7_75t_L g6273 ( 
.A(n_4568),
.Y(n_6273)
);

CKINVDCx5p33_ASAP7_75t_R g6274 ( 
.A(n_5488),
.Y(n_6274)
);

NOR2xp33_ASAP7_75t_L g6275 ( 
.A(n_4549),
.B(n_4562),
.Y(n_6275)
);

NAND2xp5_ASAP7_75t_L g6276 ( 
.A(n_4565),
.B(n_4566),
.Y(n_6276)
);

OAI22xp5_ASAP7_75t_SL g6277 ( 
.A1(n_4599),
.A2(n_4698),
.B1(n_5450),
.B2(n_5476),
.Y(n_6277)
);

OAI22xp5_ASAP7_75t_SL g6278 ( 
.A1(n_5476),
.A2(n_5316),
.B1(n_5435),
.B2(n_5213),
.Y(n_6278)
);

OAI22xp5_ASAP7_75t_L g6279 ( 
.A1(n_5196),
.A2(n_5208),
.B1(n_5225),
.B2(n_5200),
.Y(n_6279)
);

INVx3_ASAP7_75t_L g6280 ( 
.A(n_4980),
.Y(n_6280)
);

OAI21x1_ASAP7_75t_SL g6281 ( 
.A1(n_5349),
.A2(n_5052),
.B(n_5049),
.Y(n_6281)
);

BUFx8_ASAP7_75t_SL g6282 ( 
.A(n_4494),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_4873),
.Y(n_6283)
);

O2A1O1Ixp33_ASAP7_75t_L g6284 ( 
.A1(n_5485),
.A2(n_4458),
.B(n_4442),
.C(n_4438),
.Y(n_6284)
);

OAI21xp5_ASAP7_75t_L g6285 ( 
.A1(n_4901),
.A2(n_4896),
.B(n_4856),
.Y(n_6285)
);

AOI22xp5_ASAP7_75t_L g6286 ( 
.A1(n_4846),
.A2(n_5016),
.B1(n_5213),
.B2(n_5128),
.Y(n_6286)
);

OAI22xp5_ASAP7_75t_L g6287 ( 
.A1(n_5227),
.A2(n_5232),
.B1(n_5235),
.B2(n_5234),
.Y(n_6287)
);

A2O1A1Ixp33_ASAP7_75t_L g6288 ( 
.A1(n_4979),
.A2(n_5012),
.B(n_5015),
.C(n_4998),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_4876),
.Y(n_6289)
);

AND2x2_ASAP7_75t_L g6290 ( 
.A(n_4434),
.B(n_4971),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_4876),
.Y(n_6291)
);

A2O1A1Ixp33_ASAP7_75t_L g6292 ( 
.A1(n_4998),
.A2(n_5015),
.B(n_5017),
.C(n_5012),
.Y(n_6292)
);

O2A1O1Ixp33_ASAP7_75t_L g6293 ( 
.A1(n_4447),
.A2(n_4442),
.B(n_4450),
.C(n_4433),
.Y(n_6293)
);

AOI22xp33_ASAP7_75t_L g6294 ( 
.A1(n_5126),
.A2(n_5444),
.B1(n_5344),
.B2(n_5383),
.Y(n_6294)
);

NAND2xp5_ASAP7_75t_L g6295 ( 
.A(n_4565),
.B(n_4566),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_4434),
.B(n_4971),
.Y(n_6296)
);

O2A1O1Ixp5_ASAP7_75t_SL g6297 ( 
.A1(n_5182),
.A2(n_5189),
.B(n_4907),
.C(n_4908),
.Y(n_6297)
);

A2O1A1Ixp33_ASAP7_75t_L g6298 ( 
.A1(n_5012),
.A2(n_5017),
.B(n_5056),
.C(n_5015),
.Y(n_6298)
);

NAND2xp5_ASAP7_75t_L g6299 ( 
.A(n_4569),
.B(n_4575),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_4876),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_4879),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_4879),
.Y(n_6302)
);

NOR2xp33_ASAP7_75t_L g6303 ( 
.A(n_4569),
.B(n_4575),
.Y(n_6303)
);

NOR2xp33_ASAP7_75t_L g6304 ( 
.A(n_4577),
.B(n_4587),
.Y(n_6304)
);

A2O1A1Ixp33_ASAP7_75t_SL g6305 ( 
.A1(n_5515),
.A2(n_5436),
.B(n_5432),
.C(n_5344),
.Y(n_6305)
);

CKINVDCx5p33_ASAP7_75t_R g6306 ( 
.A(n_5488),
.Y(n_6306)
);

BUFx2_ASAP7_75t_L g6307 ( 
.A(n_5401),
.Y(n_6307)
);

OR2x2_ASAP7_75t_L g6308 ( 
.A(n_5355),
.B(n_4427),
.Y(n_6308)
);

NAND3xp33_ASAP7_75t_L g6309 ( 
.A(n_5515),
.B(n_5408),
.C(n_4896),
.Y(n_6309)
);

BUFx6f_ASAP7_75t_L g6310 ( 
.A(n_4559),
.Y(n_6310)
);

OAI22xp5_ASAP7_75t_L g6311 ( 
.A1(n_5227),
.A2(n_5234),
.B1(n_5235),
.B2(n_5232),
.Y(n_6311)
);

NAND2xp5_ASAP7_75t_L g6312 ( 
.A(n_4577),
.B(n_4587),
.Y(n_6312)
);

OAI22xp5_ASAP7_75t_L g6313 ( 
.A1(n_5240),
.A2(n_5246),
.B1(n_5253),
.B2(n_5245),
.Y(n_6313)
);

HB1xp67_ASAP7_75t_L g6314 ( 
.A(n_4719),
.Y(n_6314)
);

INVx3_ASAP7_75t_L g6315 ( 
.A(n_4980),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_4879),
.Y(n_6316)
);

O2A1O1Ixp33_ASAP7_75t_L g6317 ( 
.A1(n_4447),
.A2(n_4450),
.B(n_4458),
.C(n_4453),
.Y(n_6317)
);

O2A1O1Ixp33_ASAP7_75t_SL g6318 ( 
.A1(n_4453),
.A2(n_4459),
.B(n_4467),
.C(n_5417),
.Y(n_6318)
);

NAND2xp5_ASAP7_75t_L g6319 ( 
.A(n_4589),
.B(n_4591),
.Y(n_6319)
);

BUFx12f_ASAP7_75t_L g6320 ( 
.A(n_4708),
.Y(n_6320)
);

AND2x2_ASAP7_75t_L g6321 ( 
.A(n_4434),
.B(n_5070),
.Y(n_6321)
);

HB1xp67_ASAP7_75t_L g6322 ( 
.A(n_4719),
.Y(n_6322)
);

O2A1O1Ixp33_ASAP7_75t_L g6323 ( 
.A1(n_4459),
.A2(n_4467),
.B(n_5253),
.C(n_5245),
.Y(n_6323)
);

A2O1A1Ixp33_ASAP7_75t_L g6324 ( 
.A1(n_5017),
.A2(n_5056),
.B(n_4901),
.C(n_4856),
.Y(n_6324)
);

INVx3_ASAP7_75t_L g6325 ( 
.A(n_4980),
.Y(n_6325)
);

BUFx3_ASAP7_75t_L g6326 ( 
.A(n_5279),
.Y(n_6326)
);

INVx3_ASAP7_75t_L g6327 ( 
.A(n_4980),
.Y(n_6327)
);

BUFx3_ASAP7_75t_L g6328 ( 
.A(n_5279),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_SL g6329 ( 
.A(n_5056),
.B(n_4961),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_4880),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_4880),
.Y(n_6331)
);

NOR2xp33_ASAP7_75t_L g6332 ( 
.A(n_4589),
.B(n_4591),
.Y(n_6332)
);

NAND2xp5_ASAP7_75t_L g6333 ( 
.A(n_4595),
.B(n_4596),
.Y(n_6333)
);

BUFx3_ASAP7_75t_L g6334 ( 
.A(n_5279),
.Y(n_6334)
);

NAND2xp5_ASAP7_75t_L g6335 ( 
.A(n_4595),
.B(n_4596),
.Y(n_6335)
);

BUFx3_ASAP7_75t_L g6336 ( 
.A(n_5279),
.Y(n_6336)
);

NAND3xp33_ASAP7_75t_L g6337 ( 
.A(n_5151),
.B(n_5339),
.C(n_5220),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_4880),
.Y(n_6338)
);

NOR2xp33_ASAP7_75t_L g6339 ( 
.A(n_4602),
.B(n_4603),
.Y(n_6339)
);

BUFx3_ASAP7_75t_L g6340 ( 
.A(n_5293),
.Y(n_6340)
);

AOI21xp5_ASAP7_75t_L g6341 ( 
.A1(n_5201),
.A2(n_5308),
.B(n_5286),
.Y(n_6341)
);

INVx4_ASAP7_75t_L g6342 ( 
.A(n_4885),
.Y(n_6342)
);

HB1xp67_ASAP7_75t_L g6343 ( 
.A(n_4733),
.Y(n_6343)
);

HB1xp67_ASAP7_75t_L g6344 ( 
.A(n_4733),
.Y(n_6344)
);

OAI22xp5_ASAP7_75t_SL g6345 ( 
.A1(n_5316),
.A2(n_4861),
.B1(n_4468),
.B2(n_5524),
.Y(n_6345)
);

A2O1A1Ixp33_ASAP7_75t_L g6346 ( 
.A1(n_5172),
.A2(n_5218),
.B(n_5087),
.C(n_5356),
.Y(n_6346)
);

NAND2x1p5_ASAP7_75t_L g6347 ( 
.A(n_4523),
.B(n_4709),
.Y(n_6347)
);

HB1xp67_ASAP7_75t_L g6348 ( 
.A(n_4743),
.Y(n_6348)
);

NAND2xp5_ASAP7_75t_L g6349 ( 
.A(n_4602),
.B(n_4603),
.Y(n_6349)
);

BUFx3_ASAP7_75t_L g6350 ( 
.A(n_5293),
.Y(n_6350)
);

O2A1O1Ixp33_ASAP7_75t_L g6351 ( 
.A1(n_5257),
.A2(n_5284),
.B(n_5301),
.C(n_5270),
.Y(n_6351)
);

AOI21xp5_ASAP7_75t_L g6352 ( 
.A1(n_5286),
.A2(n_5317),
.B(n_5308),
.Y(n_6352)
);

CKINVDCx8_ASAP7_75t_R g6353 ( 
.A(n_4885),
.Y(n_6353)
);

NOR2xp33_ASAP7_75t_L g6354 ( 
.A(n_4605),
.B(n_4607),
.Y(n_6354)
);

NAND2xp5_ASAP7_75t_SL g6355 ( 
.A(n_4961),
.B(n_4969),
.Y(n_6355)
);

O2A1O1Ixp33_ASAP7_75t_L g6356 ( 
.A1(n_5246),
.A2(n_5302),
.B(n_5261),
.C(n_5240),
.Y(n_6356)
);

O2A1O1Ixp33_ASAP7_75t_L g6357 ( 
.A1(n_5254),
.A2(n_5255),
.B(n_5278),
.C(n_5257),
.Y(n_6357)
);

BUFx4f_ASAP7_75t_SL g6358 ( 
.A(n_4494),
.Y(n_6358)
);

OAI22xp33_ASAP7_75t_L g6359 ( 
.A1(n_5269),
.A2(n_5479),
.B1(n_5511),
.B2(n_5283),
.Y(n_6359)
);

CKINVDCx5p33_ASAP7_75t_R g6360 ( 
.A(n_5522),
.Y(n_6360)
);

BUFx2_ASAP7_75t_L g6361 ( 
.A(n_5401),
.Y(n_6361)
);

OAI22xp5_ASAP7_75t_L g6362 ( 
.A1(n_5254),
.A2(n_5256),
.B1(n_5261),
.B2(n_5255),
.Y(n_6362)
);

NAND2xp5_ASAP7_75t_SL g6363 ( 
.A(n_4961),
.B(n_4969),
.Y(n_6363)
);

AOI22xp33_ASAP7_75t_L g6364 ( 
.A1(n_5444),
.A2(n_5373),
.B1(n_5383),
.B2(n_5283),
.Y(n_6364)
);

NOR2xp33_ASAP7_75t_L g6365 ( 
.A(n_4605),
.B(n_4607),
.Y(n_6365)
);

AOI21xp33_ASAP7_75t_L g6366 ( 
.A1(n_5356),
.A2(n_5346),
.B(n_4430),
.Y(n_6366)
);

AOI22x1_ASAP7_75t_L g6367 ( 
.A1(n_5047),
.A2(n_5218),
.B1(n_5172),
.B2(n_5524),
.Y(n_6367)
);

AOI21xp5_ASAP7_75t_L g6368 ( 
.A1(n_5286),
.A2(n_5317),
.B(n_5308),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_4611),
.B(n_4617),
.Y(n_6369)
);

O2A1O1Ixp33_ASAP7_75t_L g6370 ( 
.A1(n_5276),
.A2(n_5319),
.B(n_5278),
.C(n_5256),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_4611),
.B(n_4617),
.Y(n_6371)
);

A2O1A1Ixp33_ASAP7_75t_L g6372 ( 
.A1(n_5172),
.A2(n_5218),
.B(n_5087),
.C(n_5511),
.Y(n_6372)
);

INVx4_ASAP7_75t_L g6373 ( 
.A(n_4885),
.Y(n_6373)
);

HB1xp67_ASAP7_75t_L g6374 ( 
.A(n_4743),
.Y(n_6374)
);

BUFx2_ASAP7_75t_L g6375 ( 
.A(n_5401),
.Y(n_6375)
);

A2O1A1Ixp33_ASAP7_75t_SL g6376 ( 
.A1(n_5432),
.A2(n_5436),
.B(n_5373),
.C(n_5426),
.Y(n_6376)
);

NOR2xp33_ASAP7_75t_L g6377 ( 
.A(n_4619),
.B(n_4620),
.Y(n_6377)
);

OR2x2_ASAP7_75t_L g6378 ( 
.A(n_4427),
.B(n_4430),
.Y(n_6378)
);

AO32x2_ASAP7_75t_L g6379 ( 
.A1(n_4710),
.A2(n_4932),
.A3(n_4927),
.B1(n_4871),
.B2(n_4866),
.Y(n_6379)
);

AOI22xp33_ASAP7_75t_L g6380 ( 
.A1(n_5283),
.A2(n_4944),
.B1(n_5000),
.B2(n_4723),
.Y(n_6380)
);

INVx4_ASAP7_75t_L g6381 ( 
.A(n_4885),
.Y(n_6381)
);

AOI22xp33_ASAP7_75t_L g6382 ( 
.A1(n_4723),
.A2(n_5000),
.B1(n_5084),
.B2(n_4944),
.Y(n_6382)
);

BUFx6f_ASAP7_75t_L g6383 ( 
.A(n_4568),
.Y(n_6383)
);

AOI21xp5_ASAP7_75t_L g6384 ( 
.A1(n_5317),
.A2(n_5338),
.B(n_5318),
.Y(n_6384)
);

OAI22xp5_ASAP7_75t_L g6385 ( 
.A1(n_5270),
.A2(n_5276),
.B1(n_5284),
.B2(n_5272),
.Y(n_6385)
);

INVx3_ASAP7_75t_L g6386 ( 
.A(n_5004),
.Y(n_6386)
);

BUFx2_ASAP7_75t_L g6387 ( 
.A(n_5401),
.Y(n_6387)
);

NAND2xp5_ASAP7_75t_L g6388 ( 
.A(n_4619),
.B(n_4620),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_L g6389 ( 
.A(n_4639),
.B(n_4641),
.Y(n_6389)
);

O2A1O1Ixp33_ASAP7_75t_L g6390 ( 
.A1(n_5302),
.A2(n_5328),
.B(n_5272),
.C(n_5312),
.Y(n_6390)
);

BUFx2_ASAP7_75t_L g6391 ( 
.A(n_5401),
.Y(n_6391)
);

NOR3x1_ASAP7_75t_L g6392 ( 
.A(n_5301),
.B(n_5319),
.C(n_5312),
.Y(n_6392)
);

INVx4_ASAP7_75t_L g6393 ( 
.A(n_4885),
.Y(n_6393)
);

NAND2xp5_ASAP7_75t_SL g6394 ( 
.A(n_4961),
.B(n_4969),
.Y(n_6394)
);

BUFx2_ASAP7_75t_L g6395 ( 
.A(n_4545),
.Y(n_6395)
);

INVxp67_ASAP7_75t_L g6396 ( 
.A(n_5224),
.Y(n_6396)
);

INVx1_ASAP7_75t_SL g6397 ( 
.A(n_4801),
.Y(n_6397)
);

AOI21xp5_ASAP7_75t_L g6398 ( 
.A1(n_5317),
.A2(n_5338),
.B(n_5318),
.Y(n_6398)
);

NAND2xp5_ASAP7_75t_L g6399 ( 
.A(n_4639),
.B(n_4641),
.Y(n_6399)
);

BUFx3_ASAP7_75t_L g6400 ( 
.A(n_5293),
.Y(n_6400)
);

A2O1A1Ixp33_ASAP7_75t_L g6401 ( 
.A1(n_5087),
.A2(n_4969),
.B(n_4640),
.C(n_5320),
.Y(n_6401)
);

BUFx6f_ASAP7_75t_L g6402 ( 
.A(n_4568),
.Y(n_6402)
);

BUFx12f_ASAP7_75t_L g6403 ( 
.A(n_4708),
.Y(n_6403)
);

NOR2xp33_ASAP7_75t_L g6404 ( 
.A(n_4646),
.B(n_4649),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_4646),
.B(n_4649),
.Y(n_6405)
);

CKINVDCx5p33_ASAP7_75t_R g6406 ( 
.A(n_5522),
.Y(n_6406)
);

BUFx2_ASAP7_75t_L g6407 ( 
.A(n_4545),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_4656),
.B(n_4658),
.Y(n_6408)
);

AND2x6_ASAP7_75t_L g6409 ( 
.A(n_5206),
.B(n_5229),
.Y(n_6409)
);

OR2x6_ASAP7_75t_L g6410 ( 
.A(n_5317),
.B(n_5318),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_5145),
.B(n_4466),
.Y(n_6411)
);

AOI21xp5_ASAP7_75t_L g6412 ( 
.A1(n_5317),
.A2(n_5338),
.B(n_5318),
.Y(n_6412)
);

NAND2xp5_ASAP7_75t_L g6413 ( 
.A(n_4656),
.B(n_4658),
.Y(n_6413)
);

NAND2x1_ASAP7_75t_SL g6414 ( 
.A(n_4917),
.B(n_4919),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_4666),
.B(n_4670),
.Y(n_6415)
);

A2O1A1Ixp33_ASAP7_75t_SL g6416 ( 
.A1(n_5409),
.A2(n_5427),
.B(n_5430),
.C(n_5426),
.Y(n_6416)
);

AOI21xp33_ASAP7_75t_L g6417 ( 
.A1(n_5346),
.A2(n_5412),
.B(n_5406),
.Y(n_6417)
);

NAND2x1p5_ASAP7_75t_L g6418 ( 
.A(n_4709),
.B(n_4885),
.Y(n_6418)
);

BUFx3_ASAP7_75t_L g6419 ( 
.A(n_5293),
.Y(n_6419)
);

OR2x2_ASAP7_75t_L g6420 ( 
.A(n_4917),
.B(n_4919),
.Y(n_6420)
);

NOR2xp33_ASAP7_75t_L g6421 ( 
.A(n_4666),
.B(n_4670),
.Y(n_6421)
);

AOI21xp5_ASAP7_75t_L g6422 ( 
.A1(n_5317),
.A2(n_5338),
.B(n_5318),
.Y(n_6422)
);

OAI21xp5_ASAP7_75t_L g6423 ( 
.A1(n_5047),
.A2(n_5439),
.B(n_5478),
.Y(n_6423)
);

AOI22xp5_ASAP7_75t_L g6424 ( 
.A1(n_5473),
.A2(n_5445),
.B1(n_5516),
.B2(n_5469),
.Y(n_6424)
);

BUFx12f_ASAP7_75t_L g6425 ( 
.A(n_4843),
.Y(n_6425)
);

AOI22xp33_ASAP7_75t_L g6426 ( 
.A1(n_4723),
.A2(n_5000),
.B1(n_5084),
.B2(n_4944),
.Y(n_6426)
);

O2A1O1Ixp33_ASAP7_75t_L g6427 ( 
.A1(n_5320),
.A2(n_5328),
.B(n_5329),
.C(n_5047),
.Y(n_6427)
);

CKINVDCx5p33_ASAP7_75t_R g6428 ( 
.A(n_4494),
.Y(n_6428)
);

OR2x2_ASAP7_75t_L g6429 ( 
.A(n_4930),
.B(n_5020),
.Y(n_6429)
);

A2O1A1Ixp33_ASAP7_75t_L g6430 ( 
.A1(n_5087),
.A2(n_4640),
.B(n_5329),
.C(n_5530),
.Y(n_6430)
);

AOI22xp33_ASAP7_75t_L g6431 ( 
.A1(n_4944),
.A2(n_5084),
.B1(n_5160),
.B2(n_5000),
.Y(n_6431)
);

BUFx6f_ASAP7_75t_L g6432 ( 
.A(n_4571),
.Y(n_6432)
);

AOI21xp5_ASAP7_75t_L g6433 ( 
.A1(n_5318),
.A2(n_5338),
.B(n_5144),
.Y(n_6433)
);

NAND2xp5_ASAP7_75t_SL g6434 ( 
.A(n_5479),
.B(n_5364),
.Y(n_6434)
);

BUFx3_ASAP7_75t_L g6435 ( 
.A(n_5299),
.Y(n_6435)
);

INVx3_ASAP7_75t_L g6436 ( 
.A(n_5004),
.Y(n_6436)
);

INVx3_ASAP7_75t_L g6437 ( 
.A(n_5004),
.Y(n_6437)
);

NAND2xp5_ASAP7_75t_L g6438 ( 
.A(n_4671),
.B(n_4676),
.Y(n_6438)
);

AOI22xp5_ASAP7_75t_L g6439 ( 
.A1(n_5473),
.A2(n_5445),
.B1(n_5516),
.B2(n_5469),
.Y(n_6439)
);

AOI21xp5_ASAP7_75t_L g6440 ( 
.A1(n_5318),
.A2(n_5338),
.B(n_5144),
.Y(n_6440)
);

INVx3_ASAP7_75t_L g6441 ( 
.A(n_5004),
.Y(n_6441)
);

AOI21xp5_ASAP7_75t_L g6442 ( 
.A1(n_5338),
.A2(n_5144),
.B(n_4542),
.Y(n_6442)
);

INVxp67_ASAP7_75t_L g6443 ( 
.A(n_5224),
.Y(n_6443)
);

A2O1A1Ixp33_ASAP7_75t_L g6444 ( 
.A1(n_5087),
.A2(n_4640),
.B(n_5530),
.C(n_5413),
.Y(n_6444)
);

BUFx4_ASAP7_75t_SL g6445 ( 
.A(n_4843),
.Y(n_6445)
);

INVx1_ASAP7_75t_SL g6446 ( 
.A(n_4847),
.Y(n_6446)
);

NOR2xp33_ASAP7_75t_SL g6447 ( 
.A(n_4557),
.B(n_5380),
.Y(n_6447)
);

NOR2xp33_ASAP7_75t_L g6448 ( 
.A(n_4671),
.B(n_4676),
.Y(n_6448)
);

AND2x4_ASAP7_75t_L g6449 ( 
.A(n_4780),
.B(n_4820),
.Y(n_6449)
);

AOI33xp33_ASAP7_75t_L g6450 ( 
.A1(n_5509),
.A2(n_5521),
.A3(n_4903),
.B1(n_4870),
.B2(n_4847),
.B3(n_5507),
.Y(n_6450)
);

AOI22xp33_ASAP7_75t_L g6451 ( 
.A1(n_5084),
.A2(n_5160),
.B1(n_4468),
.B2(n_4861),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_L g6452 ( 
.A(n_4678),
.B(n_4681),
.Y(n_6452)
);

OR2x6_ASAP7_75t_L g6453 ( 
.A(n_5092),
.B(n_5359),
.Y(n_6453)
);

O2A1O1Ixp33_ASAP7_75t_L g6454 ( 
.A1(n_5047),
.A2(n_5439),
.B(n_5433),
.C(n_5143),
.Y(n_6454)
);

OAI22xp5_ASAP7_75t_L g6455 ( 
.A1(n_4678),
.A2(n_4682),
.B1(n_4685),
.B2(n_4681),
.Y(n_6455)
);

BUFx3_ASAP7_75t_L g6456 ( 
.A(n_5299),
.Y(n_6456)
);

AOI22xp5_ASAP7_75t_L g6457 ( 
.A1(n_5507),
.A2(n_4468),
.B1(n_4861),
.B2(n_5046),
.Y(n_6457)
);

BUFx8_ASAP7_75t_SL g6458 ( 
.A(n_4572),
.Y(n_6458)
);

BUFx3_ASAP7_75t_L g6459 ( 
.A(n_5299),
.Y(n_6459)
);

NAND2xp5_ASAP7_75t_L g6460 ( 
.A(n_4682),
.B(n_4685),
.Y(n_6460)
);

INVx4_ASAP7_75t_L g6461 ( 
.A(n_4948),
.Y(n_6461)
);

NOR2xp33_ASAP7_75t_L g6462 ( 
.A(n_4690),
.B(n_4694),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_4690),
.B(n_4694),
.Y(n_6463)
);

BUFx2_ASAP7_75t_L g6464 ( 
.A(n_4545),
.Y(n_6464)
);

NAND3xp33_ASAP7_75t_L g6465 ( 
.A(n_5151),
.B(n_5220),
.C(n_5339),
.Y(n_6465)
);

OAI22xp5_ASAP7_75t_L g6466 ( 
.A1(n_4696),
.A2(n_4707),
.B1(n_4711),
.B2(n_4706),
.Y(n_6466)
);

OR2x6_ASAP7_75t_L g6467 ( 
.A(n_5092),
.B(n_5359),
.Y(n_6467)
);

AOI21xp5_ASAP7_75t_L g6468 ( 
.A1(n_4542),
.A2(n_5144),
.B(n_5358),
.Y(n_6468)
);

OR2x2_ASAP7_75t_L g6469 ( 
.A(n_4930),
.B(n_5020),
.Y(n_6469)
);

AOI22xp33_ASAP7_75t_L g6470 ( 
.A1(n_5160),
.A2(n_5110),
.B1(n_5433),
.B2(n_4572),
.Y(n_6470)
);

AOI22xp33_ASAP7_75t_L g6471 ( 
.A1(n_5160),
.A2(n_5110),
.B1(n_4572),
.B2(n_5410),
.Y(n_6471)
);

INVx3_ASAP7_75t_L g6472 ( 
.A(n_5005),
.Y(n_6472)
);

NAND2xp33_ASAP7_75t_L g6473 ( 
.A(n_4463),
.B(n_4865),
.Y(n_6473)
);

INVx4_ASAP7_75t_L g6474 ( 
.A(n_4948),
.Y(n_6474)
);

BUFx2_ASAP7_75t_L g6475 ( 
.A(n_4560),
.Y(n_6475)
);

INVxp67_ASAP7_75t_SL g6476 ( 
.A(n_5035),
.Y(n_6476)
);

NAND2xp5_ASAP7_75t_L g6477 ( 
.A(n_4696),
.B(n_4706),
.Y(n_6477)
);

OAI22xp5_ASAP7_75t_L g6478 ( 
.A1(n_4707),
.A2(n_4716),
.B1(n_4721),
.B2(n_4711),
.Y(n_6478)
);

AOI21xp5_ASAP7_75t_L g6479 ( 
.A1(n_4542),
.A2(n_5144),
.B(n_5358),
.Y(n_6479)
);

INVx3_ASAP7_75t_L g6480 ( 
.A(n_5005),
.Y(n_6480)
);

INVx4_ASAP7_75t_L g6481 ( 
.A(n_4986),
.Y(n_6481)
);

AOI22x1_ASAP7_75t_L g6482 ( 
.A1(n_5047),
.A2(n_5524),
.B1(n_5117),
.B2(n_5121),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_L g6483 ( 
.A(n_4716),
.B(n_4721),
.Y(n_6483)
);

INVx3_ASAP7_75t_L g6484 ( 
.A(n_5005),
.Y(n_6484)
);

INVx3_ASAP7_75t_L g6485 ( 
.A(n_5005),
.Y(n_6485)
);

AOI21x1_ASAP7_75t_L g6486 ( 
.A1(n_4941),
.A2(n_4943),
.B(n_5192),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_L g6487 ( 
.A(n_4725),
.B(n_4726),
.Y(n_6487)
);

INVxp67_ASAP7_75t_L g6488 ( 
.A(n_5224),
.Y(n_6488)
);

NAND2xp5_ASAP7_75t_L g6489 ( 
.A(n_4725),
.B(n_4726),
.Y(n_6489)
);

CKINVDCx8_ASAP7_75t_R g6490 ( 
.A(n_4948),
.Y(n_6490)
);

CKINVDCx8_ASAP7_75t_R g6491 ( 
.A(n_4948),
.Y(n_6491)
);

NAND2xp5_ASAP7_75t_L g6492 ( 
.A(n_4728),
.B(n_4734),
.Y(n_6492)
);

OAI22xp33_ASAP7_75t_L g6493 ( 
.A1(n_4557),
.A2(n_4728),
.B1(n_4739),
.B2(n_4734),
.Y(n_6493)
);

OAI22xp5_ASAP7_75t_L g6494 ( 
.A1(n_4739),
.A2(n_4762),
.B1(n_4765),
.B2(n_4754),
.Y(n_6494)
);

AOI22xp33_ASAP7_75t_L g6495 ( 
.A1(n_5110),
.A2(n_4572),
.B1(n_5410),
.B2(n_5493),
.Y(n_6495)
);

INVxp67_ASAP7_75t_SL g6496 ( 
.A(n_5035),
.Y(n_6496)
);

BUFx2_ASAP7_75t_L g6497 ( 
.A(n_4560),
.Y(n_6497)
);

AOI22xp33_ASAP7_75t_L g6498 ( 
.A1(n_5410),
.A2(n_5493),
.B1(n_5510),
.B2(n_4982),
.Y(n_6498)
);

AOI22xp33_ASAP7_75t_L g6499 ( 
.A1(n_5510),
.A2(n_4982),
.B1(n_5118),
.B2(n_5109),
.Y(n_6499)
);

A2O1A1Ixp33_ASAP7_75t_L g6500 ( 
.A1(n_4640),
.A2(n_5413),
.B(n_5395),
.C(n_4714),
.Y(n_6500)
);

O2A1O1Ixp5_ASAP7_75t_L g6501 ( 
.A1(n_5478),
.A2(n_5434),
.B(n_5417),
.C(n_5215),
.Y(n_6501)
);

INVx1_ASAP7_75t_SL g6502 ( 
.A(n_4870),
.Y(n_6502)
);

AOI21xp33_ASAP7_75t_L g6503 ( 
.A1(n_5406),
.A2(n_5412),
.B(n_4542),
.Y(n_6503)
);

NAND2x1_ASAP7_75t_L g6504 ( 
.A(n_4680),
.B(n_4448),
.Y(n_6504)
);

HB1xp67_ASAP7_75t_L g6505 ( 
.A(n_4761),
.Y(n_6505)
);

AOI22xp5_ASAP7_75t_L g6506 ( 
.A1(n_5046),
.A2(n_4652),
.B1(n_4762),
.B2(n_4754),
.Y(n_6506)
);

A2O1A1Ixp33_ASAP7_75t_L g6507 ( 
.A1(n_5395),
.A2(n_5413),
.B(n_4714),
.C(n_4814),
.Y(n_6507)
);

INVx4_ASAP7_75t_L g6508 ( 
.A(n_4948),
.Y(n_6508)
);

AOI22xp33_ASAP7_75t_L g6509 ( 
.A1(n_5109),
.A2(n_5124),
.B1(n_5226),
.B2(n_5118),
.Y(n_6509)
);

INVxp33_ASAP7_75t_SL g6510 ( 
.A(n_5447),
.Y(n_6510)
);

NOR2xp33_ASAP7_75t_L g6511 ( 
.A(n_4765),
.B(n_4768),
.Y(n_6511)
);

AOI22xp33_ASAP7_75t_L g6512 ( 
.A1(n_5124),
.A2(n_5241),
.B1(n_5263),
.B2(n_5226),
.Y(n_6512)
);

AOI22xp5_ASAP7_75t_L g6513 ( 
.A1(n_4768),
.A2(n_4769),
.B1(n_4782),
.B2(n_4770),
.Y(n_6513)
);

BUFx2_ASAP7_75t_L g6514 ( 
.A(n_4560),
.Y(n_6514)
);

O2A1O1Ixp33_ASAP7_75t_L g6515 ( 
.A1(n_5143),
.A2(n_5418),
.B(n_5434),
.C(n_5448),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_L g6516 ( 
.A(n_4769),
.B(n_4770),
.Y(n_6516)
);

INVx4_ASAP7_75t_L g6517 ( 
.A(n_4948),
.Y(n_6517)
);

A2O1A1Ixp33_ASAP7_75t_L g6518 ( 
.A1(n_5395),
.A2(n_5413),
.B(n_4714),
.C(n_4814),
.Y(n_6518)
);

INVx6_ASAP7_75t_L g6519 ( 
.A(n_5083),
.Y(n_6519)
);

BUFx12f_ASAP7_75t_L g6520 ( 
.A(n_4887),
.Y(n_6520)
);

INVx4_ASAP7_75t_L g6521 ( 
.A(n_4948),
.Y(n_6521)
);

A2O1A1Ixp33_ASAP7_75t_SL g6522 ( 
.A1(n_5409),
.A2(n_5427),
.B(n_5430),
.C(n_5426),
.Y(n_6522)
);

OR2x2_ASAP7_75t_L g6523 ( 
.A(n_5042),
.B(n_5117),
.Y(n_6523)
);

XNOR2xp5_ASAP7_75t_L g6524 ( 
.A(n_4951),
.B(n_4963),
.Y(n_6524)
);

AOI22xp33_ASAP7_75t_L g6525 ( 
.A1(n_5241),
.A2(n_5285),
.B1(n_5332),
.B2(n_5263),
.Y(n_6525)
);

CKINVDCx8_ASAP7_75t_R g6526 ( 
.A(n_4948),
.Y(n_6526)
);

BUFx2_ASAP7_75t_SL g6527 ( 
.A(n_4986),
.Y(n_6527)
);

BUFx3_ASAP7_75t_L g6528 ( 
.A(n_5299),
.Y(n_6528)
);

NAND2x1_ASAP7_75t_SL g6529 ( 
.A(n_5324),
.B(n_5340),
.Y(n_6529)
);

HB1xp67_ASAP7_75t_L g6530 ( 
.A(n_4761),
.Y(n_6530)
);

NOR2xp33_ASAP7_75t_L g6531 ( 
.A(n_4782),
.B(n_4786),
.Y(n_6531)
);

BUFx4f_ASAP7_75t_L g6532 ( 
.A(n_5206),
.Y(n_6532)
);

AOI21x1_ASAP7_75t_L g6533 ( 
.A1(n_4941),
.A2(n_5192),
.B(n_5407),
.Y(n_6533)
);

O2A1O1Ixp33_ASAP7_75t_L g6534 ( 
.A1(n_5418),
.A2(n_5448),
.B(n_5332),
.C(n_5381),
.Y(n_6534)
);

OAI22xp5_ASAP7_75t_L g6535 ( 
.A1(n_4786),
.A2(n_4789),
.B1(n_4791),
.B2(n_4788),
.Y(n_6535)
);

AOI21xp5_ASAP7_75t_L g6536 ( 
.A1(n_4542),
.A2(n_5358),
.B(n_5220),
.Y(n_6536)
);

AND3x1_ASAP7_75t_SL g6537 ( 
.A(n_5146),
.B(n_4567),
.C(n_4420),
.Y(n_6537)
);

CKINVDCx5p33_ASAP7_75t_R g6538 ( 
.A(n_4887),
.Y(n_6538)
);

OAI22xp5_ASAP7_75t_SL g6539 ( 
.A1(n_5316),
.A2(n_4909),
.B1(n_4987),
.B2(n_4958),
.Y(n_6539)
);

CKINVDCx5p33_ASAP7_75t_R g6540 ( 
.A(n_4909),
.Y(n_6540)
);

OAI21x1_ASAP7_75t_L g6541 ( 
.A1(n_5151),
.A2(n_5437),
.B(n_5339),
.Y(n_6541)
);

CKINVDCx5p33_ASAP7_75t_R g6542 ( 
.A(n_4958),
.Y(n_6542)
);

CKINVDCx8_ASAP7_75t_R g6543 ( 
.A(n_4986),
.Y(n_6543)
);

O2A1O1Ixp33_ASAP7_75t_L g6544 ( 
.A1(n_5285),
.A2(n_5391),
.B(n_5394),
.C(n_5381),
.Y(n_6544)
);

AOI22xp5_ASAP7_75t_L g6545 ( 
.A1(n_4788),
.A2(n_4789),
.B1(n_4796),
.B2(n_4791),
.Y(n_6545)
);

NOR2xp67_ASAP7_75t_L g6546 ( 
.A(n_5215),
.B(n_5222),
.Y(n_6546)
);

O2A1O1Ixp33_ASAP7_75t_L g6547 ( 
.A1(n_5391),
.A2(n_5394),
.B(n_4798),
.C(n_4799),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_SL g6548 ( 
.A(n_5364),
.B(n_5446),
.Y(n_6548)
);

INVx3_ASAP7_75t_L g6549 ( 
.A(n_5005),
.Y(n_6549)
);

AOI21xp5_ASAP7_75t_L g6550 ( 
.A1(n_5437),
.A2(n_5359),
.B(n_5092),
.Y(n_6550)
);

BUFx12f_ASAP7_75t_L g6551 ( 
.A(n_4987),
.Y(n_6551)
);

INVx4_ASAP7_75t_L g6552 ( 
.A(n_5166),
.Y(n_6552)
);

INVx8_ASAP7_75t_L g6553 ( 
.A(n_4865),
.Y(n_6553)
);

NAND2xp5_ASAP7_75t_L g6554 ( 
.A(n_4796),
.B(n_4798),
.Y(n_6554)
);

OR2x6_ASAP7_75t_L g6555 ( 
.A(n_5092),
.B(n_5359),
.Y(n_6555)
);

INVx4_ASAP7_75t_L g6556 ( 
.A(n_4986),
.Y(n_6556)
);

CKINVDCx6p67_ASAP7_75t_R g6557 ( 
.A(n_5365),
.Y(n_6557)
);

INVx1_ASAP7_75t_SL g6558 ( 
.A(n_4903),
.Y(n_6558)
);

A2O1A1Ixp33_ASAP7_75t_L g6559 ( 
.A1(n_5395),
.A2(n_5413),
.B(n_4714),
.C(n_4814),
.Y(n_6559)
);

BUFx8_ASAP7_75t_SL g6560 ( 
.A(n_5236),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_SL g6561 ( 
.A(n_5446),
.B(n_5014),
.Y(n_6561)
);

INVx4_ASAP7_75t_L g6562 ( 
.A(n_4986),
.Y(n_6562)
);

A2O1A1Ixp33_ASAP7_75t_L g6563 ( 
.A1(n_5395),
.A2(n_4714),
.B(n_4814),
.C(n_4664),
.Y(n_6563)
);

NOR2xp67_ASAP7_75t_SL g6564 ( 
.A(n_4986),
.B(n_5166),
.Y(n_6564)
);

NAND2xp5_ASAP7_75t_L g6565 ( 
.A(n_4799),
.B(n_4800),
.Y(n_6565)
);

NAND2xp5_ASAP7_75t_L g6566 ( 
.A(n_4800),
.B(n_4804),
.Y(n_6566)
);

AOI21xp5_ASAP7_75t_L g6567 ( 
.A1(n_5437),
.A2(n_5359),
.B(n_5092),
.Y(n_6567)
);

A2O1A1Ixp33_ASAP7_75t_L g6568 ( 
.A1(n_4664),
.A2(n_4966),
.B(n_5132),
.C(n_4814),
.Y(n_6568)
);

INVx1_ASAP7_75t_SL g6569 ( 
.A(n_5509),
.Y(n_6569)
);

NOR2xp33_ASAP7_75t_R g6570 ( 
.A(n_5388),
.B(n_5236),
.Y(n_6570)
);

OR2x2_ASAP7_75t_L g6571 ( 
.A(n_5121),
.B(n_5290),
.Y(n_6571)
);

HB1xp67_ASAP7_75t_L g6572 ( 
.A(n_4792),
.Y(n_6572)
);

A2O1A1Ixp33_ASAP7_75t_L g6573 ( 
.A1(n_4664),
.A2(n_5132),
.B(n_5170),
.C(n_4966),
.Y(n_6573)
);

NAND2xp5_ASAP7_75t_SL g6574 ( 
.A(n_5446),
.B(n_5014),
.Y(n_6574)
);

BUFx6f_ASAP7_75t_SL g6575 ( 
.A(n_4709),
.Y(n_6575)
);

BUFx4f_ASAP7_75t_L g6576 ( 
.A(n_5206),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_4804),
.B(n_4811),
.Y(n_6577)
);

AOI21x1_ASAP7_75t_L g6578 ( 
.A1(n_5192),
.A2(n_5407),
.B(n_5409),
.Y(n_6578)
);

INVx1_ASAP7_75t_SL g6579 ( 
.A(n_5521),
.Y(n_6579)
);

AOI22xp33_ASAP7_75t_SL g6580 ( 
.A1(n_5014),
.A2(n_5068),
.B1(n_5080),
.B2(n_5059),
.Y(n_6580)
);

NAND2x1p5_ASAP7_75t_L g6581 ( 
.A(n_4709),
.B(n_4986),
.Y(n_6581)
);

NOR2xp33_ASAP7_75t_L g6582 ( 
.A(n_4811),
.B(n_4830),
.Y(n_6582)
);

BUFx12f_ASAP7_75t_L g6583 ( 
.A(n_5415),
.Y(n_6583)
);

INVx1_ASAP7_75t_SL g6584 ( 
.A(n_5298),
.Y(n_6584)
);

OR2x6_ASAP7_75t_L g6585 ( 
.A(n_4866),
.B(n_4912),
.Y(n_6585)
);

HB1xp67_ASAP7_75t_L g6586 ( 
.A(n_4792),
.Y(n_6586)
);

O2A1O1Ixp33_ASAP7_75t_L g6587 ( 
.A1(n_4830),
.A2(n_4841),
.B(n_4845),
.C(n_4839),
.Y(n_6587)
);

NOR2xp33_ASAP7_75t_L g6588 ( 
.A(n_4839),
.B(n_4841),
.Y(n_6588)
);

AOI21x1_ASAP7_75t_L g6589 ( 
.A1(n_5427),
.A2(n_5461),
.B(n_5430),
.Y(n_6589)
);

BUFx2_ASAP7_75t_L g6590 ( 
.A(n_5514),
.Y(n_6590)
);

AOI22xp33_ASAP7_75t_L g6591 ( 
.A1(n_4845),
.A2(n_4936),
.B1(n_4950),
.B2(n_4898),
.Y(n_6591)
);

AOI21xp5_ASAP7_75t_L g6592 ( 
.A1(n_5290),
.A2(n_5295),
.B(n_5294),
.Y(n_6592)
);

BUFx2_ASAP7_75t_L g6593 ( 
.A(n_5514),
.Y(n_6593)
);

AOI22xp33_ASAP7_75t_L g6594 ( 
.A1(n_4898),
.A2(n_4906),
.B1(n_4918),
.B2(n_4899),
.Y(n_6594)
);

INVx4_ASAP7_75t_L g6595 ( 
.A(n_4986),
.Y(n_6595)
);

AOI22xp33_ASAP7_75t_SL g6596 ( 
.A1(n_5014),
.A2(n_5068),
.B1(n_5080),
.B2(n_5059),
.Y(n_6596)
);

INVx4_ASAP7_75t_L g6597 ( 
.A(n_4986),
.Y(n_6597)
);

INVxp67_ASAP7_75t_L g6598 ( 
.A(n_5298),
.Y(n_6598)
);

AOI22xp5_ASAP7_75t_L g6599 ( 
.A1(n_4854),
.A2(n_4872),
.B1(n_4878),
.B2(n_4860),
.Y(n_6599)
);

CKINVDCx20_ASAP7_75t_R g6600 ( 
.A(n_5415),
.Y(n_6600)
);

A2O1A1Ixp33_ASAP7_75t_L g6601 ( 
.A1(n_4664),
.A2(n_5132),
.B(n_5170),
.C(n_4966),
.Y(n_6601)
);

O2A1O1Ixp5_ASAP7_75t_SL g6602 ( 
.A1(n_4905),
.A2(n_4908),
.B(n_4907),
.C(n_5399),
.Y(n_6602)
);

INVx1_ASAP7_75t_SL g6603 ( 
.A(n_5298),
.Y(n_6603)
);

BUFx4f_ASAP7_75t_L g6604 ( 
.A(n_5229),
.Y(n_6604)
);

BUFx2_ASAP7_75t_L g6605 ( 
.A(n_5514),
.Y(n_6605)
);

NAND2x2_ASAP7_75t_L g6606 ( 
.A(n_4976),
.B(n_4994),
.Y(n_6606)
);

NOR2xp33_ASAP7_75t_L g6607 ( 
.A(n_4854),
.B(n_4860),
.Y(n_6607)
);

AOI21xp5_ASAP7_75t_L g6608 ( 
.A1(n_5294),
.A2(n_5296),
.B(n_5295),
.Y(n_6608)
);

AOI22xp33_ASAP7_75t_SL g6609 ( 
.A1(n_5014),
.A2(n_5068),
.B1(n_5080),
.B2(n_5059),
.Y(n_6609)
);

AOI22xp33_ASAP7_75t_L g6610 ( 
.A1(n_4914),
.A2(n_4950),
.B1(n_4970),
.B2(n_4936),
.Y(n_6610)
);

INVx1_ASAP7_75t_SL g6611 ( 
.A(n_5315),
.Y(n_6611)
);

INVx2_ASAP7_75t_L g6612 ( 
.A(n_4597),
.Y(n_6612)
);

INVx3_ASAP7_75t_L g6613 ( 
.A(n_5014),
.Y(n_6613)
);

CKINVDCx5p33_ASAP7_75t_R g6614 ( 
.A(n_5486),
.Y(n_6614)
);

INVx1_ASAP7_75t_SL g6615 ( 
.A(n_5315),
.Y(n_6615)
);

BUFx12f_ASAP7_75t_L g6616 ( 
.A(n_5486),
.Y(n_6616)
);

INVx2_ASAP7_75t_SL g6617 ( 
.A(n_5014),
.Y(n_6617)
);

A2O1A1Ixp33_ASAP7_75t_L g6618 ( 
.A1(n_4664),
.A2(n_5132),
.B(n_5170),
.C(n_4966),
.Y(n_6618)
);

NAND2xp5_ASAP7_75t_L g6619 ( 
.A(n_4872),
.B(n_4878),
.Y(n_6619)
);

INVx2_ASAP7_75t_SL g6620 ( 
.A(n_5059),
.Y(n_6620)
);

AOI22xp5_ASAP7_75t_L g6621 ( 
.A1(n_4889),
.A2(n_4899),
.B1(n_4900),
.B2(n_4891),
.Y(n_6621)
);

CKINVDCx5p33_ASAP7_75t_R g6622 ( 
.A(n_5780),
.Y(n_6622)
);

AND2x4_ASAP7_75t_L g6623 ( 
.A(n_5795),
.B(n_4925),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_L g6624 ( 
.A(n_5673),
.B(n_5121),
.Y(n_6624)
);

AND2x4_ASAP7_75t_L g6625 ( 
.A(n_5795),
.B(n_4925),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_5546),
.Y(n_6626)
);

INVx2_ASAP7_75t_SL g6627 ( 
.A(n_5566),
.Y(n_6627)
);

NAND2xp5_ASAP7_75t_L g6628 ( 
.A(n_5673),
.B(n_5788),
.Y(n_6628)
);

NAND2xp5_ASAP7_75t_L g6629 ( 
.A(n_5788),
.B(n_4905),
.Y(n_6629)
);

INVx2_ASAP7_75t_SL g6630 ( 
.A(n_5566),
.Y(n_6630)
);

BUFx6f_ASAP7_75t_L g6631 ( 
.A(n_6097),
.Y(n_6631)
);

BUFx3_ASAP7_75t_L g6632 ( 
.A(n_5704),
.Y(n_6632)
);

INVx2_ASAP7_75t_SL g6633 ( 
.A(n_5566),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_5885),
.B(n_4609),
.Y(n_6634)
);

INVx3_ASAP7_75t_L g6635 ( 
.A(n_6097),
.Y(n_6635)
);

HAxp5_ASAP7_75t_L g6636 ( 
.A(n_5897),
.B(n_4420),
.CON(n_6636),
.SN(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_5546),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_5546),
.Y(n_6638)
);

NAND2xp5_ASAP7_75t_L g6639 ( 
.A(n_5843),
.B(n_4907),
.Y(n_6639)
);

INVx4_ASAP7_75t_L g6640 ( 
.A(n_5704),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_5546),
.Y(n_6641)
);

BUFx2_ASAP7_75t_SL g6642 ( 
.A(n_6353),
.Y(n_6642)
);

INVxp67_ASAP7_75t_L g6643 ( 
.A(n_6127),
.Y(n_6643)
);

HB1xp67_ASAP7_75t_L g6644 ( 
.A(n_5580),
.Y(n_6644)
);

INVx3_ASAP7_75t_L g6645 ( 
.A(n_6097),
.Y(n_6645)
);

AND2x4_ASAP7_75t_L g6646 ( 
.A(n_5795),
.B(n_4925),
.Y(n_6646)
);

OAI22xp5_ASAP7_75t_L g6647 ( 
.A1(n_5841),
.A2(n_4914),
.B1(n_4938),
.B2(n_4900),
.Y(n_6647)
);

INVx3_ASAP7_75t_SL g6648 ( 
.A(n_6557),
.Y(n_6648)
);

INVx5_ASAP7_75t_L g6649 ( 
.A(n_6383),
.Y(n_6649)
);

INVx1_ASAP7_75t_SL g6650 ( 
.A(n_5969),
.Y(n_6650)
);

NOR2xp33_ASAP7_75t_SL g6651 ( 
.A(n_5897),
.B(n_5166),
.Y(n_6651)
);

NAND2xp5_ASAP7_75t_L g6652 ( 
.A(n_5843),
.B(n_4822),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_L g6653 ( 
.A(n_5870),
.B(n_4822),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5551),
.Y(n_6654)
);

OAI22xp33_ASAP7_75t_L g6655 ( 
.A1(n_5841),
.A2(n_5068),
.B1(n_5080),
.B2(n_5059),
.Y(n_6655)
);

NAND2x1p5_ASAP7_75t_L g6656 ( 
.A(n_6564),
.B(n_5166),
.Y(n_6656)
);

BUFx3_ASAP7_75t_L g6657 ( 
.A(n_5704),
.Y(n_6657)
);

AND2x4_ASAP7_75t_L g6658 ( 
.A(n_5885),
.B(n_5059),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_5551),
.Y(n_6659)
);

AOI22xp5_ASAP7_75t_L g6660 ( 
.A1(n_5542),
.A2(n_4963),
.B1(n_4974),
.B2(n_4951),
.Y(n_6660)
);

NAND2xp5_ASAP7_75t_L g6661 ( 
.A(n_5870),
.B(n_4692),
.Y(n_6661)
);

AOI21xp5_ASAP7_75t_L g6662 ( 
.A1(n_5802),
.A2(n_5295),
.B(n_5294),
.Y(n_6662)
);

BUFx6f_ASAP7_75t_L g6663 ( 
.A(n_6097),
.Y(n_6663)
);

CKINVDCx20_ASAP7_75t_R g6664 ( 
.A(n_5665),
.Y(n_6664)
);

NAND3xp33_ASAP7_75t_L g6665 ( 
.A(n_5918),
.B(n_5466),
.C(n_5461),
.Y(n_6665)
);

INVx1_ASAP7_75t_L g6666 ( 
.A(n_5551),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_5551),
.Y(n_6667)
);

AOI21xp5_ASAP7_75t_L g6668 ( 
.A1(n_5802),
.A2(n_5297),
.B(n_5296),
.Y(n_6668)
);

OAI22xp33_ASAP7_75t_L g6669 ( 
.A1(n_5851),
.A2(n_5068),
.B1(n_5080),
.B2(n_5059),
.Y(n_6669)
);

BUFx6f_ASAP7_75t_L g6670 ( 
.A(n_6097),
.Y(n_6670)
);

CKINVDCx5p33_ASAP7_75t_R g6671 ( 
.A(n_5780),
.Y(n_6671)
);

NAND2xp5_ASAP7_75t_L g6672 ( 
.A(n_5957),
.B(n_4692),
.Y(n_6672)
);

HB1xp67_ASAP7_75t_L g6673 ( 
.A(n_5580),
.Y(n_6673)
);

AOI22xp33_ASAP7_75t_L g6674 ( 
.A1(n_5542),
.A2(n_4891),
.B1(n_4906),
.B2(n_4889),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_L g6675 ( 
.A(n_5957),
.B(n_4692),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_5885),
.B(n_4609),
.Y(n_6676)
);

AOI21xp5_ASAP7_75t_L g6677 ( 
.A1(n_5559),
.A2(n_5303),
.B(n_5297),
.Y(n_6677)
);

A2O1A1Ixp33_ASAP7_75t_L g6678 ( 
.A1(n_5918),
.A2(n_5324),
.B(n_5388),
.C(n_5132),
.Y(n_6678)
);

NAND2xp5_ASAP7_75t_L g6679 ( 
.A(n_5961),
.B(n_4815),
.Y(n_6679)
);

AOI21xp5_ASAP7_75t_L g6680 ( 
.A1(n_5559),
.A2(n_5562),
.B(n_5958),
.Y(n_6680)
);

INVx2_ASAP7_75t_L g6681 ( 
.A(n_5560),
.Y(n_6681)
);

BUFx3_ASAP7_75t_L g6682 ( 
.A(n_5704),
.Y(n_6682)
);

NAND2xp5_ASAP7_75t_SL g6683 ( 
.A(n_5616),
.B(n_5941),
.Y(n_6683)
);

AOI21xp5_ASAP7_75t_L g6684 ( 
.A1(n_5562),
.A2(n_5303),
.B(n_5297),
.Y(n_6684)
);

BUFx2_ASAP7_75t_L g6685 ( 
.A(n_6529),
.Y(n_6685)
);

INVx5_ASAP7_75t_L g6686 ( 
.A(n_6383),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_5560),
.Y(n_6687)
);

BUFx6f_ASAP7_75t_L g6688 ( 
.A(n_6097),
.Y(n_6688)
);

AOI22xp33_ASAP7_75t_L g6689 ( 
.A1(n_5906),
.A2(n_4911),
.B1(n_4923),
.B2(n_4918),
.Y(n_6689)
);

AOI22xp33_ASAP7_75t_L g6690 ( 
.A1(n_5906),
.A2(n_5671),
.B1(n_5884),
.B2(n_5902),
.Y(n_6690)
);

OAI21xp5_ASAP7_75t_L g6691 ( 
.A1(n_5616),
.A2(n_5487),
.B(n_5468),
.Y(n_6691)
);

BUFx3_ASAP7_75t_L g6692 ( 
.A(n_5704),
.Y(n_6692)
);

AND2x4_ASAP7_75t_L g6693 ( 
.A(n_5937),
.B(n_5068),
.Y(n_6693)
);

AND2x2_ASAP7_75t_SL g6694 ( 
.A(n_6000),
.B(n_5324),
.Y(n_6694)
);

NAND2x1p5_ASAP7_75t_L g6695 ( 
.A(n_6564),
.B(n_5166),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_5560),
.Y(n_6696)
);

CKINVDCx5p33_ASAP7_75t_R g6697 ( 
.A(n_5987),
.Y(n_6697)
);

BUFx2_ASAP7_75t_L g6698 ( 
.A(n_6529),
.Y(n_6698)
);

INVx1_ASAP7_75t_SL g6699 ( 
.A(n_5969),
.Y(n_6699)
);

INVx2_ASAP7_75t_SL g6700 ( 
.A(n_5566),
.Y(n_6700)
);

AND2x4_ASAP7_75t_L g6701 ( 
.A(n_5937),
.B(n_5068),
.Y(n_6701)
);

INVx2_ASAP7_75t_L g6702 ( 
.A(n_5560),
.Y(n_6702)
);

INVx3_ASAP7_75t_L g6703 ( 
.A(n_6097),
.Y(n_6703)
);

BUFx3_ASAP7_75t_L g6704 ( 
.A(n_5704),
.Y(n_6704)
);

AOI21xp5_ASAP7_75t_L g6705 ( 
.A1(n_5958),
.A2(n_5305),
.B(n_5303),
.Y(n_6705)
);

BUFx6f_ASAP7_75t_SL g6706 ( 
.A(n_6157),
.Y(n_6706)
);

AOI21xp5_ASAP7_75t_L g6707 ( 
.A1(n_5565),
.A2(n_5311),
.B(n_5305),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_5561),
.Y(n_6708)
);

AOI21xp5_ASAP7_75t_L g6709 ( 
.A1(n_5565),
.A2(n_5311),
.B(n_5305),
.Y(n_6709)
);

NOR2xp33_ASAP7_75t_L g6710 ( 
.A(n_5979),
.B(n_5146),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_5561),
.Y(n_6711)
);

INVxp67_ASAP7_75t_L g6712 ( 
.A(n_6127),
.Y(n_6712)
);

BUFx2_ASAP7_75t_L g6713 ( 
.A(n_6379),
.Y(n_6713)
);

AOI22xp5_ASAP7_75t_L g6714 ( 
.A1(n_5851),
.A2(n_4963),
.B1(n_4974),
.B2(n_4951),
.Y(n_6714)
);

AND2x4_ASAP7_75t_L g6715 ( 
.A(n_5937),
.B(n_5896),
.Y(n_6715)
);

NAND3xp33_ASAP7_75t_L g6716 ( 
.A(n_5695),
.B(n_5468),
.C(n_5466),
.Y(n_6716)
);

AND2x4_ASAP7_75t_L g6717 ( 
.A(n_5896),
.B(n_5068),
.Y(n_6717)
);

BUFx6f_ASAP7_75t_L g6718 ( 
.A(n_6101),
.Y(n_6718)
);

A2O1A1Ixp33_ASAP7_75t_L g6719 ( 
.A1(n_5695),
.A2(n_5324),
.B(n_5170),
.C(n_4966),
.Y(n_6719)
);

AOI21xp5_ASAP7_75t_L g6720 ( 
.A1(n_5570),
.A2(n_5321),
.B(n_5311),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_5571),
.Y(n_6721)
);

AOI221xp5_ASAP7_75t_L g6722 ( 
.A1(n_5612),
.A2(n_4926),
.B1(n_4931),
.B2(n_4923),
.C(n_4911),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_5531),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_5531),
.Y(n_6724)
);

O2A1O1Ixp5_ASAP7_75t_SL g6725 ( 
.A1(n_5926),
.A2(n_5468),
.B(n_5487),
.C(n_5482),
.Y(n_6725)
);

CKINVDCx5p33_ASAP7_75t_R g6726 ( 
.A(n_5987),
.Y(n_6726)
);

AND2x4_ASAP7_75t_L g6727 ( 
.A(n_5896),
.B(n_5059),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_SL g6728 ( 
.A(n_5941),
.B(n_5059),
.Y(n_6728)
);

NOR2xp33_ASAP7_75t_L g6729 ( 
.A(n_5979),
.B(n_5440),
.Y(n_6729)
);

BUFx2_ASAP7_75t_L g6730 ( 
.A(n_6379),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_5533),
.Y(n_6731)
);

AND2x4_ASAP7_75t_L g6732 ( 
.A(n_5896),
.B(n_5068),
.Y(n_6732)
);

BUFx6f_ASAP7_75t_L g6733 ( 
.A(n_6101),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_5571),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_5533),
.Y(n_6735)
);

HB1xp67_ASAP7_75t_L g6736 ( 
.A(n_5590),
.Y(n_6736)
);

AND2x4_ASAP7_75t_L g6737 ( 
.A(n_5896),
.B(n_5080),
.Y(n_6737)
);

AOI21x1_ASAP7_75t_L g6738 ( 
.A1(n_6237),
.A2(n_5187),
.B(n_5185),
.Y(n_6738)
);

NAND2xp33_ASAP7_75t_L g6739 ( 
.A(n_5650),
.B(n_4463),
.Y(n_6739)
);

BUFx4_ASAP7_75t_SL g6740 ( 
.A(n_6235),
.Y(n_6740)
);

NAND2xp5_ASAP7_75t_L g6741 ( 
.A(n_5956),
.B(n_5315),
.Y(n_6741)
);

INVx2_ASAP7_75t_L g6742 ( 
.A(n_5571),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6411),
.B(n_4609),
.Y(n_6743)
);

INVx4_ASAP7_75t_L g6744 ( 
.A(n_5997),
.Y(n_6744)
);

NOR2x1_ASAP7_75t_SL g6745 ( 
.A(n_6527),
.B(n_5324),
.Y(n_6745)
);

INVx2_ASAP7_75t_L g6746 ( 
.A(n_5571),
.Y(n_6746)
);

BUFx2_ASAP7_75t_L g6747 ( 
.A(n_6379),
.Y(n_6747)
);

NAND2xp5_ASAP7_75t_L g6748 ( 
.A(n_5956),
.B(n_5361),
.Y(n_6748)
);

INVxp67_ASAP7_75t_L g6749 ( 
.A(n_5590),
.Y(n_6749)
);

BUFx12f_ASAP7_75t_L g6750 ( 
.A(n_5593),
.Y(n_6750)
);

AND2x6_ASAP7_75t_L g6751 ( 
.A(n_5579),
.B(n_5229),
.Y(n_6751)
);

INVx2_ASAP7_75t_L g6752 ( 
.A(n_5596),
.Y(n_6752)
);

AOI22xp5_ASAP7_75t_L g6753 ( 
.A1(n_5884),
.A2(n_4963),
.B1(n_4974),
.B2(n_4951),
.Y(n_6753)
);

AOI21xp5_ASAP7_75t_L g6754 ( 
.A1(n_5570),
.A2(n_5943),
.B(n_6337),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_5596),
.Y(n_6755)
);

AOI21xp5_ASAP7_75t_L g6756 ( 
.A1(n_5943),
.A2(n_5326),
.B(n_5321),
.Y(n_6756)
);

INVx3_ASAP7_75t_SL g6757 ( 
.A(n_6557),
.Y(n_6757)
);

AOI21xp5_ASAP7_75t_L g6758 ( 
.A1(n_6337),
.A2(n_5326),
.B(n_5321),
.Y(n_6758)
);

NAND2x1p5_ASAP7_75t_L g6759 ( 
.A(n_6564),
.B(n_5166),
.Y(n_6759)
);

BUFx10_ASAP7_75t_L g6760 ( 
.A(n_5679),
.Y(n_6760)
);

INVxp67_ASAP7_75t_L g6761 ( 
.A(n_5597),
.Y(n_6761)
);

INVx2_ASAP7_75t_SL g6762 ( 
.A(n_5566),
.Y(n_6762)
);

O2A1O1Ixp33_ASAP7_75t_L g6763 ( 
.A1(n_5650),
.A2(n_5612),
.B(n_6305),
.C(n_5925),
.Y(n_6763)
);

CKINVDCx20_ASAP7_75t_R g6764 ( 
.A(n_5665),
.Y(n_6764)
);

INVxp67_ASAP7_75t_L g6765 ( 
.A(n_5597),
.Y(n_6765)
);

INVx3_ASAP7_75t_L g6766 ( 
.A(n_6101),
.Y(n_6766)
);

NOR2xp33_ASAP7_75t_L g6767 ( 
.A(n_5666),
.B(n_5440),
.Y(n_6767)
);

AND2x2_ASAP7_75t_L g6768 ( 
.A(n_6411),
.B(n_4609),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_5540),
.Y(n_6769)
);

AOI21xp5_ASAP7_75t_L g6770 ( 
.A1(n_6465),
.A2(n_5883),
.B(n_5875),
.Y(n_6770)
);

AOI21xp5_ASAP7_75t_L g6771 ( 
.A1(n_6465),
.A2(n_5883),
.B(n_5875),
.Y(n_6771)
);

BUFx6f_ASAP7_75t_L g6772 ( 
.A(n_6101),
.Y(n_6772)
);

NOR2xp67_ASAP7_75t_L g6773 ( 
.A(n_5754),
.B(n_5222),
.Y(n_6773)
);

NAND2x1p5_ASAP7_75t_L g6774 ( 
.A(n_5754),
.B(n_5166),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_5540),
.Y(n_6775)
);

AND2x4_ASAP7_75t_L g6776 ( 
.A(n_5896),
.B(n_5080),
.Y(n_6776)
);

NAND2xp5_ASAP7_75t_L g6777 ( 
.A(n_5961),
.B(n_4815),
.Y(n_6777)
);

OAI22xp33_ASAP7_75t_SL g6778 ( 
.A1(n_5905),
.A2(n_5502),
.B1(n_5504),
.B2(n_5500),
.Y(n_6778)
);

AOI22xp5_ASAP7_75t_L g6779 ( 
.A1(n_5671),
.A2(n_4963),
.B1(n_4974),
.B2(n_4951),
.Y(n_6779)
);

NAND2xp5_ASAP7_75t_SL g6780 ( 
.A(n_5953),
.B(n_5080),
.Y(n_6780)
);

INVx3_ASAP7_75t_SL g6781 ( 
.A(n_6557),
.Y(n_6781)
);

NAND2xp33_ASAP7_75t_L g6782 ( 
.A(n_5889),
.B(n_4865),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_5596),
.Y(n_6783)
);

INVx2_ASAP7_75t_SL g6784 ( 
.A(n_5566),
.Y(n_6784)
);

BUFx6f_ASAP7_75t_L g6785 ( 
.A(n_6116),
.Y(n_6785)
);

NAND2xp5_ASAP7_75t_L g6786 ( 
.A(n_6378),
.B(n_6323),
.Y(n_6786)
);

NAND2xp5_ASAP7_75t_L g6787 ( 
.A(n_6378),
.B(n_6323),
.Y(n_6787)
);

CKINVDCx20_ASAP7_75t_R g6788 ( 
.A(n_5815),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_5544),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_L g6790 ( 
.A(n_6378),
.B(n_4815),
.Y(n_6790)
);

INVx2_ASAP7_75t_SL g6791 ( 
.A(n_5566),
.Y(n_6791)
);

BUFx2_ASAP7_75t_L g6792 ( 
.A(n_6379),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_L g6793 ( 
.A(n_6200),
.B(n_4794),
.Y(n_6793)
);

BUFx4_ASAP7_75t_SL g6794 ( 
.A(n_6235),
.Y(n_6794)
);

BUFx12f_ASAP7_75t_L g6795 ( 
.A(n_5593),
.Y(n_6795)
);

INVx5_ASAP7_75t_L g6796 ( 
.A(n_6383),
.Y(n_6796)
);

BUFx2_ASAP7_75t_L g6797 ( 
.A(n_6379),
.Y(n_6797)
);

HB1xp67_ASAP7_75t_L g6798 ( 
.A(n_6395),
.Y(n_6798)
);

AND2x2_ASAP7_75t_L g6799 ( 
.A(n_6411),
.B(n_4609),
.Y(n_6799)
);

INVxp67_ASAP7_75t_L g6800 ( 
.A(n_6003),
.Y(n_6800)
);

NAND2xp5_ASAP7_75t_L g6801 ( 
.A(n_6200),
.B(n_6366),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_5544),
.Y(n_6802)
);

HB1xp67_ASAP7_75t_L g6803 ( 
.A(n_6395),
.Y(n_6803)
);

AOI21xp5_ASAP7_75t_L g6804 ( 
.A1(n_6550),
.A2(n_5327),
.B(n_5326),
.Y(n_6804)
);

O2A1O1Ixp5_ASAP7_75t_SL g6805 ( 
.A1(n_5926),
.A2(n_5482),
.B(n_5495),
.C(n_5487),
.Y(n_6805)
);

BUFx6f_ASAP7_75t_L g6806 ( 
.A(n_6116),
.Y(n_6806)
);

INVx8_ASAP7_75t_L g6807 ( 
.A(n_6553),
.Y(n_6807)
);

AOI22xp5_ASAP7_75t_L g6808 ( 
.A1(n_5902),
.A2(n_4963),
.B1(n_4974),
.B2(n_4951),
.Y(n_6808)
);

AOI22xp5_ASAP7_75t_L g6809 ( 
.A1(n_5904),
.A2(n_5007),
.B1(n_5018),
.B2(n_4974),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_5552),
.Y(n_6810)
);

BUFx12f_ASAP7_75t_L g6811 ( 
.A(n_5593),
.Y(n_6811)
);

BUFx2_ASAP7_75t_L g6812 ( 
.A(n_6379),
.Y(n_6812)
);

AOI22xp33_ASAP7_75t_L g6813 ( 
.A1(n_5938),
.A2(n_4931),
.B1(n_4934),
.B2(n_4926),
.Y(n_6813)
);

CKINVDCx5p33_ASAP7_75t_R g6814 ( 
.A(n_6560),
.Y(n_6814)
);

CKINVDCx11_ASAP7_75t_R g6815 ( 
.A(n_5815),
.Y(n_6815)
);

INVx1_ASAP7_75t_SL g6816 ( 
.A(n_6414),
.Y(n_6816)
);

AND2x6_ASAP7_75t_L g6817 ( 
.A(n_5579),
.B(n_5229),
.Y(n_6817)
);

OR2x2_ASAP7_75t_L g6818 ( 
.A(n_6308),
.B(n_6148),
.Y(n_6818)
);

OAI22xp5_ASAP7_75t_L g6819 ( 
.A1(n_5889),
.A2(n_4977),
.B1(n_5027),
.B2(n_4934),
.Y(n_6819)
);

BUFx2_ASAP7_75t_L g6820 ( 
.A(n_6379),
.Y(n_6820)
);

AOI21xp5_ASAP7_75t_L g6821 ( 
.A1(n_6550),
.A2(n_6567),
.B(n_5905),
.Y(n_6821)
);

INVx1_ASAP7_75t_SL g6822 ( 
.A(n_6414),
.Y(n_6822)
);

CKINVDCx8_ASAP7_75t_R g6823 ( 
.A(n_5583),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_5552),
.Y(n_6824)
);

NOR2xp33_ASAP7_75t_L g6825 ( 
.A(n_5666),
.B(n_5440),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_5577),
.Y(n_6826)
);

AND2x4_ASAP7_75t_L g6827 ( 
.A(n_5734),
.B(n_5096),
.Y(n_6827)
);

NAND2xp5_ASAP7_75t_L g6828 ( 
.A(n_6366),
.B(n_5907),
.Y(n_6828)
);

AND2x4_ASAP7_75t_L g6829 ( 
.A(n_5734),
.B(n_5096),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_5907),
.B(n_4794),
.Y(n_6830)
);

NAND2xp5_ASAP7_75t_L g6831 ( 
.A(n_6293),
.B(n_4803),
.Y(n_6831)
);

INVx2_ASAP7_75t_L g6832 ( 
.A(n_5596),
.Y(n_6832)
);

BUFx6f_ASAP7_75t_L g6833 ( 
.A(n_6116),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6290),
.B(n_4612),
.Y(n_6834)
);

CKINVDCx6p67_ASAP7_75t_R g6835 ( 
.A(n_5644),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_5604),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_5577),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6293),
.B(n_4803),
.Y(n_6838)
);

CKINVDCx20_ASAP7_75t_R g6839 ( 
.A(n_6041),
.Y(n_6839)
);

NOR2x1_ASAP7_75t_L g6840 ( 
.A(n_6003),
.B(n_5340),
.Y(n_6840)
);

AOI22xp33_ASAP7_75t_L g6841 ( 
.A1(n_5938),
.A2(n_4942),
.B1(n_4968),
.B2(n_4938),
.Y(n_6841)
);

AOI22xp33_ASAP7_75t_L g6842 ( 
.A1(n_6209),
.A2(n_4968),
.B1(n_4970),
.B2(n_4942),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_5604),
.Y(n_6843)
);

BUFx6f_ASAP7_75t_L g6844 ( 
.A(n_6116),
.Y(n_6844)
);

AOI21xp5_ASAP7_75t_L g6845 ( 
.A1(n_6567),
.A2(n_5337),
.B(n_5327),
.Y(n_6845)
);

INVx3_ASAP7_75t_L g6846 ( 
.A(n_6116),
.Y(n_6846)
);

BUFx2_ASAP7_75t_L g6847 ( 
.A(n_6379),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_5578),
.Y(n_6848)
);

INVx3_ASAP7_75t_L g6849 ( 
.A(n_6116),
.Y(n_6849)
);

AOI21xp5_ASAP7_75t_L g6850 ( 
.A1(n_5942),
.A2(n_5337),
.B(n_5327),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_5578),
.Y(n_6851)
);

BUFx2_ASAP7_75t_L g6852 ( 
.A(n_6395),
.Y(n_6852)
);

AND2x4_ASAP7_75t_L g6853 ( 
.A(n_5734),
.B(n_5096),
.Y(n_6853)
);

INVx8_ASAP7_75t_L g6854 ( 
.A(n_6553),
.Y(n_6854)
);

BUFx4_ASAP7_75t_SL g6855 ( 
.A(n_5603),
.Y(n_6855)
);

INVx3_ASAP7_75t_L g6856 ( 
.A(n_6116),
.Y(n_6856)
);

AOI22xp33_ASAP7_75t_L g6857 ( 
.A1(n_6209),
.A2(n_4977),
.B1(n_4978),
.B2(n_4972),
.Y(n_6857)
);

OAI22xp5_ASAP7_75t_L g6858 ( 
.A1(n_5915),
.A2(n_5027),
.B1(n_4978),
.B2(n_4984),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_SL g6859 ( 
.A(n_5953),
.B(n_5096),
.Y(n_6859)
);

INVx2_ASAP7_75t_L g6860 ( 
.A(n_5604),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_SL g6861 ( 
.A(n_5976),
.B(n_5096),
.Y(n_6861)
);

O2A1O1Ixp33_ASAP7_75t_L g6862 ( 
.A1(n_6305),
.A2(n_4984),
.B(n_4985),
.C(n_4972),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_6317),
.B(n_4827),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_5604),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_5584),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_5584),
.Y(n_6866)
);

CKINVDCx5p33_ASAP7_75t_R g6867 ( 
.A(n_6560),
.Y(n_6867)
);

INVx3_ASAP7_75t_L g6868 ( 
.A(n_6116),
.Y(n_6868)
);

AOI21x1_ASAP7_75t_L g6869 ( 
.A1(n_6237),
.A2(n_5187),
.B(n_5185),
.Y(n_6869)
);

AO21x1_ASAP7_75t_L g6870 ( 
.A1(n_6220),
.A2(n_5399),
.B(n_4700),
.Y(n_6870)
);

INVx2_ASAP7_75t_L g6871 ( 
.A(n_5625),
.Y(n_6871)
);

INVx3_ASAP7_75t_L g6872 ( 
.A(n_6119),
.Y(n_6872)
);

OAI22xp5_ASAP7_75t_L g6873 ( 
.A1(n_5915),
.A2(n_5044),
.B1(n_5058),
.B2(n_4985),
.Y(n_6873)
);

OAI22xp5_ASAP7_75t_L g6874 ( 
.A1(n_5910),
.A2(n_5021),
.B1(n_4988),
.B2(n_4997),
.Y(n_6874)
);

AOI22xp5_ASAP7_75t_L g6875 ( 
.A1(n_5904),
.A2(n_5018),
.B1(n_5072),
.B2(n_5007),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6290),
.B(n_4612),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6290),
.B(n_4612),
.Y(n_6877)
);

CKINVDCx5p33_ASAP7_75t_R g6878 ( 
.A(n_5971),
.Y(n_6878)
);

AOI21xp5_ASAP7_75t_L g6879 ( 
.A1(n_5942),
.A2(n_5341),
.B(n_5337),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_5600),
.Y(n_6880)
);

AOI21xp5_ASAP7_75t_L g6881 ( 
.A1(n_5587),
.A2(n_5608),
.B(n_6433),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_5600),
.Y(n_6882)
);

AOI22xp33_ASAP7_75t_L g6883 ( 
.A1(n_5910),
.A2(n_4995),
.B1(n_4997),
.B2(n_4988),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_6317),
.B(n_4827),
.Y(n_6884)
);

INVx1_ASAP7_75t_SL g6885 ( 
.A(n_6523),
.Y(n_6885)
);

O2A1O1Ixp33_ASAP7_75t_SL g6886 ( 
.A1(n_5966),
.A2(n_5006),
.B(n_5010),
.C(n_4995),
.Y(n_6886)
);

INVx1_ASAP7_75t_SL g6887 ( 
.A(n_6523),
.Y(n_6887)
);

AND2x2_ASAP7_75t_L g6888 ( 
.A(n_6296),
.B(n_4612),
.Y(n_6888)
);

INVx1_ASAP7_75t_L g6889 ( 
.A(n_5614),
.Y(n_6889)
);

HB1xp67_ASAP7_75t_L g6890 ( 
.A(n_6407),
.Y(n_6890)
);

AOI21xp5_ASAP7_75t_L g6891 ( 
.A1(n_5587),
.A2(n_5347),
.B(n_5341),
.Y(n_6891)
);

INVx2_ASAP7_75t_SL g6892 ( 
.A(n_5566),
.Y(n_6892)
);

INVx2_ASAP7_75t_L g6893 ( 
.A(n_5625),
.Y(n_6893)
);

NAND2xp5_ASAP7_75t_L g6894 ( 
.A(n_6009),
.B(n_5361),
.Y(n_6894)
);

INVx5_ASAP7_75t_L g6895 ( 
.A(n_6383),
.Y(n_6895)
);

AOI22xp33_ASAP7_75t_L g6896 ( 
.A1(n_5931),
.A2(n_5006),
.B1(n_5013),
.B2(n_5010),
.Y(n_6896)
);

AOI22xp5_ASAP7_75t_L g6897 ( 
.A1(n_5931),
.A2(n_5018),
.B1(n_5072),
.B2(n_5007),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_5625),
.Y(n_6898)
);

AOI22xp33_ASAP7_75t_L g6899 ( 
.A1(n_5927),
.A2(n_5021),
.B1(n_5025),
.B2(n_5013),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_5625),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6296),
.B(n_4612),
.Y(n_6901)
);

INVx1_ASAP7_75t_SL g6902 ( 
.A(n_6523),
.Y(n_6902)
);

INVx2_ASAP7_75t_L g6903 ( 
.A(n_5633),
.Y(n_6903)
);

AOI22xp33_ASAP7_75t_L g6904 ( 
.A1(n_5927),
.A2(n_5028),
.B1(n_5029),
.B2(n_5025),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_5614),
.Y(n_6905)
);

BUFx2_ASAP7_75t_L g6906 ( 
.A(n_6407),
.Y(n_6906)
);

BUFx10_ASAP7_75t_L g6907 ( 
.A(n_5679),
.Y(n_6907)
);

INVx5_ASAP7_75t_L g6908 ( 
.A(n_6383),
.Y(n_6908)
);

HB1xp67_ASAP7_75t_L g6909 ( 
.A(n_6407),
.Y(n_6909)
);

AOI21x1_ASAP7_75t_SL g6910 ( 
.A1(n_6009),
.A2(n_4593),
.B(n_5360),
.Y(n_6910)
);

AND2x4_ASAP7_75t_L g6911 ( 
.A(n_5576),
.B(n_5096),
.Y(n_6911)
);

INVx4_ASAP7_75t_L g6912 ( 
.A(n_6519),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_5619),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6245),
.B(n_5361),
.Y(n_6914)
);

NAND2xp5_ASAP7_75t_L g6915 ( 
.A(n_6245),
.B(n_5374),
.Y(n_6915)
);

AND2x4_ASAP7_75t_L g6916 ( 
.A(n_5576),
.B(n_5096),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_5619),
.Y(n_6917)
);

AND2x2_ASAP7_75t_L g6918 ( 
.A(n_6296),
.B(n_4612),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_5635),
.Y(n_6919)
);

NOR2xp33_ASAP7_75t_L g6920 ( 
.A(n_6063),
.B(n_5028),
.Y(n_6920)
);

AOI22xp33_ASAP7_75t_L g6921 ( 
.A1(n_5558),
.A2(n_5031),
.B1(n_5036),
.B2(n_5029),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_5635),
.Y(n_6922)
);

INVx2_ASAP7_75t_SL g6923 ( 
.A(n_5576),
.Y(n_6923)
);

INVx3_ASAP7_75t_L g6924 ( 
.A(n_6119),
.Y(n_6924)
);

CKINVDCx5p33_ASAP7_75t_R g6925 ( 
.A(n_5971),
.Y(n_6925)
);

INVx2_ASAP7_75t_L g6926 ( 
.A(n_5633),
.Y(n_6926)
);

NAND2xp5_ASAP7_75t_L g6927 ( 
.A(n_5700),
.B(n_5374),
.Y(n_6927)
);

INVx2_ASAP7_75t_SL g6928 ( 
.A(n_5576),
.Y(n_6928)
);

INVx2_ASAP7_75t_SL g6929 ( 
.A(n_5576),
.Y(n_6929)
);

INVx2_ASAP7_75t_L g6930 ( 
.A(n_5633),
.Y(n_6930)
);

NAND2xp5_ASAP7_75t_L g6931 ( 
.A(n_5700),
.B(n_6146),
.Y(n_6931)
);

OAI22xp5_ASAP7_75t_L g6932 ( 
.A1(n_5982),
.A2(n_5036),
.B1(n_5044),
.B2(n_5031),
.Y(n_6932)
);

NAND3xp33_ASAP7_75t_L g6933 ( 
.A(n_5925),
.B(n_5495),
.C(n_5482),
.Y(n_6933)
);

NAND2xp5_ASAP7_75t_L g6934 ( 
.A(n_6146),
.B(n_5374),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_5633),
.Y(n_6935)
);

BUFx6f_ASAP7_75t_L g6936 ( 
.A(n_6119),
.Y(n_6936)
);

NAND2x1p5_ASAP7_75t_L g6937 ( 
.A(n_5754),
.B(n_5166),
.Y(n_6937)
);

CKINVDCx20_ASAP7_75t_R g6938 ( 
.A(n_6041),
.Y(n_6938)
);

INVx4_ASAP7_75t_L g6939 ( 
.A(n_6519),
.Y(n_6939)
);

INVx2_ASAP7_75t_L g6940 ( 
.A(n_5638),
.Y(n_6940)
);

BUFx6f_ASAP7_75t_L g6941 ( 
.A(n_6119),
.Y(n_6941)
);

AND2x4_ASAP7_75t_L g6942 ( 
.A(n_5576),
.B(n_5594),
.Y(n_6942)
);

OAI21x1_ASAP7_75t_L g6943 ( 
.A1(n_6536),
.A2(n_4432),
.B(n_5185),
.Y(n_6943)
);

BUFx3_ASAP7_75t_L g6944 ( 
.A(n_5844),
.Y(n_6944)
);

INVx2_ASAP7_75t_L g6945 ( 
.A(n_5638),
.Y(n_6945)
);

BUFx3_ASAP7_75t_L g6946 ( 
.A(n_5844),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_5638),
.Y(n_6947)
);

BUFx6f_ASAP7_75t_L g6948 ( 
.A(n_6119),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_5643),
.Y(n_6949)
);

INVx4_ASAP7_75t_L g6950 ( 
.A(n_6519),
.Y(n_6950)
);

BUFx6f_ASAP7_75t_L g6951 ( 
.A(n_6119),
.Y(n_6951)
);

NAND2x1p5_ASAP7_75t_L g6952 ( 
.A(n_5754),
.B(n_5166),
.Y(n_6952)
);

BUFx3_ASAP7_75t_L g6953 ( 
.A(n_5844),
.Y(n_6953)
);

AOI22xp33_ASAP7_75t_L g6954 ( 
.A1(n_5558),
.A2(n_5057),
.B1(n_5058),
.B2(n_5055),
.Y(n_6954)
);

NAND2xp5_ASAP7_75t_L g6955 ( 
.A(n_5888),
.B(n_5396),
.Y(n_6955)
);

NAND2x1p5_ASAP7_75t_L g6956 ( 
.A(n_5754),
.B(n_5153),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_5643),
.Y(n_6957)
);

NAND2xp5_ASAP7_75t_SL g6958 ( 
.A(n_5976),
.B(n_5104),
.Y(n_6958)
);

NAND2xp5_ASAP7_75t_L g6959 ( 
.A(n_5888),
.B(n_5396),
.Y(n_6959)
);

AOI22xp33_ASAP7_75t_L g6960 ( 
.A1(n_6036),
.A2(n_5057),
.B1(n_5055),
.B2(n_5007),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_5638),
.Y(n_6961)
);

BUFx3_ASAP7_75t_L g6962 ( 
.A(n_5887),
.Y(n_6962)
);

INVx2_ASAP7_75t_L g6963 ( 
.A(n_5641),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6321),
.B(n_4612),
.Y(n_6964)
);

INVx6_ASAP7_75t_L g6965 ( 
.A(n_5557),
.Y(n_6965)
);

BUFx3_ASAP7_75t_L g6966 ( 
.A(n_5887),
.Y(n_6966)
);

INVx4_ASAP7_75t_L g6967 ( 
.A(n_6519),
.Y(n_6967)
);

AOI22xp33_ASAP7_75t_L g6968 ( 
.A1(n_6036),
.A2(n_6028),
.B1(n_5543),
.B2(n_5981),
.Y(n_6968)
);

AND2x4_ASAP7_75t_L g6969 ( 
.A(n_5576),
.B(n_5113),
.Y(n_6969)
);

NAND2xp5_ASAP7_75t_L g6970 ( 
.A(n_5994),
.B(n_5396),
.Y(n_6970)
);

BUFx3_ASAP7_75t_L g6971 ( 
.A(n_5887),
.Y(n_6971)
);

INVx5_ASAP7_75t_L g6972 ( 
.A(n_6383),
.Y(n_6972)
);

CKINVDCx20_ASAP7_75t_R g6973 ( 
.A(n_6272),
.Y(n_6973)
);

HB1xp67_ASAP7_75t_L g6974 ( 
.A(n_6464),
.Y(n_6974)
);

INVx2_ASAP7_75t_SL g6975 ( 
.A(n_5576),
.Y(n_6975)
);

NAND2xp5_ASAP7_75t_L g6976 ( 
.A(n_5994),
.B(n_5405),
.Y(n_6976)
);

A2O1A1Ixp33_ASAP7_75t_L g6977 ( 
.A1(n_5966),
.A2(n_5170),
.B(n_5446),
.C(n_5023),
.Y(n_6977)
);

INVx2_ASAP7_75t_SL g6978 ( 
.A(n_5594),
.Y(n_6978)
);

NOR2xp67_ASAP7_75t_SL g6979 ( 
.A(n_5944),
.B(n_5498),
.Y(n_6979)
);

AND2x2_ASAP7_75t_SL g6980 ( 
.A(n_6000),
.B(n_5446),
.Y(n_6980)
);

INVx1_ASAP7_75t_SL g6981 ( 
.A(n_6571),
.Y(n_6981)
);

BUFx4f_ASAP7_75t_L g6982 ( 
.A(n_5656),
.Y(n_6982)
);

NAND2xp5_ASAP7_75t_SL g6983 ( 
.A(n_5981),
.B(n_5982),
.Y(n_6983)
);

INVx3_ASAP7_75t_L g6984 ( 
.A(n_6119),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_5657),
.Y(n_6985)
);

INVx3_ASAP7_75t_L g6986 ( 
.A(n_6119),
.Y(n_6986)
);

INVx3_ASAP7_75t_R g6987 ( 
.A(n_6044),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_5657),
.Y(n_6988)
);

BUFx6f_ASAP7_75t_L g6989 ( 
.A(n_6134),
.Y(n_6989)
);

NAND2xp5_ASAP7_75t_L g6990 ( 
.A(n_6002),
.B(n_5405),
.Y(n_6990)
);

CKINVDCx5p33_ASAP7_75t_R g6991 ( 
.A(n_6445),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_5660),
.Y(n_6992)
);

BUFx12f_ASAP7_75t_L g6993 ( 
.A(n_5632),
.Y(n_6993)
);

AOI21xp5_ASAP7_75t_L g6994 ( 
.A1(n_6433),
.A2(n_5357),
.B(n_5354),
.Y(n_6994)
);

CKINVDCx20_ASAP7_75t_R g6995 ( 
.A(n_6272),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_5660),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_5664),
.Y(n_6997)
);

AND2x2_ASAP7_75t_L g6998 ( 
.A(n_5721),
.B(n_4623),
.Y(n_6998)
);

CKINVDCx11_ASAP7_75t_R g6999 ( 
.A(n_5632),
.Y(n_6999)
);

BUFx2_ASAP7_75t_L g7000 ( 
.A(n_6464),
.Y(n_7000)
);

BUFx3_ASAP7_75t_L g7001 ( 
.A(n_6504),
.Y(n_7001)
);

A2O1A1Ixp33_ASAP7_75t_L g7002 ( 
.A1(n_6444),
.A2(n_5023),
.B(n_5026),
.C(n_4994),
.Y(n_7002)
);

NOR2x1_ASAP7_75t_L g7003 ( 
.A(n_6064),
.B(n_5179),
.Y(n_7003)
);

BUFx2_ASAP7_75t_L g7004 ( 
.A(n_6464),
.Y(n_7004)
);

NOR2xp33_ASAP7_75t_L g7005 ( 
.A(n_6063),
.B(n_4422),
.Y(n_7005)
);

AOI22xp33_ASAP7_75t_L g7006 ( 
.A1(n_6028),
.A2(n_5007),
.B1(n_5072),
.B2(n_5018),
.Y(n_7006)
);

INVx4_ASAP7_75t_L g7007 ( 
.A(n_6519),
.Y(n_7007)
);

CKINVDCx20_ASAP7_75t_R g7008 ( 
.A(n_6600),
.Y(n_7008)
);

BUFx6f_ASAP7_75t_L g7009 ( 
.A(n_6134),
.Y(n_7009)
);

NOR2xp33_ASAP7_75t_L g7010 ( 
.A(n_6019),
.B(n_4422),
.Y(n_7010)
);

AND2x2_ASAP7_75t_L g7011 ( 
.A(n_5721),
.B(n_4623),
.Y(n_7011)
);

HB1xp67_ASAP7_75t_L g7012 ( 
.A(n_6475),
.Y(n_7012)
);

AOI21xp5_ASAP7_75t_L g7013 ( 
.A1(n_6440),
.A2(n_5362),
.B(n_5357),
.Y(n_7013)
);

INVx1_ASAP7_75t_SL g7014 ( 
.A(n_6571),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_5901),
.B(n_4868),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_5664),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_5721),
.B(n_4623),
.Y(n_7017)
);

O2A1O1Ixp33_ASAP7_75t_L g7018 ( 
.A1(n_6376),
.A2(n_5525),
.B(n_5502),
.C(n_5504),
.Y(n_7018)
);

BUFx6f_ASAP7_75t_L g7019 ( 
.A(n_6134),
.Y(n_7019)
);

BUFx3_ASAP7_75t_L g7020 ( 
.A(n_6504),
.Y(n_7020)
);

AOI22xp33_ASAP7_75t_L g7021 ( 
.A1(n_5543),
.A2(n_5007),
.B1(n_5072),
.B2(n_5018),
.Y(n_7021)
);

OA21x2_ASAP7_75t_L g7022 ( 
.A1(n_6442),
.A2(n_5187),
.B(n_5185),
.Y(n_7022)
);

BUFx3_ASAP7_75t_L g7023 ( 
.A(n_6504),
.Y(n_7023)
);

OAI22xp33_ASAP7_75t_L g7024 ( 
.A1(n_6037),
.A2(n_5113),
.B1(n_5147),
.B2(n_5104),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_5674),
.Y(n_7025)
);

OAI22xp5_ASAP7_75t_L g7026 ( 
.A1(n_6430),
.A2(n_5505),
.B1(n_5523),
.B2(n_5500),
.Y(n_7026)
);

INVx3_ASAP7_75t_L g7027 ( 
.A(n_6134),
.Y(n_7027)
);

AOI21xp5_ASAP7_75t_L g7028 ( 
.A1(n_6440),
.A2(n_5362),
.B(n_5357),
.Y(n_7028)
);

AOI22xp33_ASAP7_75t_L g7029 ( 
.A1(n_5536),
.A2(n_5018),
.B1(n_5114),
.B2(n_5072),
.Y(n_7029)
);

OR2x2_ASAP7_75t_L g7030 ( 
.A(n_6190),
.B(n_5920),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_5674),
.Y(n_7031)
);

AND2x2_ASAP7_75t_L g7032 ( 
.A(n_5730),
.B(n_4623),
.Y(n_7032)
);

AO21x1_ASAP7_75t_L g7033 ( 
.A1(n_6220),
.A2(n_5399),
.B(n_4700),
.Y(n_7033)
);

NAND2xp5_ASAP7_75t_L g7034 ( 
.A(n_5901),
.B(n_4868),
.Y(n_7034)
);

AND2x2_ASAP7_75t_L g7035 ( 
.A(n_5730),
.B(n_4623),
.Y(n_7035)
);

INVx3_ASAP7_75t_L g7036 ( 
.A(n_6134),
.Y(n_7036)
);

AND2x4_ASAP7_75t_L g7037 ( 
.A(n_5594),
.B(n_5104),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_5683),
.Y(n_7038)
);

INVx4_ASAP7_75t_L g7039 ( 
.A(n_6519),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_L g7040 ( 
.A(n_5575),
.B(n_4886),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_L g7041 ( 
.A1(n_5536),
.A2(n_5114),
.B1(n_5072),
.B2(n_5113),
.Y(n_7041)
);

BUFx10_ASAP7_75t_L g7042 ( 
.A(n_5679),
.Y(n_7042)
);

OAI22xp5_ASAP7_75t_L g7043 ( 
.A1(n_6430),
.A2(n_5505),
.B1(n_5523),
.B2(n_5520),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_5683),
.Y(n_7044)
);

CKINVDCx20_ASAP7_75t_R g7045 ( 
.A(n_6600),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_5684),
.Y(n_7046)
);

OAI22xp5_ASAP7_75t_L g7047 ( 
.A1(n_6262),
.A2(n_5525),
.B1(n_5520),
.B2(n_5375),
.Y(n_7047)
);

INVx3_ASAP7_75t_L g7048 ( 
.A(n_6134),
.Y(n_7048)
);

AOI21xp5_ASAP7_75t_L g7049 ( 
.A1(n_5970),
.A2(n_6001),
.B(n_5980),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_5684),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_5696),
.Y(n_7051)
);

OAI22xp5_ASAP7_75t_L g7052 ( 
.A1(n_6262),
.A2(n_5375),
.B1(n_5376),
.B2(n_5368),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_5696),
.Y(n_7053)
);

HB1xp67_ASAP7_75t_L g7054 ( 
.A(n_6475),
.Y(n_7054)
);

INVx3_ASAP7_75t_L g7055 ( 
.A(n_6134),
.Y(n_7055)
);

NOR2xp33_ASAP7_75t_L g7056 ( 
.A(n_6019),
.B(n_4558),
.Y(n_7056)
);

INVx3_ASAP7_75t_L g7057 ( 
.A(n_6134),
.Y(n_7057)
);

INVx2_ASAP7_75t_SL g7058 ( 
.A(n_5594),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_5575),
.B(n_4886),
.Y(n_7059)
);

HAxp5_ASAP7_75t_L g7060 ( 
.A(n_5892),
.B(n_4567),
.CON(n_7060),
.SN(n_7060)
);

CKINVDCx8_ASAP7_75t_R g7061 ( 
.A(n_5583),
.Y(n_7061)
);

NAND2xp5_ASAP7_75t_L g7062 ( 
.A(n_6247),
.B(n_4902),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_SL g7063 ( 
.A(n_5947),
.B(n_5104),
.Y(n_7063)
);

HB1xp67_ASAP7_75t_L g7064 ( 
.A(n_6475),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_5698),
.Y(n_7065)
);

INVxp67_ASAP7_75t_L g7066 ( 
.A(n_6046),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6247),
.B(n_4902),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_5698),
.Y(n_7068)
);

NOR2xp33_ASAP7_75t_L g7069 ( 
.A(n_6043),
.B(n_4558),
.Y(n_7069)
);

INVx2_ASAP7_75t_SL g7070 ( 
.A(n_5594),
.Y(n_7070)
);

O2A1O1Ixp33_ASAP7_75t_L g7071 ( 
.A1(n_6376),
.A2(n_5894),
.B(n_5947),
.C(n_5964),
.Y(n_7071)
);

INVx1_ASAP7_75t_L g7072 ( 
.A(n_5710),
.Y(n_7072)
);

BUFx6f_ASAP7_75t_L g7073 ( 
.A(n_6137),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_5710),
.Y(n_7074)
);

INVxp67_ASAP7_75t_SL g7075 ( 
.A(n_6571),
.Y(n_7075)
);

AO21x2_ASAP7_75t_L g7076 ( 
.A1(n_6442),
.A2(n_5187),
.B(n_5362),
.Y(n_7076)
);

NAND2xp5_ASAP7_75t_L g7077 ( 
.A(n_6255),
.B(n_5371),
.Y(n_7077)
);

BUFx12f_ASAP7_75t_L g7078 ( 
.A(n_5632),
.Y(n_7078)
);

AND2x6_ASAP7_75t_L g7079 ( 
.A(n_5535),
.B(n_5229),
.Y(n_7079)
);

HB1xp67_ASAP7_75t_L g7080 ( 
.A(n_6497),
.Y(n_7080)
);

AND2x4_ASAP7_75t_L g7081 ( 
.A(n_5594),
.B(n_5623),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_5718),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_5718),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_5723),
.Y(n_7084)
);

AND2x4_ASAP7_75t_L g7085 ( 
.A(n_5594),
.B(n_5104),
.Y(n_7085)
);

AND2x2_ASAP7_75t_L g7086 ( 
.A(n_5721),
.B(n_4623),
.Y(n_7086)
);

AND2x4_ASAP7_75t_L g7087 ( 
.A(n_5594),
.B(n_5104),
.Y(n_7087)
);

INVxp67_ASAP7_75t_SL g7088 ( 
.A(n_6153),
.Y(n_7088)
);

AOI221xp5_ASAP7_75t_L g7089 ( 
.A1(n_5894),
.A2(n_5231),
.B1(n_5376),
.B2(n_5378),
.C(n_5368),
.Y(n_7089)
);

NAND2xp5_ASAP7_75t_L g7090 ( 
.A(n_6255),
.B(n_5371),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_SL g7091 ( 
.A(n_6064),
.B(n_5104),
.Y(n_7091)
);

INVx1_ASAP7_75t_SL g7092 ( 
.A(n_6497),
.Y(n_7092)
);

OAI22xp5_ASAP7_75t_L g7093 ( 
.A1(n_6056),
.A2(n_5378),
.B1(n_4435),
.B2(n_4503),
.Y(n_7093)
);

BUFx6f_ASAP7_75t_L g7094 ( 
.A(n_6137),
.Y(n_7094)
);

INVx1_ASAP7_75t_L g7095 ( 
.A(n_5723),
.Y(n_7095)
);

HB1xp67_ASAP7_75t_L g7096 ( 
.A(n_6497),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_SL g7097 ( 
.A(n_6006),
.B(n_5104),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_L g7098 ( 
.A(n_6264),
.B(n_5379),
.Y(n_7098)
);

AOI21xp5_ASAP7_75t_L g7099 ( 
.A1(n_5980),
.A2(n_5397),
.B(n_5495),
.Y(n_7099)
);

NOR2xp33_ASAP7_75t_L g7100 ( 
.A(n_6043),
.B(n_4663),
.Y(n_7100)
);

CKINVDCx16_ASAP7_75t_R g7101 ( 
.A(n_5986),
.Y(n_7101)
);

NOR2x1_ASAP7_75t_L g7102 ( 
.A(n_6454),
.B(n_5948),
.Y(n_7102)
);

AOI22xp33_ASAP7_75t_L g7103 ( 
.A1(n_6012),
.A2(n_5114),
.B1(n_5147),
.B2(n_5113),
.Y(n_7103)
);

INVx2_ASAP7_75t_SL g7104 ( 
.A(n_5623),
.Y(n_7104)
);

AOI22xp5_ASAP7_75t_L g7105 ( 
.A1(n_5892),
.A2(n_5114),
.B1(n_5074),
.B2(n_5113),
.Y(n_7105)
);

INVx3_ASAP7_75t_L g7106 ( 
.A(n_6137),
.Y(n_7106)
);

INVx2_ASAP7_75t_SL g7107 ( 
.A(n_5623),
.Y(n_7107)
);

NAND2xp5_ASAP7_75t_L g7108 ( 
.A(n_6002),
.B(n_5405),
.Y(n_7108)
);

INVx2_ASAP7_75t_SL g7109 ( 
.A(n_5623),
.Y(n_7109)
);

INVx3_ASAP7_75t_L g7110 ( 
.A(n_6137),
.Y(n_7110)
);

BUFx6f_ASAP7_75t_L g7111 ( 
.A(n_6137),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_5727),
.Y(n_7112)
);

NAND2xp5_ASAP7_75t_SL g7113 ( 
.A(n_6006),
.B(n_5113),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_5727),
.Y(n_7114)
);

NOR2xp33_ASAP7_75t_L g7115 ( 
.A(n_6067),
.B(n_4663),
.Y(n_7115)
);

AOI21xp5_ASAP7_75t_L g7116 ( 
.A1(n_6001),
.A2(n_5397),
.B(n_5506),
.Y(n_7116)
);

INVx5_ASAP7_75t_L g7117 ( 
.A(n_6383),
.Y(n_7117)
);

INVx2_ASAP7_75t_SL g7118 ( 
.A(n_5623),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_5738),
.Y(n_7119)
);

HB1xp67_ASAP7_75t_L g7120 ( 
.A(n_6514),
.Y(n_7120)
);

BUFx3_ASAP7_75t_L g7121 ( 
.A(n_5801),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_L g7122 ( 
.A(n_6264),
.B(n_6275),
.Y(n_7122)
);

INVx1_ASAP7_75t_SL g7123 ( 
.A(n_6514),
.Y(n_7123)
);

INVx1_ASAP7_75t_SL g7124 ( 
.A(n_6514),
.Y(n_7124)
);

OAI22xp5_ASAP7_75t_L g7125 ( 
.A1(n_6056),
.A2(n_4435),
.B1(n_4503),
.B2(n_4471),
.Y(n_7125)
);

INVx1_ASAP7_75t_L g7126 ( 
.A(n_5738),
.Y(n_7126)
);

OAI22xp5_ASAP7_75t_L g7127 ( 
.A1(n_6037),
.A2(n_4435),
.B1(n_4503),
.B2(n_4471),
.Y(n_7127)
);

NAND2xp5_ASAP7_75t_L g7128 ( 
.A(n_6275),
.B(n_4536),
.Y(n_7128)
);

CKINVDCx20_ASAP7_75t_R g7129 ( 
.A(n_5648),
.Y(n_7129)
);

A2O1A1Ixp33_ASAP7_75t_L g7130 ( 
.A1(n_6444),
.A2(n_5023),
.B(n_5026),
.C(n_4994),
.Y(n_7130)
);

O2A1O1Ixp33_ASAP7_75t_L g7131 ( 
.A1(n_5948),
.A2(n_4704),
.B(n_4730),
.C(n_4689),
.Y(n_7131)
);

INVx3_ASAP7_75t_L g7132 ( 
.A(n_6137),
.Y(n_7132)
);

INVx5_ASAP7_75t_L g7133 ( 
.A(n_6383),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_L g7134 ( 
.A(n_6303),
.B(n_4536),
.Y(n_7134)
);

CKINVDCx5p33_ASAP7_75t_R g7135 ( 
.A(n_6445),
.Y(n_7135)
);

BUFx6f_ASAP7_75t_L g7136 ( 
.A(n_6137),
.Y(n_7136)
);

O2A1O1Ixp33_ASAP7_75t_L g7137 ( 
.A1(n_5989),
.A2(n_4704),
.B(n_4730),
.C(n_4689),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_5771),
.Y(n_7138)
);

INVx6_ASAP7_75t_L g7139 ( 
.A(n_5557),
.Y(n_7139)
);

BUFx4f_ASAP7_75t_L g7140 ( 
.A(n_5656),
.Y(n_7140)
);

BUFx6f_ASAP7_75t_L g7141 ( 
.A(n_6137),
.Y(n_7141)
);

INVx4_ASAP7_75t_L g7142 ( 
.A(n_5656),
.Y(n_7142)
);

INVxp67_ASAP7_75t_SL g7143 ( 
.A(n_6153),
.Y(n_7143)
);

AOI22xp5_ASAP7_75t_L g7144 ( 
.A1(n_6067),
.A2(n_5114),
.B1(n_5074),
.B2(n_5113),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_L g7145 ( 
.A(n_6303),
.B(n_4556),
.Y(n_7145)
);

OAI22xp5_ASAP7_75t_L g7146 ( 
.A1(n_6099),
.A2(n_4435),
.B1(n_4503),
.B2(n_4471),
.Y(n_7146)
);

BUFx6f_ASAP7_75t_L g7147 ( 
.A(n_6171),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_SL g7148 ( 
.A(n_6107),
.B(n_5147),
.Y(n_7148)
);

NOR2xp33_ASAP7_75t_L g7149 ( 
.A(n_6107),
.B(n_4745),
.Y(n_7149)
);

OAI22xp5_ASAP7_75t_L g7150 ( 
.A1(n_6099),
.A2(n_4435),
.B1(n_4503),
.B2(n_4471),
.Y(n_7150)
);

AOI22xp33_ASAP7_75t_L g7151 ( 
.A1(n_6012),
.A2(n_5114),
.B1(n_5148),
.B2(n_5147),
.Y(n_7151)
);

O2A1O1Ixp5_ASAP7_75t_L g7152 ( 
.A1(n_6076),
.A2(n_5506),
.B(n_5519),
.C(n_5508),
.Y(n_7152)
);

CKINVDCx6p67_ASAP7_75t_R g7153 ( 
.A(n_5644),
.Y(n_7153)
);

OR2x6_ASAP7_75t_L g7154 ( 
.A(n_6095),
.B(n_6585),
.Y(n_7154)
);

BUFx3_ASAP7_75t_L g7155 ( 
.A(n_5801),
.Y(n_7155)
);

HB1xp67_ASAP7_75t_L g7156 ( 
.A(n_6546),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_6304),
.B(n_4556),
.Y(n_7157)
);

INVx3_ASAP7_75t_L g7158 ( 
.A(n_6171),
.Y(n_7158)
);

NOR2xp33_ASAP7_75t_L g7159 ( 
.A(n_6007),
.B(n_4745),
.Y(n_7159)
);

NAND2xp5_ASAP7_75t_L g7160 ( 
.A(n_6304),
.B(n_4556),
.Y(n_7160)
);

AND3x1_ASAP7_75t_SL g7161 ( 
.A(n_6537),
.B(n_5330),
.C(n_5447),
.Y(n_7161)
);

OAI22xp5_ASAP7_75t_L g7162 ( 
.A1(n_6372),
.A2(n_4576),
.B1(n_4471),
.B2(n_4838),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_5771),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_SL g7164 ( 
.A(n_6020),
.B(n_5147),
.Y(n_7164)
);

O2A1O1Ixp33_ASAP7_75t_L g7165 ( 
.A1(n_5989),
.A2(n_4838),
.B(n_4877),
.C(n_5414),
.Y(n_7165)
);

INVx4_ASAP7_75t_L g7166 ( 
.A(n_5656),
.Y(n_7166)
);

INVx4_ASAP7_75t_L g7167 ( 
.A(n_5647),
.Y(n_7167)
);

HB1xp67_ASAP7_75t_L g7168 ( 
.A(n_6546),
.Y(n_7168)
);

BUFx6f_ASAP7_75t_L g7169 ( 
.A(n_6171),
.Y(n_7169)
);

OAI21xp33_ASAP7_75t_L g7170 ( 
.A1(n_6020),
.A2(n_5416),
.B(n_5414),
.Y(n_7170)
);

INVxp67_ASAP7_75t_SL g7171 ( 
.A(n_6284),
.Y(n_7171)
);

OAI21xp5_ASAP7_75t_L g7172 ( 
.A1(n_6076),
.A2(n_5508),
.B(n_5506),
.Y(n_7172)
);

AOI22xp33_ASAP7_75t_L g7173 ( 
.A1(n_5573),
.A2(n_5148),
.B1(n_5147),
.B2(n_5398),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_L g7174 ( 
.A(n_6332),
.B(n_4583),
.Y(n_7174)
);

BUFx6f_ASAP7_75t_L g7175 ( 
.A(n_6171),
.Y(n_7175)
);

NAND2xp5_ASAP7_75t_L g7176 ( 
.A(n_6332),
.B(n_4583),
.Y(n_7176)
);

AOI22xp33_ASAP7_75t_L g7177 ( 
.A1(n_5573),
.A2(n_5148),
.B1(n_5147),
.B2(n_5398),
.Y(n_7177)
);

O2A1O1Ixp5_ASAP7_75t_L g7178 ( 
.A1(n_6211),
.A2(n_5951),
.B(n_5993),
.C(n_6040),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_5777),
.Y(n_7179)
);

NOR2xp33_ASAP7_75t_SL g7180 ( 
.A(n_6353),
.B(n_4462),
.Y(n_7180)
);

NAND2xp5_ASAP7_75t_L g7181 ( 
.A(n_6339),
.B(n_4583),
.Y(n_7181)
);

NOR2xp33_ASAP7_75t_R g7182 ( 
.A(n_6152),
.B(n_5330),
.Y(n_7182)
);

AOI22xp33_ASAP7_75t_SL g7183 ( 
.A1(n_6018),
.A2(n_5148),
.B1(n_5147),
.B2(n_5153),
.Y(n_7183)
);

BUFx3_ASAP7_75t_L g7184 ( 
.A(n_5801),
.Y(n_7184)
);

OAI22xp33_ASAP7_75t_L g7185 ( 
.A1(n_6286),
.A2(n_5148),
.B1(n_5023),
.B2(n_5026),
.Y(n_7185)
);

CKINVDCx11_ASAP7_75t_R g7186 ( 
.A(n_5912),
.Y(n_7186)
);

INVx2_ASAP7_75t_SL g7187 ( 
.A(n_5663),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_5777),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_5800),
.Y(n_7189)
);

NAND2xp5_ASAP7_75t_L g7190 ( 
.A(n_5913),
.B(n_4771),
.Y(n_7190)
);

INVx1_ASAP7_75t_SL g7191 ( 
.A(n_5920),
.Y(n_7191)
);

AOI21xp5_ASAP7_75t_L g7192 ( 
.A1(n_6005),
.A2(n_5519),
.B(n_5508),
.Y(n_7192)
);

NOR2xp33_ASAP7_75t_L g7193 ( 
.A(n_6007),
.B(n_4877),
.Y(n_7193)
);

AOI22xp5_ASAP7_75t_L g7194 ( 
.A1(n_6018),
.A2(n_5148),
.B1(n_5512),
.B2(n_5398),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_5800),
.Y(n_7195)
);

NAND2xp5_ASAP7_75t_SL g7196 ( 
.A(n_6033),
.B(n_5148),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_5806),
.Y(n_7197)
);

INVx3_ASAP7_75t_SL g7198 ( 
.A(n_5541),
.Y(n_7198)
);

INVx5_ASAP7_75t_L g7199 ( 
.A(n_6402),
.Y(n_7199)
);

AOI21xp5_ASAP7_75t_L g7200 ( 
.A1(n_6005),
.A2(n_5519),
.B(n_4677),
.Y(n_7200)
);

INVx1_ASAP7_75t_SL g7201 ( 
.A(n_5920),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_5806),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_5807),
.Y(n_7203)
);

OAI22xp5_ASAP7_75t_L g7204 ( 
.A1(n_6372),
.A2(n_4576),
.B1(n_5148),
.B2(n_4437),
.Y(n_7204)
);

OR2x6_ASAP7_75t_L g7205 ( 
.A(n_6095),
.B(n_4680),
.Y(n_7205)
);

BUFx6f_ASAP7_75t_L g7206 ( 
.A(n_6171),
.Y(n_7206)
);

HB1xp67_ASAP7_75t_L g7207 ( 
.A(n_6314),
.Y(n_7207)
);

NAND2xp5_ASAP7_75t_L g7208 ( 
.A(n_5929),
.B(n_4774),
.Y(n_7208)
);

NOR2x1_ASAP7_75t_L g7209 ( 
.A(n_6454),
.B(n_6288),
.Y(n_7209)
);

OAI21xp5_ASAP7_75t_L g7210 ( 
.A1(n_6211),
.A2(n_5360),
.B(n_5419),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_5807),
.Y(n_7211)
);

AOI21xp5_ASAP7_75t_L g7212 ( 
.A1(n_6015),
.A2(n_6049),
.B(n_6034),
.Y(n_7212)
);

AOI222xp33_ASAP7_75t_L g7213 ( 
.A1(n_6029),
.A2(n_5416),
.B1(n_5420),
.B2(n_5442),
.C1(n_5441),
.C2(n_5428),
.Y(n_7213)
);

AOI21xp5_ASAP7_75t_L g7214 ( 
.A1(n_6015),
.A2(n_4677),
.B(n_5199),
.Y(n_7214)
);

INVx1_ASAP7_75t_SL g7215 ( 
.A(n_5945),
.Y(n_7215)
);

CKINVDCx5p33_ASAP7_75t_R g7216 ( 
.A(n_6010),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_5816),
.Y(n_7217)
);

INVx3_ASAP7_75t_L g7218 ( 
.A(n_6171),
.Y(n_7218)
);

INVxp67_ASAP7_75t_L g7219 ( 
.A(n_6046),
.Y(n_7219)
);

NOR2xp33_ASAP7_75t_L g7220 ( 
.A(n_6187),
.B(n_5148),
.Y(n_7220)
);

BUFx6f_ASAP7_75t_L g7221 ( 
.A(n_6171),
.Y(n_7221)
);

NOR2xp33_ASAP7_75t_L g7222 ( 
.A(n_6187),
.B(n_5231),
.Y(n_7222)
);

O2A1O1Ixp5_ASAP7_75t_L g7223 ( 
.A1(n_5951),
.A2(n_4729),
.B(n_5199),
.C(n_4576),
.Y(n_7223)
);

INVx3_ASAP7_75t_L g7224 ( 
.A(n_6171),
.Y(n_7224)
);

INVx5_ASAP7_75t_L g7225 ( 
.A(n_6402),
.Y(n_7225)
);

OR2x6_ASAP7_75t_L g7226 ( 
.A(n_6095),
.B(n_4994),
.Y(n_7226)
);

AOI222xp33_ASAP7_75t_L g7227 ( 
.A1(n_6029),
.A2(n_5428),
.B1(n_5420),
.B2(n_5449),
.C1(n_5442),
.C2(n_5441),
.Y(n_7227)
);

OAI21xp5_ASAP7_75t_L g7228 ( 
.A1(n_6033),
.A2(n_5438),
.B(n_5419),
.Y(n_7228)
);

AOI22xp5_ASAP7_75t_L g7229 ( 
.A1(n_6123),
.A2(n_5512),
.B1(n_5398),
.B2(n_4920),
.Y(n_7229)
);

HB1xp67_ASAP7_75t_L g7230 ( 
.A(n_6314),
.Y(n_7230)
);

INVx2_ASAP7_75t_SL g7231 ( 
.A(n_5663),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_5816),
.Y(n_7232)
);

NOR2xp33_ASAP7_75t_L g7233 ( 
.A(n_5983),
.B(n_5231),
.Y(n_7233)
);

NAND2xp5_ASAP7_75t_L g7234 ( 
.A(n_5929),
.B(n_6339),
.Y(n_7234)
);

INVxp67_ASAP7_75t_L g7235 ( 
.A(n_6121),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_6354),
.B(n_4776),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_5817),
.Y(n_7237)
);

AOI22xp33_ASAP7_75t_L g7238 ( 
.A1(n_6032),
.A2(n_5398),
.B1(n_5233),
.B2(n_5129),
.Y(n_7238)
);

HB1xp67_ASAP7_75t_L g7239 ( 
.A(n_6322),
.Y(n_7239)
);

INVxp67_ASAP7_75t_SL g7240 ( 
.A(n_6284),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_6354),
.B(n_4776),
.Y(n_7241)
);

INVx1_ASAP7_75t_SL g7242 ( 
.A(n_5945),
.Y(n_7242)
);

NOR2xp33_ASAP7_75t_L g7243 ( 
.A(n_5983),
.B(n_5494),
.Y(n_7243)
);

INVx3_ASAP7_75t_SL g7244 ( 
.A(n_5541),
.Y(n_7244)
);

INVx1_ASAP7_75t_SL g7245 ( 
.A(n_5968),
.Y(n_7245)
);

CKINVDCx5p33_ASAP7_75t_R g7246 ( 
.A(n_6039),
.Y(n_7246)
);

NOR2xp67_ASAP7_75t_L g7247 ( 
.A(n_5754),
.B(n_4776),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_5817),
.Y(n_7248)
);

NOR2xp33_ASAP7_75t_SL g7249 ( 
.A(n_6353),
.B(n_4462),
.Y(n_7249)
);

NAND2x1_ASAP7_75t_L g7250 ( 
.A(n_5801),
.B(n_6083),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_5824),
.Y(n_7251)
);

CKINVDCx5p33_ASAP7_75t_R g7252 ( 
.A(n_6138),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_6365),
.B(n_4629),
.Y(n_7253)
);

INVx5_ASAP7_75t_L g7254 ( 
.A(n_6402),
.Y(n_7254)
);

AOI21xp5_ASAP7_75t_L g7255 ( 
.A1(n_6049),
.A2(n_4929),
.B(n_4921),
.Y(n_7255)
);

NOR2xp33_ASAP7_75t_L g7256 ( 
.A(n_5975),
.B(n_5494),
.Y(n_7256)
);

INVx1_ASAP7_75t_SL g7257 ( 
.A(n_5968),
.Y(n_7257)
);

INVx2_ASAP7_75t_SL g7258 ( 
.A(n_5663),
.Y(n_7258)
);

BUFx12f_ASAP7_75t_L g7259 ( 
.A(n_5644),
.Y(n_7259)
);

INVx2_ASAP7_75t_SL g7260 ( 
.A(n_5688),
.Y(n_7260)
);

INVx4_ASAP7_75t_L g7261 ( 
.A(n_5647),
.Y(n_7261)
);

INVx5_ASAP7_75t_L g7262 ( 
.A(n_6402),
.Y(n_7262)
);

NOR2xp33_ASAP7_75t_L g7263 ( 
.A(n_5975),
.B(n_5494),
.Y(n_7263)
);

BUFx2_ASAP7_75t_R g7264 ( 
.A(n_6282),
.Y(n_7264)
);

NAND2xp5_ASAP7_75t_L g7265 ( 
.A(n_6365),
.B(n_4629),
.Y(n_7265)
);

NOR2xp33_ASAP7_75t_L g7266 ( 
.A(n_5975),
.B(n_5494),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_5824),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_5825),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_6377),
.B(n_4629),
.Y(n_7269)
);

OAI22xp33_ASAP7_75t_L g7270 ( 
.A1(n_6286),
.A2(n_5129),
.B1(n_5026),
.B2(n_5153),
.Y(n_7270)
);

AOI221xp5_ASAP7_75t_L g7271 ( 
.A1(n_6123),
.A2(n_5449),
.B1(n_5463),
.B2(n_5460),
.C(n_5457),
.Y(n_7271)
);

BUFx10_ASAP7_75t_L g7272 ( 
.A(n_5679),
.Y(n_7272)
);

NAND2xp5_ASAP7_75t_L g7273 ( 
.A(n_6377),
.B(n_4637),
.Y(n_7273)
);

CKINVDCx20_ASAP7_75t_R g7274 ( 
.A(n_6263),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_L g7275 ( 
.A(n_6404),
.B(n_4637),
.Y(n_7275)
);

OAI21x1_ASAP7_75t_L g7276 ( 
.A1(n_6536),
.A2(n_6479),
.B(n_6468),
.Y(n_7276)
);

BUFx6f_ASAP7_75t_L g7277 ( 
.A(n_6192),
.Y(n_7277)
);

AND2x6_ASAP7_75t_L g7278 ( 
.A(n_5535),
.B(n_5229),
.Y(n_7278)
);

AOI22xp5_ASAP7_75t_L g7279 ( 
.A1(n_6032),
.A2(n_5398),
.B1(n_4928),
.B2(n_5233),
.Y(n_7279)
);

INVx3_ASAP7_75t_L g7280 ( 
.A(n_6192),
.Y(n_7280)
);

AOI221xp5_ASAP7_75t_L g7281 ( 
.A1(n_5539),
.A2(n_5457),
.B1(n_5477),
.B2(n_5463),
.C(n_5460),
.Y(n_7281)
);

BUFx6f_ASAP7_75t_L g7282 ( 
.A(n_6192),
.Y(n_7282)
);

NAND2xp5_ASAP7_75t_L g7283 ( 
.A(n_6404),
.B(n_4776),
.Y(n_7283)
);

INVxp67_ASAP7_75t_SL g7284 ( 
.A(n_5724),
.Y(n_7284)
);

HB1xp67_ASAP7_75t_L g7285 ( 
.A(n_6322),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_L g7286 ( 
.A(n_6421),
.B(n_4637),
.Y(n_7286)
);

INVx3_ASAP7_75t_L g7287 ( 
.A(n_6192),
.Y(n_7287)
);

CKINVDCx8_ASAP7_75t_R g7288 ( 
.A(n_5631),
.Y(n_7288)
);

BUFx3_ASAP7_75t_L g7289 ( 
.A(n_5801),
.Y(n_7289)
);

INVx5_ASAP7_75t_L g7290 ( 
.A(n_6402),
.Y(n_7290)
);

AOI22xp5_ASAP7_75t_L g7291 ( 
.A1(n_6160),
.A2(n_6278),
.B1(n_6218),
.B2(n_5645),
.Y(n_7291)
);

NAND2x1p5_ASAP7_75t_L g7292 ( 
.A(n_5754),
.B(n_5153),
.Y(n_7292)
);

BUFx2_ASAP7_75t_R g7293 ( 
.A(n_6282),
.Y(n_7293)
);

INVx3_ASAP7_75t_L g7294 ( 
.A(n_6192),
.Y(n_7294)
);

INVx2_ASAP7_75t_SL g7295 ( 
.A(n_5688),
.Y(n_7295)
);

AND2x4_ASAP7_75t_L g7296 ( 
.A(n_5688),
.B(n_5702),
.Y(n_7296)
);

CKINVDCx8_ASAP7_75t_R g7297 ( 
.A(n_5631),
.Y(n_7297)
);

AND2x4_ASAP7_75t_L g7298 ( 
.A(n_5688),
.B(n_5702),
.Y(n_7298)
);

O2A1O1Ixp33_ASAP7_75t_L g7299 ( 
.A1(n_5988),
.A2(n_5480),
.B(n_5483),
.C(n_5477),
.Y(n_7299)
);

INVx3_ASAP7_75t_L g7300 ( 
.A(n_6192),
.Y(n_7300)
);

INVx3_ASAP7_75t_SL g7301 ( 
.A(n_5541),
.Y(n_7301)
);

NAND2xp5_ASAP7_75t_L g7302 ( 
.A(n_6421),
.B(n_4672),
.Y(n_7302)
);

INVx5_ASAP7_75t_L g7303 ( 
.A(n_6402),
.Y(n_7303)
);

BUFx6f_ASAP7_75t_L g7304 ( 
.A(n_6192),
.Y(n_7304)
);

NAND2xp5_ASAP7_75t_L g7305 ( 
.A(n_6448),
.B(n_4778),
.Y(n_7305)
);

INVx5_ASAP7_75t_L g7306 ( 
.A(n_6402),
.Y(n_7306)
);

OR2x6_ASAP7_75t_L g7307 ( 
.A(n_6095),
.B(n_5129),
.Y(n_7307)
);

INVx3_ASAP7_75t_L g7308 ( 
.A(n_6192),
.Y(n_7308)
);

AOI22xp5_ASAP7_75t_L g7309 ( 
.A1(n_6160),
.A2(n_5398),
.B1(n_4928),
.B2(n_5233),
.Y(n_7309)
);

AOI21xp5_ASAP7_75t_L g7310 ( 
.A1(n_6053),
.A2(n_4929),
.B(n_4921),
.Y(n_7310)
);

O2A1O1Ixp5_ASAP7_75t_L g7311 ( 
.A1(n_5993),
.A2(n_4729),
.B(n_4576),
.C(n_5197),
.Y(n_7311)
);

INVx3_ASAP7_75t_L g7312 ( 
.A(n_6196),
.Y(n_7312)
);

INVx3_ASAP7_75t_L g7313 ( 
.A(n_6196),
.Y(n_7313)
);

OR2x6_ASAP7_75t_L g7314 ( 
.A(n_6585),
.B(n_5129),
.Y(n_7314)
);

OAI221xp5_ASAP7_75t_L g7315 ( 
.A1(n_6048),
.A2(n_5480),
.B1(n_5497),
.B2(n_5496),
.C(n_5483),
.Y(n_7315)
);

BUFx8_ASAP7_75t_SL g7316 ( 
.A(n_5912),
.Y(n_7316)
);

INVx3_ASAP7_75t_L g7317 ( 
.A(n_6196),
.Y(n_7317)
);

INVx4_ASAP7_75t_SL g7318 ( 
.A(n_5801),
.Y(n_7318)
);

NOR3xp33_ASAP7_75t_L g7319 ( 
.A(n_5545),
.B(n_5497),
.C(n_5496),
.Y(n_7319)
);

HB1xp67_ASAP7_75t_L g7320 ( 
.A(n_6343),
.Y(n_7320)
);

INVx4_ASAP7_75t_L g7321 ( 
.A(n_5647),
.Y(n_7321)
);

BUFx3_ASAP7_75t_L g7322 ( 
.A(n_5801),
.Y(n_7322)
);

AOI22xp5_ASAP7_75t_SL g7323 ( 
.A1(n_6121),
.A2(n_4748),
.B1(n_4608),
.B2(n_4865),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_6448),
.B(n_4778),
.Y(n_7324)
);

AOI21xp5_ASAP7_75t_L g7325 ( 
.A1(n_6053),
.A2(n_4921),
.B(n_5153),
.Y(n_7325)
);

INVx2_ASAP7_75t_SL g7326 ( 
.A(n_5702),
.Y(n_7326)
);

INVx3_ASAP7_75t_L g7327 ( 
.A(n_6196),
.Y(n_7327)
);

INVxp67_ASAP7_75t_SL g7328 ( 
.A(n_5724),
.Y(n_7328)
);

NAND2x1p5_ASAP7_75t_L g7329 ( 
.A(n_5754),
.B(n_5829),
.Y(n_7329)
);

INVx2_ASAP7_75t_SL g7330 ( 
.A(n_5702),
.Y(n_7330)
);

NAND2x2_ASAP7_75t_L g7331 ( 
.A(n_5535),
.B(n_5556),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_6462),
.B(n_4778),
.Y(n_7332)
);

INVx3_ASAP7_75t_L g7333 ( 
.A(n_6196),
.Y(n_7333)
);

AO21x2_ASAP7_75t_L g7334 ( 
.A1(n_6468),
.A2(n_4425),
.B(n_4424),
.Y(n_7334)
);

INVx4_ASAP7_75t_L g7335 ( 
.A(n_5647),
.Y(n_7335)
);

AND2x2_ASAP7_75t_L g7336 ( 
.A(n_5784),
.B(n_5770),
.Y(n_7336)
);

NOR2xp33_ASAP7_75t_L g7337 ( 
.A(n_5975),
.B(n_5150),
.Y(n_7337)
);

INVx2_ASAP7_75t_SL g7338 ( 
.A(n_5702),
.Y(n_7338)
);

AND3x2_ASAP7_75t_L g7339 ( 
.A(n_6447),
.B(n_5475),
.C(n_5474),
.Y(n_7339)
);

OAI22xp5_ASAP7_75t_L g7340 ( 
.A1(n_6048),
.A2(n_4576),
.B1(n_4437),
.B2(n_4550),
.Y(n_7340)
);

OAI22xp5_ASAP7_75t_L g7341 ( 
.A1(n_6401),
.A2(n_4437),
.B1(n_4550),
.B2(n_4487),
.Y(n_7341)
);

AND2x4_ASAP7_75t_L g7342 ( 
.A(n_5702),
.B(n_5708),
.Y(n_7342)
);

AOI21xp5_ASAP7_75t_L g7343 ( 
.A1(n_6054),
.A2(n_5153),
.B(n_4662),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_L g7344 ( 
.A(n_6462),
.B(n_4778),
.Y(n_7344)
);

AOI22xp5_ASAP7_75t_L g7345 ( 
.A1(n_6278),
.A2(n_5398),
.B1(n_5499),
.B2(n_4448),
.Y(n_7345)
);

BUFx12f_ASAP7_75t_L g7346 ( 
.A(n_5798),
.Y(n_7346)
);

BUFx6f_ASAP7_75t_L g7347 ( 
.A(n_6196),
.Y(n_7347)
);

BUFx3_ASAP7_75t_L g7348 ( 
.A(n_5801),
.Y(n_7348)
);

AOI22xp5_ASAP7_75t_L g7349 ( 
.A1(n_6218),
.A2(n_5398),
.B1(n_5499),
.B2(n_4448),
.Y(n_7349)
);

BUFx6f_ASAP7_75t_L g7350 ( 
.A(n_6196),
.Y(n_7350)
);

BUFx12f_ASAP7_75t_L g7351 ( 
.A(n_5798),
.Y(n_7351)
);

AOI22xp5_ASAP7_75t_L g7352 ( 
.A1(n_5645),
.A2(n_5398),
.B1(n_4448),
.B2(n_5330),
.Y(n_7352)
);

BUFx3_ASAP7_75t_L g7353 ( 
.A(n_6083),
.Y(n_7353)
);

NAND2xp5_ASAP7_75t_L g7354 ( 
.A(n_6511),
.B(n_4790),
.Y(n_7354)
);

CKINVDCx11_ASAP7_75t_R g7355 ( 
.A(n_5912),
.Y(n_7355)
);

NAND2xp5_ASAP7_75t_L g7356 ( 
.A(n_6511),
.B(n_6531),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_6531),
.B(n_4672),
.Y(n_7357)
);

NOR2xp33_ASAP7_75t_L g7358 ( 
.A(n_6424),
.B(n_5150),
.Y(n_7358)
);

AOI22xp5_ASAP7_75t_L g7359 ( 
.A1(n_6359),
.A2(n_5398),
.B1(n_4448),
.B2(n_5330),
.Y(n_7359)
);

INVx4_ASAP7_75t_L g7360 ( 
.A(n_5647),
.Y(n_7360)
);

NAND2xp5_ASAP7_75t_L g7361 ( 
.A(n_6582),
.B(n_4672),
.Y(n_7361)
);

NAND2xp5_ASAP7_75t_L g7362 ( 
.A(n_6582),
.B(n_4687),
.Y(n_7362)
);

HB1xp67_ASAP7_75t_L g7363 ( 
.A(n_6343),
.Y(n_7363)
);

INVx1_ASAP7_75t_SL g7364 ( 
.A(n_6270),
.Y(n_7364)
);

AOI22xp33_ASAP7_75t_L g7365 ( 
.A1(n_5545),
.A2(n_5330),
.B1(n_5153),
.B2(n_4550),
.Y(n_7365)
);

BUFx6f_ASAP7_75t_L g7366 ( 
.A(n_6197),
.Y(n_7366)
);

NOR3xp33_ASAP7_75t_L g7367 ( 
.A(n_5598),
.B(n_4967),
.C(n_4933),
.Y(n_7367)
);

HB1xp67_ASAP7_75t_L g7368 ( 
.A(n_6344),
.Y(n_7368)
);

AOI22xp33_ASAP7_75t_L g7369 ( 
.A1(n_5598),
.A2(n_5153),
.B1(n_4487),
.B2(n_5150),
.Y(n_7369)
);

AOI22xp33_ASAP7_75t_L g7370 ( 
.A1(n_5605),
.A2(n_5153),
.B1(n_4487),
.B2(n_5150),
.Y(n_7370)
);

BUFx6f_ASAP7_75t_L g7371 ( 
.A(n_6197),
.Y(n_7371)
);

HB1xp67_ASAP7_75t_L g7372 ( 
.A(n_6344),
.Y(n_7372)
);

AOI22xp5_ASAP7_75t_L g7373 ( 
.A1(n_6359),
.A2(n_5250),
.B1(n_5262),
.B2(n_5150),
.Y(n_7373)
);

CKINVDCx5p33_ASAP7_75t_R g7374 ( 
.A(n_5933),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_6588),
.B(n_4687),
.Y(n_7375)
);

INVx6_ASAP7_75t_L g7376 ( 
.A(n_5557),
.Y(n_7376)
);

OAI22xp5_ASAP7_75t_L g7377 ( 
.A1(n_6401),
.A2(n_5060),
.B1(n_5071),
.B2(n_5040),
.Y(n_7377)
);

NAND2xp5_ASAP7_75t_L g7378 ( 
.A(n_6588),
.B(n_4687),
.Y(n_7378)
);

NOR2xp33_ASAP7_75t_L g7379 ( 
.A(n_6424),
.B(n_5150),
.Y(n_7379)
);

AOI21xp5_ASAP7_75t_L g7380 ( 
.A1(n_6054),
.A2(n_4662),
.B(n_4651),
.Y(n_7380)
);

INVxp67_ASAP7_75t_L g7381 ( 
.A(n_6281),
.Y(n_7381)
);

OAI22xp5_ASAP7_75t_L g7382 ( 
.A1(n_5986),
.A2(n_5060),
.B1(n_5071),
.B2(n_5040),
.Y(n_7382)
);

NOR2x1_ASAP7_75t_R g7383 ( 
.A(n_5798),
.B(n_4462),
.Y(n_7383)
);

BUFx3_ASAP7_75t_L g7384 ( 
.A(n_6083),
.Y(n_7384)
);

CKINVDCx5p33_ASAP7_75t_R g7385 ( 
.A(n_5933),
.Y(n_7385)
);

OAI22xp5_ASAP7_75t_L g7386 ( 
.A1(n_5986),
.A2(n_5060),
.B1(n_5071),
.B2(n_5040),
.Y(n_7386)
);

OAI22xp5_ASAP7_75t_L g7387 ( 
.A1(n_6346),
.A2(n_5090),
.B1(n_5095),
.B2(n_5076),
.Y(n_7387)
);

NAND2xp5_ASAP7_75t_SL g7388 ( 
.A(n_6251),
.B(n_5171),
.Y(n_7388)
);

BUFx3_ASAP7_75t_L g7389 ( 
.A(n_6083),
.Y(n_7389)
);

AND2x2_ASAP7_75t_L g7390 ( 
.A(n_5784),
.B(n_5793),
.Y(n_7390)
);

CKINVDCx20_ASAP7_75t_R g7391 ( 
.A(n_6263),
.Y(n_7391)
);

AOI22xp33_ASAP7_75t_L g7392 ( 
.A1(n_5605),
.A2(n_5250),
.B1(n_5262),
.B2(n_5237),
.Y(n_7392)
);

OAI21x1_ASAP7_75t_L g7393 ( 
.A1(n_6479),
.A2(n_4795),
.B(n_4790),
.Y(n_7393)
);

BUFx4_ASAP7_75t_SL g7394 ( 
.A(n_5744),
.Y(n_7394)
);

AOI21xp33_ASAP7_75t_SL g7395 ( 
.A1(n_6140),
.A2(n_5365),
.B(n_5184),
.Y(n_7395)
);

BUFx12f_ASAP7_75t_L g7396 ( 
.A(n_6428),
.Y(n_7396)
);

CKINVDCx5p33_ASAP7_75t_R g7397 ( 
.A(n_5933),
.Y(n_7397)
);

BUFx10_ASAP7_75t_L g7398 ( 
.A(n_5679),
.Y(n_7398)
);

NAND2xp5_ASAP7_75t_L g7399 ( 
.A(n_6607),
.B(n_4790),
.Y(n_7399)
);

AOI22xp5_ASAP7_75t_L g7400 ( 
.A1(n_6074),
.A2(n_5262),
.B1(n_5250),
.B2(n_4638),
.Y(n_7400)
);

OAI22xp5_ASAP7_75t_L g7401 ( 
.A1(n_6346),
.A2(n_6294),
.B1(n_5988),
.B2(n_5639),
.Y(n_7401)
);

HAxp5_ASAP7_75t_L g7402 ( 
.A(n_6537),
.B(n_5513),
.CON(n_7402),
.SN(n_7402)
);

INVx2_ASAP7_75t_SL g7403 ( 
.A(n_5708),
.Y(n_7403)
);

CKINVDCx5p33_ASAP7_75t_R g7404 ( 
.A(n_5946),
.Y(n_7404)
);

CKINVDCx8_ASAP7_75t_R g7405 ( 
.A(n_5729),
.Y(n_7405)
);

CKINVDCx5p33_ASAP7_75t_R g7406 ( 
.A(n_5946),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_L g7407 ( 
.A(n_6607),
.B(n_4790),
.Y(n_7407)
);

CKINVDCx20_ASAP7_75t_R g7408 ( 
.A(n_6458),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_6591),
.B(n_6594),
.Y(n_7409)
);

NAND2xp5_ASAP7_75t_L g7410 ( 
.A(n_6591),
.B(n_4795),
.Y(n_7410)
);

AOI21xp5_ASAP7_75t_L g7411 ( 
.A1(n_6060),
.A2(n_4665),
.B(n_4662),
.Y(n_7411)
);

NOR2xp33_ASAP7_75t_L g7412 ( 
.A(n_6439),
.B(n_6011),
.Y(n_7412)
);

OAI22xp33_ASAP7_75t_L g7413 ( 
.A1(n_5629),
.A2(n_5230),
.B1(n_5268),
.B2(n_5229),
.Y(n_7413)
);

INVx2_ASAP7_75t_SL g7414 ( 
.A(n_5768),
.Y(n_7414)
);

OAI21xp33_ASAP7_75t_SL g7415 ( 
.A1(n_5939),
.A2(n_5090),
.B(n_5076),
.Y(n_7415)
);

CKINVDCx5p33_ASAP7_75t_R g7416 ( 
.A(n_5946),
.Y(n_7416)
);

NAND2xp5_ASAP7_75t_L g7417 ( 
.A(n_6594),
.B(n_4795),
.Y(n_7417)
);

AOI22xp5_ASAP7_75t_L g7418 ( 
.A1(n_6074),
.A2(n_6201),
.B1(n_6185),
.B2(n_5977),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_L g7419 ( 
.A(n_6610),
.B(n_6513),
.Y(n_7419)
);

AO32x2_ASAP7_75t_L g7420 ( 
.A1(n_6205),
.A2(n_4927),
.A3(n_4932),
.B1(n_4871),
.B2(n_4710),
.Y(n_7420)
);

NAND2xp5_ASAP7_75t_L g7421 ( 
.A(n_6569),
.B(n_4809),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_6569),
.B(n_4809),
.Y(n_7422)
);

INVx2_ASAP7_75t_SL g7423 ( 
.A(n_5768),
.Y(n_7423)
);

AOI22xp5_ASAP7_75t_L g7424 ( 
.A1(n_6185),
.A2(n_5262),
.B1(n_5250),
.B2(n_4638),
.Y(n_7424)
);

INVx1_ASAP7_75t_SL g7425 ( 
.A(n_6270),
.Y(n_7425)
);

BUFx3_ASAP7_75t_L g7426 ( 
.A(n_6083),
.Y(n_7426)
);

NOR4xp25_ASAP7_75t_L g7427 ( 
.A(n_6258),
.B(n_6251),
.C(n_6047),
.D(n_6052),
.Y(n_7427)
);

INVx2_ASAP7_75t_SL g7428 ( 
.A(n_5768),
.Y(n_7428)
);

INVx5_ASAP7_75t_L g7429 ( 
.A(n_6432),
.Y(n_7429)
);

O2A1O1Ixp33_ASAP7_75t_SL g7430 ( 
.A1(n_5692),
.A2(n_4729),
.B(n_5184),
.C(n_4953),
.Y(n_7430)
);

BUFx6f_ASAP7_75t_L g7431 ( 
.A(n_6216),
.Y(n_7431)
);

NAND2xp5_ASAP7_75t_SL g7432 ( 
.A(n_6493),
.B(n_5171),
.Y(n_7432)
);

NAND2x1p5_ASAP7_75t_L g7433 ( 
.A(n_5754),
.B(n_4462),
.Y(n_7433)
);

INVx1_ASAP7_75t_SL g7434 ( 
.A(n_6270),
.Y(n_7434)
);

AOI21xp5_ASAP7_75t_L g7435 ( 
.A1(n_6078),
.A2(n_4665),
.B(n_4662),
.Y(n_7435)
);

CKINVDCx5p33_ASAP7_75t_R g7436 ( 
.A(n_5753),
.Y(n_7436)
);

BUFx6f_ASAP7_75t_L g7437 ( 
.A(n_6216),
.Y(n_7437)
);

INVx4_ASAP7_75t_L g7438 ( 
.A(n_5647),
.Y(n_7438)
);

CKINVDCx5p33_ASAP7_75t_R g7439 ( 
.A(n_5775),
.Y(n_7439)
);

NAND2x1p5_ASAP7_75t_L g7440 ( 
.A(n_5829),
.B(n_4462),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_L g7441 ( 
.A(n_6579),
.B(n_4809),
.Y(n_7441)
);

INVx2_ASAP7_75t_SL g7442 ( 
.A(n_5768),
.Y(n_7442)
);

NOR2xp33_ASAP7_75t_L g7443 ( 
.A(n_6439),
.B(n_5250),
.Y(n_7443)
);

O2A1O1Ixp33_ASAP7_75t_L g7444 ( 
.A1(n_5617),
.A2(n_5184),
.B(n_5365),
.C(n_5251),
.Y(n_7444)
);

AOI21xp5_ASAP7_75t_L g7445 ( 
.A1(n_6078),
.A2(n_4665),
.B(n_4662),
.Y(n_7445)
);

OA21x2_ASAP7_75t_L g7446 ( 
.A1(n_6592),
.A2(n_4831),
.B(n_4813),
.Y(n_7446)
);

AOI22xp33_ASAP7_75t_L g7447 ( 
.A1(n_6294),
.A2(n_5250),
.B1(n_5262),
.B2(n_5237),
.Y(n_7447)
);

OAI22xp33_ASAP7_75t_L g7448 ( 
.A1(n_5629),
.A2(n_5268),
.B1(n_5314),
.B2(n_5230),
.Y(n_7448)
);

NOR2x1_ASAP7_75t_L g7449 ( 
.A(n_6288),
.B(n_5179),
.Y(n_7449)
);

O2A1O1Ixp33_ASAP7_75t_L g7450 ( 
.A1(n_5617),
.A2(n_6040),
.B(n_6085),
.C(n_6258),
.Y(n_7450)
);

INVx1_ASAP7_75t_SL g7451 ( 
.A(n_5932),
.Y(n_7451)
);

CKINVDCx5p33_ASAP7_75t_R g7452 ( 
.A(n_5805),
.Y(n_7452)
);

BUFx6f_ASAP7_75t_L g7453 ( 
.A(n_6236),
.Y(n_7453)
);

CKINVDCx20_ASAP7_75t_R g7454 ( 
.A(n_6458),
.Y(n_7454)
);

AOI22xp33_ASAP7_75t_L g7455 ( 
.A1(n_5639),
.A2(n_5262),
.B1(n_5291),
.B2(n_5237),
.Y(n_7455)
);

AOI22xp33_ASAP7_75t_L g7456 ( 
.A1(n_6140),
.A2(n_5300),
.B1(n_5304),
.B2(n_5291),
.Y(n_7456)
);

NAND2xp5_ASAP7_75t_L g7457 ( 
.A(n_6610),
.B(n_6513),
.Y(n_7457)
);

BUFx2_ASAP7_75t_SL g7458 ( 
.A(n_6490),
.Y(n_7458)
);

AOI21xp5_ASAP7_75t_L g7459 ( 
.A1(n_6091),
.A2(n_4665),
.B(n_4662),
.Y(n_7459)
);

INVx4_ASAP7_75t_L g7460 ( 
.A(n_5647),
.Y(n_7460)
);

BUFx6f_ASAP7_75t_L g7461 ( 
.A(n_6236),
.Y(n_7461)
);

AOI22xp33_ASAP7_75t_L g7462 ( 
.A1(n_6170),
.A2(n_6162),
.B1(n_6201),
.B2(n_5572),
.Y(n_7462)
);

AOI22xp33_ASAP7_75t_L g7463 ( 
.A1(n_6170),
.A2(n_5300),
.B1(n_5304),
.B2(n_5291),
.Y(n_7463)
);

BUFx3_ASAP7_75t_L g7464 ( 
.A(n_6083),
.Y(n_7464)
);

BUFx3_ASAP7_75t_L g7465 ( 
.A(n_6083),
.Y(n_7465)
);

INVx2_ASAP7_75t_SL g7466 ( 
.A(n_5779),
.Y(n_7466)
);

HB1xp67_ASAP7_75t_L g7467 ( 
.A(n_6348),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_6545),
.B(n_4813),
.Y(n_7468)
);

CKINVDCx5p33_ASAP7_75t_R g7469 ( 
.A(n_6274),
.Y(n_7469)
);

AOI21x1_ASAP7_75t_L g7470 ( 
.A1(n_6486),
.A2(n_5438),
.B(n_5474),
.Y(n_7470)
);

NOR2xp33_ASAP7_75t_L g7471 ( 
.A(n_6011),
.B(n_4650),
.Y(n_7471)
);

CKINVDCx20_ASAP7_75t_R g7472 ( 
.A(n_6306),
.Y(n_7472)
);

NAND2xp5_ASAP7_75t_L g7473 ( 
.A(n_6545),
.B(n_4831),
.Y(n_7473)
);

OR2x6_ASAP7_75t_SL g7474 ( 
.A(n_6309),
.B(n_5049),
.Y(n_7474)
);

NAND3xp33_ASAP7_75t_L g7475 ( 
.A(n_6224),
.B(n_5205),
.C(n_5202),
.Y(n_7475)
);

CKINVDCx5p33_ASAP7_75t_R g7476 ( 
.A(n_6360),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_SL g7477 ( 
.A(n_6493),
.B(n_5171),
.Y(n_7477)
);

AOI22xp33_ASAP7_75t_L g7478 ( 
.A1(n_6162),
.A2(n_5304),
.B1(n_5300),
.B2(n_5239),
.Y(n_7478)
);

OR2x6_ASAP7_75t_SL g7479 ( 
.A(n_6309),
.B(n_5049),
.Y(n_7479)
);

NAND2xp5_ASAP7_75t_L g7480 ( 
.A(n_6579),
.B(n_4831),
.Y(n_7480)
);

BUFx6f_ASAP7_75t_L g7481 ( 
.A(n_6236),
.Y(n_7481)
);

OAI21xp5_ASAP7_75t_L g7482 ( 
.A1(n_5939),
.A2(n_5249),
.B(n_5238),
.Y(n_7482)
);

INVx8_ASAP7_75t_L g7483 ( 
.A(n_5842),
.Y(n_7483)
);

AOI22xp33_ASAP7_75t_L g7484 ( 
.A1(n_5572),
.A2(n_5239),
.B1(n_5266),
.B2(n_5242),
.Y(n_7484)
);

AOI22xp33_ASAP7_75t_SL g7485 ( 
.A1(n_6482),
.A2(n_5431),
.B1(n_5268),
.B2(n_5314),
.Y(n_7485)
);

NOR2xp67_ASAP7_75t_L g7486 ( 
.A(n_5829),
.B(n_4832),
.Y(n_7486)
);

AOI21xp5_ASAP7_75t_L g7487 ( 
.A1(n_6091),
.A2(n_4675),
.B(n_4665),
.Y(n_7487)
);

AOI222xp33_ASAP7_75t_L g7488 ( 
.A1(n_6277),
.A2(n_5549),
.B1(n_5539),
.B2(n_5634),
.C1(n_5720),
.C2(n_5685),
.Y(n_7488)
);

BUFx3_ASAP7_75t_L g7489 ( 
.A(n_6083),
.Y(n_7489)
);

BUFx8_ASAP7_75t_SL g7490 ( 
.A(n_5973),
.Y(n_7490)
);

NAND2xp5_ASAP7_75t_L g7491 ( 
.A(n_6599),
.B(n_4832),
.Y(n_7491)
);

BUFx6f_ASAP7_75t_L g7492 ( 
.A(n_6236),
.Y(n_7492)
);

BUFx4_ASAP7_75t_SL g7493 ( 
.A(n_6406),
.Y(n_7493)
);

AOI22xp33_ASAP7_75t_SL g7494 ( 
.A1(n_6482),
.A2(n_5431),
.B1(n_5268),
.B2(n_5314),
.Y(n_7494)
);

AOI21xp5_ASAP7_75t_L g7495 ( 
.A1(n_6104),
.A2(n_4679),
.B(n_4675),
.Y(n_7495)
);

NAND2xp5_ASAP7_75t_SL g7496 ( 
.A(n_6030),
.B(n_5171),
.Y(n_7496)
);

NAND2xp33_ASAP7_75t_L g7497 ( 
.A(n_6570),
.B(n_4865),
.Y(n_7497)
);

NOR2xp33_ASAP7_75t_L g7498 ( 
.A(n_6094),
.B(n_4650),
.Y(n_7498)
);

AOI22xp33_ASAP7_75t_L g7499 ( 
.A1(n_6145),
.A2(n_5239),
.B1(n_5266),
.B2(n_5242),
.Y(n_7499)
);

BUFx12f_ASAP7_75t_L g7500 ( 
.A(n_6038),
.Y(n_7500)
);

AND2x2_ASAP7_75t_L g7501 ( 
.A(n_5822),
.B(n_5833),
.Y(n_7501)
);

AOI22xp5_ASAP7_75t_L g7502 ( 
.A1(n_5974),
.A2(n_4644),
.B1(n_4654),
.B2(n_4638),
.Y(n_7502)
);

OAI22xp5_ASAP7_75t_L g7503 ( 
.A1(n_6364),
.A2(n_5090),
.B1(n_5095),
.B2(n_5076),
.Y(n_7503)
);

BUFx3_ASAP7_75t_L g7504 ( 
.A(n_6409),
.Y(n_7504)
);

BUFx3_ASAP7_75t_L g7505 ( 
.A(n_6409),
.Y(n_7505)
);

AOI21xp5_ASAP7_75t_L g7506 ( 
.A1(n_6104),
.A2(n_4679),
.B(n_4675),
.Y(n_7506)
);

NOR2xp33_ASAP7_75t_L g7507 ( 
.A(n_6094),
.B(n_4650),
.Y(n_7507)
);

BUFx3_ASAP7_75t_L g7508 ( 
.A(n_6409),
.Y(n_7508)
);

A2O1A1Ixp33_ASAP7_75t_L g7509 ( 
.A1(n_5874),
.A2(n_4472),
.B(n_5193),
.C(n_5179),
.Y(n_7509)
);

AND2x4_ASAP7_75t_L g7510 ( 
.A(n_5779),
.B(n_5787),
.Y(n_7510)
);

NOR2xp67_ASAP7_75t_L g7511 ( 
.A(n_5829),
.B(n_4834),
.Y(n_7511)
);

INVxp67_ASAP7_75t_L g7512 ( 
.A(n_6281),
.Y(n_7512)
);

AOI222xp33_ASAP7_75t_L g7513 ( 
.A1(n_6277),
.A2(n_5219),
.B1(n_5202),
.B2(n_5223),
.C1(n_5216),
.C2(n_5205),
.Y(n_7513)
);

BUFx4_ASAP7_75t_SL g7514 ( 
.A(n_6261),
.Y(n_7514)
);

BUFx6f_ASAP7_75t_L g7515 ( 
.A(n_6252),
.Y(n_7515)
);

AOI22xp33_ASAP7_75t_L g7516 ( 
.A1(n_6145),
.A2(n_5242),
.B1(n_5275),
.B2(n_5266),
.Y(n_7516)
);

O2A1O1Ixp5_ASAP7_75t_L g7517 ( 
.A1(n_6244),
.A2(n_5287),
.B(n_5363),
.C(n_5197),
.Y(n_7517)
);

OAI22xp33_ASAP7_75t_L g7518 ( 
.A1(n_5624),
.A2(n_5268),
.B1(n_5314),
.B2(n_5230),
.Y(n_7518)
);

AOI22xp5_ASAP7_75t_L g7519 ( 
.A1(n_5974),
.A2(n_4654),
.B1(n_4660),
.B2(n_4644),
.Y(n_7519)
);

A2O1A1Ixp33_ASAP7_75t_L g7520 ( 
.A1(n_5874),
.A2(n_4472),
.B(n_5193),
.C(n_5179),
.Y(n_7520)
);

BUFx3_ASAP7_75t_L g7521 ( 
.A(n_6409),
.Y(n_7521)
);

NAND2xp5_ASAP7_75t_L g7522 ( 
.A(n_6599),
.B(n_4834),
.Y(n_7522)
);

AND2x4_ASAP7_75t_SL g7523 ( 
.A(n_6157),
.B(n_5230),
.Y(n_7523)
);

INVx1_ASAP7_75t_SL g7524 ( 
.A(n_5932),
.Y(n_7524)
);

CKINVDCx20_ASAP7_75t_R g7525 ( 
.A(n_6358),
.Y(n_7525)
);

BUFx3_ASAP7_75t_L g7526 ( 
.A(n_6409),
.Y(n_7526)
);

BUFx6f_ASAP7_75t_L g7527 ( 
.A(n_6252),
.Y(n_7527)
);

INVx2_ASAP7_75t_SL g7528 ( 
.A(n_5779),
.Y(n_7528)
);

AOI22xp5_ASAP7_75t_L g7529 ( 
.A1(n_5977),
.A2(n_4654),
.B1(n_4660),
.B2(n_4644),
.Y(n_7529)
);

AOI22xp33_ASAP7_75t_L g7530 ( 
.A1(n_6364),
.A2(n_5289),
.B1(n_5275),
.B2(n_5249),
.Y(n_7530)
);

OAI21xp33_ASAP7_75t_L g7531 ( 
.A1(n_6085),
.A2(n_6115),
.B(n_5624),
.Y(n_7531)
);

BUFx3_ASAP7_75t_L g7532 ( 
.A(n_6409),
.Y(n_7532)
);

CKINVDCx8_ASAP7_75t_R g7533 ( 
.A(n_5729),
.Y(n_7533)
);

INVxp67_ASAP7_75t_SL g7534 ( 
.A(n_5985),
.Y(n_7534)
);

BUFx6f_ASAP7_75t_L g7535 ( 
.A(n_6252),
.Y(n_7535)
);

INVxp67_ASAP7_75t_L g7536 ( 
.A(n_6281),
.Y(n_7536)
);

AOI22xp33_ASAP7_75t_L g7537 ( 
.A1(n_6122),
.A2(n_5289),
.B1(n_5275),
.B2(n_5249),
.Y(n_7537)
);

OAI22xp5_ASAP7_75t_L g7538 ( 
.A1(n_6271),
.A2(n_5099),
.B1(n_5103),
.B2(n_5095),
.Y(n_7538)
);

AOI22xp5_ASAP7_75t_L g7539 ( 
.A1(n_5685),
.A2(n_4654),
.B1(n_4660),
.B2(n_4644),
.Y(n_7539)
);

OAI22xp33_ASAP7_75t_L g7540 ( 
.A1(n_6447),
.A2(n_5268),
.B1(n_5314),
.B2(n_5230),
.Y(n_7540)
);

AOI21xp5_ASAP7_75t_L g7541 ( 
.A1(n_6106),
.A2(n_4679),
.B(n_4675),
.Y(n_7541)
);

AOI22xp33_ASAP7_75t_L g7542 ( 
.A1(n_6122),
.A2(n_5289),
.B1(n_5249),
.B2(n_5260),
.Y(n_7542)
);

BUFx3_ASAP7_75t_L g7543 ( 
.A(n_6409),
.Y(n_7543)
);

NAND2xp5_ASAP7_75t_SL g7544 ( 
.A(n_6030),
.B(n_5171),
.Y(n_7544)
);

AOI22xp5_ASAP7_75t_L g7545 ( 
.A1(n_5720),
.A2(n_4654),
.B1(n_4660),
.B2(n_4644),
.Y(n_7545)
);

NAND2x1p5_ASAP7_75t_L g7546 ( 
.A(n_5829),
.B(n_4462),
.Y(n_7546)
);

AND2x2_ASAP7_75t_SL g7547 ( 
.A(n_6000),
.B(n_4472),
.Y(n_7547)
);

INVx1_ASAP7_75t_SL g7548 ( 
.A(n_5932),
.Y(n_7548)
);

BUFx3_ASAP7_75t_L g7549 ( 
.A(n_6409),
.Y(n_7549)
);

NOR2xp67_ASAP7_75t_SL g7550 ( 
.A(n_5701),
.B(n_5707),
.Y(n_7550)
);

CKINVDCx5p33_ASAP7_75t_R g7551 ( 
.A(n_5990),
.Y(n_7551)
);

NOR2xp33_ASAP7_75t_L g7552 ( 
.A(n_6231),
.B(n_4650),
.Y(n_7552)
);

NOR2xp33_ASAP7_75t_L g7553 ( 
.A(n_6231),
.B(n_4650),
.Y(n_7553)
);

AOI22xp5_ASAP7_75t_L g7554 ( 
.A1(n_5797),
.A2(n_4660),
.B1(n_4668),
.B2(n_4654),
.Y(n_7554)
);

CKINVDCx5p33_ASAP7_75t_R g7555 ( 
.A(n_5991),
.Y(n_7555)
);

AOI22xp5_ASAP7_75t_L g7556 ( 
.A1(n_5797),
.A2(n_4674),
.B1(n_4691),
.B2(n_4668),
.Y(n_7556)
);

CKINVDCx5p33_ASAP7_75t_R g7557 ( 
.A(n_5903),
.Y(n_7557)
);

AOI21xp5_ASAP7_75t_L g7558 ( 
.A1(n_6106),
.A2(n_4679),
.B(n_4675),
.Y(n_7558)
);

INVxp67_ASAP7_75t_SL g7559 ( 
.A(n_5985),
.Y(n_7559)
);

CKINVDCx5p33_ASAP7_75t_R g7560 ( 
.A(n_5950),
.Y(n_7560)
);

NOR2x1_ASAP7_75t_L g7561 ( 
.A(n_6292),
.B(n_5193),
.Y(n_7561)
);

OAI22xp5_ASAP7_75t_L g7562 ( 
.A1(n_6271),
.A2(n_5103),
.B1(n_5115),
.B2(n_5099),
.Y(n_7562)
);

CKINVDCx5p33_ASAP7_75t_R g7563 ( 
.A(n_5955),
.Y(n_7563)
);

BUFx4f_ASAP7_75t_L g7564 ( 
.A(n_5860),
.Y(n_7564)
);

NOR2x1_ASAP7_75t_L g7565 ( 
.A(n_6292),
.B(n_5193),
.Y(n_7565)
);

OAI22xp5_ASAP7_75t_L g7566 ( 
.A1(n_6500),
.A2(n_5103),
.B1(n_5115),
.B2(n_5099),
.Y(n_7566)
);

NAND2xp5_ASAP7_75t_L g7567 ( 
.A(n_6621),
.B(n_4842),
.Y(n_7567)
);

NAND2xp5_ASAP7_75t_L g7568 ( 
.A(n_6621),
.B(n_4842),
.Y(n_7568)
);

AND2x4_ASAP7_75t_L g7569 ( 
.A(n_5787),
.B(n_5810),
.Y(n_7569)
);

INVx3_ASAP7_75t_SL g7570 ( 
.A(n_5541),
.Y(n_7570)
);

BUFx12f_ASAP7_75t_L g7571 ( 
.A(n_6038),
.Y(n_7571)
);

NOR2xp33_ASAP7_75t_L g7572 ( 
.A(n_6150),
.B(n_4650),
.Y(n_7572)
);

INVx6_ASAP7_75t_L g7573 ( 
.A(n_5557),
.Y(n_7573)
);

AOI22xp5_ASAP7_75t_L g7574 ( 
.A1(n_5745),
.A2(n_4674),
.B1(n_4691),
.B2(n_4668),
.Y(n_7574)
);

BUFx3_ASAP7_75t_L g7575 ( 
.A(n_6409),
.Y(n_7575)
);

HB1xp67_ASAP7_75t_L g7576 ( 
.A(n_6348),
.Y(n_7576)
);

AOI22xp33_ASAP7_75t_L g7577 ( 
.A1(n_5549),
.A2(n_5260),
.B1(n_5265),
.B2(n_5238),
.Y(n_7577)
);

NOR3xp33_ASAP7_75t_L g7578 ( 
.A(n_5532),
.B(n_4967),
.C(n_4933),
.Y(n_7578)
);

NAND2xp5_ASAP7_75t_SL g7579 ( 
.A(n_6047),
.B(n_5171),
.Y(n_7579)
);

AOI21xp5_ASAP7_75t_L g7580 ( 
.A1(n_6118),
.A2(n_4684),
.B(n_4679),
.Y(n_7580)
);

INVx2_ASAP7_75t_SL g7581 ( 
.A(n_5787),
.Y(n_7581)
);

INVxp67_ASAP7_75t_L g7582 ( 
.A(n_6150),
.Y(n_7582)
);

BUFx3_ASAP7_75t_L g7583 ( 
.A(n_6490),
.Y(n_7583)
);

AOI21xp5_ASAP7_75t_L g7584 ( 
.A1(n_6118),
.A2(n_4684),
.B(n_4679),
.Y(n_7584)
);

OAI22xp5_ASAP7_75t_L g7585 ( 
.A1(n_6500),
.A2(n_5116),
.B1(n_5119),
.B2(n_5115),
.Y(n_7585)
);

BUFx6f_ASAP7_75t_L g7586 ( 
.A(n_6268),
.Y(n_7586)
);

INVx2_ASAP7_75t_SL g7587 ( 
.A(n_5787),
.Y(n_7587)
);

INVx1_ASAP7_75t_SL g7588 ( 
.A(n_5952),
.Y(n_7588)
);

NOR2xp33_ASAP7_75t_L g7589 ( 
.A(n_6159),
.B(n_4722),
.Y(n_7589)
);

BUFx3_ASAP7_75t_L g7590 ( 
.A(n_6490),
.Y(n_7590)
);

INVx2_ASAP7_75t_SL g7591 ( 
.A(n_5810),
.Y(n_7591)
);

AOI222xp33_ASAP7_75t_L g7592 ( 
.A1(n_5634),
.A2(n_5219),
.B1(n_5202),
.B2(n_5223),
.C1(n_5216),
.C2(n_5205),
.Y(n_7592)
);

CKINVDCx5p33_ASAP7_75t_R g7593 ( 
.A(n_5965),
.Y(n_7593)
);

NAND3xp33_ASAP7_75t_L g7594 ( 
.A(n_6224),
.B(n_5219),
.C(n_5216),
.Y(n_7594)
);

O2A1O1Ixp33_ASAP7_75t_L g7595 ( 
.A1(n_5569),
.A2(n_5365),
.B(n_5251),
.C(n_5333),
.Y(n_7595)
);

INVx1_ASAP7_75t_SL g7596 ( 
.A(n_5952),
.Y(n_7596)
);

O2A1O1Ixp5_ASAP7_75t_L g7597 ( 
.A1(n_5752),
.A2(n_5287),
.B(n_5363),
.C(n_5197),
.Y(n_7597)
);

NAND2xp5_ASAP7_75t_SL g7598 ( 
.A(n_6052),
.B(n_5171),
.Y(n_7598)
);

AOI22xp5_ASAP7_75t_L g7599 ( 
.A1(n_5745),
.A2(n_4691),
.B1(n_4702),
.B2(n_4674),
.Y(n_7599)
);

OAI22xp5_ASAP7_75t_L g7600 ( 
.A1(n_6115),
.A2(n_5119),
.B1(n_5127),
.B2(n_5116),
.Y(n_7600)
);

BUFx12f_ASAP7_75t_L g7601 ( 
.A(n_6038),
.Y(n_7601)
);

AOI21xp5_ASAP7_75t_L g7602 ( 
.A1(n_6131),
.A2(n_4686),
.B(n_4684),
.Y(n_7602)
);

BUFx5_ASAP7_75t_L g7603 ( 
.A(n_5547),
.Y(n_7603)
);

OAI22xp5_ASAP7_75t_L g7604 ( 
.A1(n_5828),
.A2(n_5119),
.B1(n_5127),
.B2(n_5116),
.Y(n_7604)
);

BUFx10_ASAP7_75t_L g7605 ( 
.A(n_5891),
.Y(n_7605)
);

INVxp67_ASAP7_75t_L g7606 ( 
.A(n_6159),
.Y(n_7606)
);

NAND3xp33_ASAP7_75t_L g7607 ( 
.A(n_5939),
.B(n_5223),
.C(n_4693),
.Y(n_7607)
);

INVx1_ASAP7_75t_SL g7608 ( 
.A(n_5952),
.Y(n_7608)
);

OAI22xp33_ASAP7_75t_L g7609 ( 
.A1(n_5814),
.A2(n_5268),
.B1(n_5314),
.B2(n_5230),
.Y(n_7609)
);

OR2x2_ASAP7_75t_L g7610 ( 
.A(n_5652),
.B(n_5658),
.Y(n_7610)
);

INVxp67_ASAP7_75t_L g7611 ( 
.A(n_6590),
.Y(n_7611)
);

BUFx3_ASAP7_75t_L g7612 ( 
.A(n_6491),
.Y(n_7612)
);

NOR2xp33_ASAP7_75t_L g7613 ( 
.A(n_6227),
.B(n_4722),
.Y(n_7613)
);

AOI22xp5_ASAP7_75t_L g7614 ( 
.A1(n_5755),
.A2(n_4691),
.B1(n_4702),
.B2(n_4674),
.Y(n_7614)
);

BUFx12f_ASAP7_75t_L g7615 ( 
.A(n_6109),
.Y(n_7615)
);

OAI22xp5_ASAP7_75t_SL g7616 ( 
.A1(n_6345),
.A2(n_4825),
.B1(n_4844),
.B2(n_4819),
.Y(n_7616)
);

CKINVDCx5p33_ASAP7_75t_R g7617 ( 
.A(n_5973),
.Y(n_7617)
);

AOI21xp5_ASAP7_75t_L g7618 ( 
.A1(n_6131),
.A2(n_4693),
.B(n_4686),
.Y(n_7618)
);

NOR2xp67_ASAP7_75t_L g7619 ( 
.A(n_5829),
.B(n_4852),
.Y(n_7619)
);

BUFx2_ASAP7_75t_SL g7620 ( 
.A(n_6491),
.Y(n_7620)
);

AOI221xp5_ASAP7_75t_L g7621 ( 
.A1(n_6100),
.A2(n_5135),
.B1(n_5142),
.B2(n_5133),
.C(n_5127),
.Y(n_7621)
);

AOI21xp5_ASAP7_75t_L g7622 ( 
.A1(n_6165),
.A2(n_6176),
.B(n_6166),
.Y(n_7622)
);

INVxp67_ASAP7_75t_SL g7623 ( 
.A(n_6476),
.Y(n_7623)
);

AOI21xp5_ASAP7_75t_L g7624 ( 
.A1(n_6165),
.A2(n_4693),
.B(n_4686),
.Y(n_7624)
);

AND3x4_ASAP7_75t_L g7625 ( 
.A(n_5819),
.B(n_4702),
.C(n_4691),
.Y(n_7625)
);

AOI21x1_ASAP7_75t_SL g7626 ( 
.A1(n_5585),
.A2(n_4593),
.B(n_5307),
.Y(n_7626)
);

CKINVDCx5p33_ASAP7_75t_R g7627 ( 
.A(n_5973),
.Y(n_7627)
);

NOR2xp67_ASAP7_75t_SL g7628 ( 
.A(n_5701),
.B(n_5498),
.Y(n_7628)
);

AOI22xp33_ASAP7_75t_L g7629 ( 
.A1(n_5743),
.A2(n_5678),
.B1(n_5676),
.B2(n_5752),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_5911),
.B(n_5916),
.Y(n_7630)
);

CKINVDCx5p33_ASAP7_75t_R g7631 ( 
.A(n_5978),
.Y(n_7631)
);

INVx8_ASAP7_75t_L g7632 ( 
.A(n_5547),
.Y(n_7632)
);

NAND2xp5_ASAP7_75t_SL g7633 ( 
.A(n_6100),
.B(n_5171),
.Y(n_7633)
);

INVx4_ASAP7_75t_L g7634 ( 
.A(n_5586),
.Y(n_7634)
);

NOR2xp33_ASAP7_75t_L g7635 ( 
.A(n_6227),
.B(n_4722),
.Y(n_7635)
);

BUFx2_ASAP7_75t_SL g7636 ( 
.A(n_6491),
.Y(n_7636)
);

NAND2xp5_ASAP7_75t_L g7637 ( 
.A(n_6455),
.B(n_6466),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_SL g7638 ( 
.A(n_5659),
.B(n_6427),
.Y(n_7638)
);

NOR2xp33_ASAP7_75t_L g7639 ( 
.A(n_6253),
.B(n_6254),
.Y(n_7639)
);

O2A1O1Ixp33_ASAP7_75t_L g7640 ( 
.A1(n_5569),
.A2(n_5251),
.B(n_5333),
.C(n_5203),
.Y(n_7640)
);

CKINVDCx5p33_ASAP7_75t_R g7641 ( 
.A(n_5978),
.Y(n_7641)
);

AOI21xp5_ASAP7_75t_L g7642 ( 
.A1(n_6166),
.A2(n_4693),
.B(n_4686),
.Y(n_7642)
);

AOI222xp33_ASAP7_75t_L g7643 ( 
.A1(n_5678),
.A2(n_5211),
.B1(n_5212),
.B2(n_5173),
.C1(n_5135),
.C2(n_5133),
.Y(n_7643)
);

BUFx3_ASAP7_75t_L g7644 ( 
.A(n_6526),
.Y(n_7644)
);

CKINVDCx5p33_ASAP7_75t_R g7645 ( 
.A(n_5978),
.Y(n_7645)
);

NAND2xp5_ASAP7_75t_SL g7646 ( 
.A(n_5659),
.B(n_5171),
.Y(n_7646)
);

BUFx3_ASAP7_75t_L g7647 ( 
.A(n_6526),
.Y(n_7647)
);

AOI21xp5_ASAP7_75t_L g7648 ( 
.A1(n_6176),
.A2(n_4693),
.B(n_4686),
.Y(n_7648)
);

AOI22xp33_ASAP7_75t_L g7649 ( 
.A1(n_5743),
.A2(n_5260),
.B1(n_5265),
.B2(n_5238),
.Y(n_7649)
);

INVx4_ASAP7_75t_L g7650 ( 
.A(n_5586),
.Y(n_7650)
);

AOI21xp5_ASAP7_75t_L g7651 ( 
.A1(n_6180),
.A2(n_4693),
.B(n_4686),
.Y(n_7651)
);

HB1xp67_ASAP7_75t_L g7652 ( 
.A(n_6374),
.Y(n_7652)
);

INVxp67_ASAP7_75t_SL g7653 ( 
.A(n_6476),
.Y(n_7653)
);

INVx2_ASAP7_75t_SL g7654 ( 
.A(n_5810),
.Y(n_7654)
);

NAND2xp5_ASAP7_75t_SL g7655 ( 
.A(n_6427),
.B(n_5180),
.Y(n_7655)
);

INVxp67_ASAP7_75t_L g7656 ( 
.A(n_6590),
.Y(n_7656)
);

BUFx6f_ASAP7_75t_L g7657 ( 
.A(n_6310),
.Y(n_7657)
);

AOI22xp5_ASAP7_75t_L g7658 ( 
.A1(n_5755),
.A2(n_4828),
.B1(n_4829),
.B2(n_4785),
.Y(n_7658)
);

HB1xp67_ASAP7_75t_L g7659 ( 
.A(n_6374),
.Y(n_7659)
);

AOI22xp33_ASAP7_75t_L g7660 ( 
.A1(n_5676),
.A2(n_5260),
.B1(n_5265),
.B2(n_5238),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_6253),
.B(n_4722),
.Y(n_7661)
);

CKINVDCx5p33_ASAP7_75t_R g7662 ( 
.A(n_6008),
.Y(n_7662)
);

NOR2xp33_ASAP7_75t_L g7663 ( 
.A(n_6254),
.B(n_4722),
.Y(n_7663)
);

NAND2xp33_ASAP7_75t_L g7664 ( 
.A(n_6570),
.B(n_4865),
.Y(n_7664)
);

OAI22xp5_ASAP7_75t_L g7665 ( 
.A1(n_5828),
.A2(n_5804),
.B1(n_5786),
.B2(n_5814),
.Y(n_7665)
);

NAND2xp5_ASAP7_75t_L g7666 ( 
.A(n_6455),
.B(n_4859),
.Y(n_7666)
);

AOI21xp5_ASAP7_75t_L g7667 ( 
.A1(n_6180),
.A2(n_6203),
.B(n_6199),
.Y(n_7667)
);

BUFx2_ASAP7_75t_SL g7668 ( 
.A(n_6526),
.Y(n_7668)
);

BUFx6f_ASAP7_75t_SL g7669 ( 
.A(n_6157),
.Y(n_7669)
);

AOI21xp5_ASAP7_75t_L g7670 ( 
.A1(n_6199),
.A2(n_4741),
.B(n_4693),
.Y(n_7670)
);

INVx2_ASAP7_75t_SL g7671 ( 
.A(n_5812),
.Y(n_7671)
);

CKINVDCx16_ASAP7_75t_R g7672 ( 
.A(n_6345),
.Y(n_7672)
);

INVx1_ASAP7_75t_SL g7673 ( 
.A(n_5962),
.Y(n_7673)
);

NOR2xp33_ASAP7_75t_SL g7674 ( 
.A(n_6543),
.B(n_4474),
.Y(n_7674)
);

CKINVDCx20_ASAP7_75t_R g7675 ( 
.A(n_6358),
.Y(n_7675)
);

AOI21xp5_ASAP7_75t_L g7676 ( 
.A1(n_6203),
.A2(n_4741),
.B(n_4693),
.Y(n_7676)
);

O2A1O1Ixp33_ASAP7_75t_L g7677 ( 
.A1(n_5599),
.A2(n_5333),
.B(n_5350),
.C(n_5203),
.Y(n_7677)
);

CKINVDCx20_ASAP7_75t_R g7678 ( 
.A(n_6538),
.Y(n_7678)
);

CKINVDCx5p33_ASAP7_75t_R g7679 ( 
.A(n_6008),
.Y(n_7679)
);

AND2x4_ASAP7_75t_L g7680 ( 
.A(n_5812),
.B(n_5850),
.Y(n_7680)
);

NAND2x1p5_ASAP7_75t_L g7681 ( 
.A(n_5829),
.B(n_4474),
.Y(n_7681)
);

HB1xp67_ASAP7_75t_L g7682 ( 
.A(n_6505),
.Y(n_7682)
);

OAI221xp5_ASAP7_75t_L g7683 ( 
.A1(n_5602),
.A2(n_5492),
.B1(n_5475),
.B2(n_5474),
.C(n_5386),
.Y(n_7683)
);

CKINVDCx20_ASAP7_75t_R g7684 ( 
.A(n_6540),
.Y(n_7684)
);

BUFx2_ASAP7_75t_SL g7685 ( 
.A(n_6543),
.Y(n_7685)
);

INVxp67_ASAP7_75t_SL g7686 ( 
.A(n_6496),
.Y(n_7686)
);

NAND2xp5_ASAP7_75t_L g7687 ( 
.A(n_6466),
.B(n_4859),
.Y(n_7687)
);

AOI21xp5_ASAP7_75t_L g7688 ( 
.A1(n_6225),
.A2(n_6250),
.B(n_6238),
.Y(n_7688)
);

NAND2xp5_ASAP7_75t_L g7689 ( 
.A(n_6478),
.B(n_4859),
.Y(n_7689)
);

CKINVDCx20_ASAP7_75t_R g7690 ( 
.A(n_6542),
.Y(n_7690)
);

AOI22xp5_ASAP7_75t_L g7691 ( 
.A1(n_5757),
.A2(n_4828),
.B1(n_4829),
.B2(n_4785),
.Y(n_7691)
);

AOI21x1_ASAP7_75t_L g7692 ( 
.A1(n_6486),
.A2(n_5492),
.B(n_5475),
.Y(n_7692)
);

CKINVDCx5p33_ASAP7_75t_R g7693 ( 
.A(n_6008),
.Y(n_7693)
);

AOI22xp33_ASAP7_75t_L g7694 ( 
.A1(n_5736),
.A2(n_5271),
.B1(n_5265),
.B2(n_4825),
.Y(n_7694)
);

NAND2x1p5_ASAP7_75t_L g7695 ( 
.A(n_5829),
.B(n_4474),
.Y(n_7695)
);

HB1xp67_ASAP7_75t_L g7696 ( 
.A(n_6505),
.Y(n_7696)
);

AOI222xp33_ASAP7_75t_L g7697 ( 
.A1(n_5759),
.A2(n_5826),
.B1(n_5765),
.B2(n_5882),
.C1(n_6510),
.C2(n_5741),
.Y(n_7697)
);

NAND2xp5_ASAP7_75t_L g7698 ( 
.A(n_6478),
.B(n_4859),
.Y(n_7698)
);

AOI22xp33_ASAP7_75t_L g7699 ( 
.A1(n_5736),
.A2(n_5271),
.B1(n_4825),
.B2(n_4844),
.Y(n_7699)
);

NOR2xp33_ASAP7_75t_L g7700 ( 
.A(n_6266),
.B(n_4722),
.Y(n_7700)
);

BUFx4f_ASAP7_75t_SL g7701 ( 
.A(n_6109),
.Y(n_7701)
);

AOI21xp5_ASAP7_75t_L g7702 ( 
.A1(n_6225),
.A2(n_4747),
.B(n_4741),
.Y(n_7702)
);

OAI21x1_ASAP7_75t_L g7703 ( 
.A1(n_6238),
.A2(n_4875),
.B(n_4862),
.Y(n_7703)
);

OAI22xp33_ASAP7_75t_L g7704 ( 
.A1(n_6457),
.A2(n_5268),
.B1(n_5314),
.B2(n_5230),
.Y(n_7704)
);

AOI21xp5_ASAP7_75t_L g7705 ( 
.A1(n_6680),
.A2(n_6754),
.B(n_6881),
.Y(n_7705)
);

OAI21x1_ASAP7_75t_L g7706 ( 
.A1(n_6943),
.A2(n_6341),
.B(n_6250),
.Y(n_7706)
);

AO31x2_ASAP7_75t_L g7707 ( 
.A1(n_6754),
.A2(n_5832),
.A3(n_6229),
.B(n_5785),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_6723),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_6723),
.Y(n_7709)
);

AOI222xp33_ASAP7_75t_L g7710 ( 
.A1(n_6690),
.A2(n_5882),
.B1(n_5759),
.B2(n_5826),
.C1(n_5765),
.C2(n_5537),
.Y(n_7710)
);

BUFx6f_ASAP7_75t_L g7711 ( 
.A(n_7329),
.Y(n_7711)
);

OR2x6_ASAP7_75t_L g7712 ( 
.A(n_7632),
.B(n_6410),
.Y(n_7712)
);

OAI21xp5_ASAP7_75t_L g7713 ( 
.A1(n_7071),
.A2(n_6501),
.B(n_6128),
.Y(n_7713)
);

OAI22xp5_ASAP7_75t_L g7714 ( 
.A1(n_6690),
.A2(n_6457),
.B1(n_5773),
.B2(n_5804),
.Y(n_7714)
);

OA21x2_ASAP7_75t_L g7715 ( 
.A1(n_7276),
.A2(n_6608),
.B(n_6592),
.Y(n_7715)
);

INVx1_ASAP7_75t_L g7716 ( 
.A(n_6723),
.Y(n_7716)
);

OR2x2_ASAP7_75t_L g7717 ( 
.A(n_6713),
.B(n_6420),
.Y(n_7717)
);

OAI21x1_ASAP7_75t_L g7718 ( 
.A1(n_6943),
.A2(n_7276),
.B(n_6869),
.Y(n_7718)
);

BUFx3_ASAP7_75t_L g7719 ( 
.A(n_6751),
.Y(n_7719)
);

INVx2_ASAP7_75t_L g7720 ( 
.A(n_6721),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_6724),
.Y(n_7721)
);

AO31x2_ASAP7_75t_L g7722 ( 
.A1(n_6870),
.A2(n_5832),
.A3(n_6229),
.B(n_5785),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_6724),
.Y(n_7723)
);

OAI21x1_ASAP7_75t_L g7724 ( 
.A1(n_6943),
.A2(n_6352),
.B(n_6341),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_6724),
.Y(n_7725)
);

OAI21x1_ASAP7_75t_L g7726 ( 
.A1(n_6943),
.A2(n_6368),
.B(n_6352),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_6731),
.Y(n_7727)
);

AOI22xp33_ASAP7_75t_L g7728 ( 
.A1(n_6983),
.A2(n_5819),
.B1(n_6367),
.B2(n_6434),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_6731),
.Y(n_7729)
);

CKINVDCx20_ASAP7_75t_R g7730 ( 
.A(n_6973),
.Y(n_7730)
);

AND2x2_ASAP7_75t_L g7731 ( 
.A(n_6713),
.B(n_6027),
.Y(n_7731)
);

AND2x4_ASAP7_75t_L g7732 ( 
.A(n_7318),
.B(n_5812),
.Y(n_7732)
);

OAI21x1_ASAP7_75t_L g7733 ( 
.A1(n_7276),
.A2(n_6384),
.B(n_6368),
.Y(n_7733)
);

OAI21x1_ASAP7_75t_L g7734 ( 
.A1(n_7276),
.A2(n_6398),
.B(n_6384),
.Y(n_7734)
);

INVx1_ASAP7_75t_L g7735 ( 
.A(n_6731),
.Y(n_7735)
);

NAND2xp5_ASAP7_75t_L g7736 ( 
.A(n_6786),
.B(n_6547),
.Y(n_7736)
);

INVx2_ASAP7_75t_L g7737 ( 
.A(n_6721),
.Y(n_7737)
);

AOI21xp33_ASAP7_75t_L g7738 ( 
.A1(n_6763),
.A2(n_6128),
.B(n_6113),
.Y(n_7738)
);

OAI21x1_ASAP7_75t_L g7739 ( 
.A1(n_6738),
.A2(n_6412),
.B(n_6398),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6735),
.Y(n_7740)
);

OA21x2_ASAP7_75t_L g7741 ( 
.A1(n_7343),
.A2(n_6608),
.B(n_6503),
.Y(n_7741)
);

NAND2xp5_ASAP7_75t_SL g7742 ( 
.A(n_7071),
.B(n_7427),
.Y(n_7742)
);

OAI21x1_ASAP7_75t_L g7743 ( 
.A1(n_6738),
.A2(n_6422),
.B(n_6412),
.Y(n_7743)
);

AOI21xp5_ASAP7_75t_L g7744 ( 
.A1(n_6680),
.A2(n_6422),
.B(n_5611),
.Y(n_7744)
);

INVx2_ASAP7_75t_L g7745 ( 
.A(n_6721),
.Y(n_7745)
);

OAI21xp5_ASAP7_75t_SL g7746 ( 
.A1(n_7291),
.A2(n_6506),
.B(n_5537),
.Y(n_7746)
);

OA21x2_ASAP7_75t_L g7747 ( 
.A1(n_7343),
.A2(n_7411),
.B(n_7380),
.Y(n_7747)
);

A2O1A1Ixp33_ASAP7_75t_L g7748 ( 
.A1(n_6763),
.A2(n_5534),
.B(n_5786),
.C(n_6059),
.Y(n_7748)
);

AND2x4_ASAP7_75t_L g7749 ( 
.A(n_7318),
.B(n_5812),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_6735),
.Y(n_7750)
);

OA21x2_ASAP7_75t_L g7751 ( 
.A1(n_7380),
.A2(n_6503),
.B(n_6501),
.Y(n_7751)
);

AND2x2_ASAP7_75t_L g7752 ( 
.A(n_6713),
.B(n_6027),
.Y(n_7752)
);

OAI21x1_ASAP7_75t_L g7753 ( 
.A1(n_6869),
.A2(n_6541),
.B(n_6589),
.Y(n_7753)
);

NOR2xp33_ASAP7_75t_L g7754 ( 
.A(n_6710),
.B(n_6168),
.Y(n_7754)
);

AO21x2_ASAP7_75t_L g7755 ( 
.A1(n_6881),
.A2(n_6110),
.B(n_6079),
.Y(n_7755)
);

AOI21xp5_ASAP7_75t_SL g7756 ( 
.A1(n_7450),
.A2(n_6113),
.B(n_6175),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_6735),
.Y(n_7757)
);

HB1xp67_ASAP7_75t_L g7758 ( 
.A(n_6798),
.Y(n_7758)
);

OA21x2_ASAP7_75t_L g7759 ( 
.A1(n_7411),
.A2(n_6059),
.B(n_6298),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_6769),
.Y(n_7760)
);

AO21x2_ASAP7_75t_L g7761 ( 
.A1(n_6821),
.A2(n_6110),
.B(n_6079),
.Y(n_7761)
);

INVxp67_ASAP7_75t_SL g7762 ( 
.A(n_6870),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_6769),
.Y(n_7763)
);

OAI22xp5_ASAP7_75t_L g7764 ( 
.A1(n_7291),
.A2(n_5773),
.B1(n_6226),
.B2(n_6151),
.Y(n_7764)
);

AND2x2_ASAP7_75t_L g7765 ( 
.A(n_6730),
.B(n_6027),
.Y(n_7765)
);

NAND2x1p5_ASAP7_75t_L g7766 ( 
.A(n_7628),
.B(n_5586),
.Y(n_7766)
);

AOI22xp33_ASAP7_75t_SL g7767 ( 
.A1(n_7401),
.A2(n_6000),
.B1(n_6367),
.B2(n_5919),
.Y(n_7767)
);

INVx3_ASAP7_75t_L g7768 ( 
.A(n_6631),
.Y(n_7768)
);

AOI22xp5_ASAP7_75t_L g7769 ( 
.A1(n_7291),
.A2(n_5839),
.B1(n_6506),
.B2(n_5791),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_L g7770 ( 
.A(n_6786),
.B(n_6547),
.Y(n_7770)
);

INVx6_ASAP7_75t_L g7771 ( 
.A(n_7318),
.Y(n_7771)
);

OR2x2_ASAP7_75t_L g7772 ( 
.A(n_6730),
.B(n_6420),
.Y(n_7772)
);

NAND2xp33_ASAP7_75t_SL g7773 ( 
.A(n_6979),
.B(n_5649),
.Y(n_7773)
);

NOR2x1_ASAP7_75t_SL g7774 ( 
.A(n_7382),
.B(n_5747),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_6786),
.B(n_6417),
.Y(n_7775)
);

O2A1O1Ixp33_ASAP7_75t_SL g7776 ( 
.A1(n_6683),
.A2(n_5692),
.B(n_5846),
.C(n_5646),
.Y(n_7776)
);

INVx2_ASAP7_75t_L g7777 ( 
.A(n_6721),
.Y(n_7777)
);

AO21x2_ASAP7_75t_L g7778 ( 
.A1(n_6821),
.A2(n_6110),
.B(n_6079),
.Y(n_7778)
);

OAI21x1_ASAP7_75t_L g7779 ( 
.A1(n_7255),
.A2(n_6589),
.B(n_6578),
.Y(n_7779)
);

OAI21x1_ASAP7_75t_L g7780 ( 
.A1(n_7255),
.A2(n_6578),
.B(n_6533),
.Y(n_7780)
);

OAI21x1_ASAP7_75t_L g7781 ( 
.A1(n_7310),
.A2(n_6578),
.B(n_6533),
.Y(n_7781)
);

AOI21xp5_ASAP7_75t_L g7782 ( 
.A1(n_6770),
.A2(n_5611),
.B(n_6242),
.Y(n_7782)
);

AOI22xp33_ASAP7_75t_L g7783 ( 
.A1(n_6983),
.A2(n_6434),
.B1(n_5602),
.B2(n_5613),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_6769),
.Y(n_7784)
);

AO21x2_ASAP7_75t_L g7785 ( 
.A1(n_6770),
.A2(n_6522),
.B(n_6416),
.Y(n_7785)
);

AO32x2_ASAP7_75t_L g7786 ( 
.A1(n_7382),
.A2(n_6205),
.A3(n_6620),
.B1(n_6617),
.B2(n_5909),
.Y(n_7786)
);

HB1xp67_ASAP7_75t_L g7787 ( 
.A(n_6798),
.Y(n_7787)
);

AND3x2_ASAP7_75t_L g7788 ( 
.A(n_7427),
.B(n_7240),
.C(n_7171),
.Y(n_7788)
);

INVx2_ASAP7_75t_L g7789 ( 
.A(n_6734),
.Y(n_7789)
);

AOI22xp33_ASAP7_75t_L g7790 ( 
.A1(n_7462),
.A2(n_5613),
.B1(n_5757),
.B2(n_5758),
.Y(n_7790)
);

O2A1O1Ixp33_ASAP7_75t_SL g7791 ( 
.A1(n_6683),
.A2(n_5846),
.B(n_5646),
.C(n_5703),
.Y(n_7791)
);

AND2x4_ASAP7_75t_L g7792 ( 
.A(n_7318),
.B(n_5812),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_6775),
.Y(n_7793)
);

CKINVDCx5p33_ASAP7_75t_R g7794 ( 
.A(n_6855),
.Y(n_7794)
);

AO21x1_ASAP7_75t_L g7795 ( 
.A1(n_7171),
.A2(n_5534),
.B(n_6175),
.Y(n_7795)
);

OA21x2_ASAP7_75t_L g7796 ( 
.A1(n_7435),
.A2(n_6298),
.B(n_6090),
.Y(n_7796)
);

OAI22xp5_ASAP7_75t_L g7797 ( 
.A1(n_7629),
.A2(n_6226),
.B1(n_6151),
.B2(n_6183),
.Y(n_7797)
);

AOI22xp33_ASAP7_75t_L g7798 ( 
.A1(n_7462),
.A2(n_5758),
.B1(n_5778),
.B2(n_5654),
.Y(n_7798)
);

NAND4xp25_ASAP7_75t_L g7799 ( 
.A(n_7450),
.B(n_6392),
.C(n_5599),
.D(n_5532),
.Y(n_7799)
);

INVx2_ASAP7_75t_L g7800 ( 
.A(n_6734),
.Y(n_7800)
);

NAND2xp5_ASAP7_75t_L g7801 ( 
.A(n_6787),
.B(n_6417),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_6775),
.Y(n_7802)
);

OAI21xp5_ASAP7_75t_L g7803 ( 
.A1(n_7427),
.A2(n_6090),
.B(n_5582),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_6775),
.Y(n_7804)
);

OAI21x1_ASAP7_75t_L g7805 ( 
.A1(n_7445),
.A2(n_5555),
.B(n_6602),
.Y(n_7805)
);

OAI21xp5_ASAP7_75t_L g7806 ( 
.A1(n_7401),
.A2(n_5582),
.B(n_5654),
.Y(n_7806)
);

NOR3xp33_ASAP7_75t_SL g7807 ( 
.A(n_6622),
.B(n_6614),
.C(n_5741),
.Y(n_7807)
);

AO21x2_ASAP7_75t_L g7808 ( 
.A1(n_6771),
.A2(n_6522),
.B(n_6416),
.Y(n_7808)
);

INVx2_ASAP7_75t_L g7809 ( 
.A(n_6734),
.Y(n_7809)
);

AO21x2_ASAP7_75t_L g7810 ( 
.A1(n_6771),
.A2(n_6423),
.B(n_5621),
.Y(n_7810)
);

HB1xp67_ASAP7_75t_L g7811 ( 
.A(n_6803),
.Y(n_7811)
);

OAI21x1_ASAP7_75t_L g7812 ( 
.A1(n_7445),
.A2(n_5555),
.B(n_6602),
.Y(n_7812)
);

OAI21x1_ASAP7_75t_L g7813 ( 
.A1(n_7459),
.A2(n_6602),
.B(n_6004),
.Y(n_7813)
);

NOR2xp33_ASAP7_75t_L g7814 ( 
.A(n_6710),
.B(n_6168),
.Y(n_7814)
);

OA21x2_ASAP7_75t_L g7815 ( 
.A1(n_7459),
.A2(n_6324),
.B(n_6423),
.Y(n_7815)
);

OAI21x1_ASAP7_75t_L g7816 ( 
.A1(n_7487),
.A2(n_6004),
.B(n_6156),
.Y(n_7816)
);

CKINVDCx9p33_ASAP7_75t_R g7817 ( 
.A(n_6740),
.Y(n_7817)
);

OAI21x1_ASAP7_75t_L g7818 ( 
.A1(n_7487),
.A2(n_6004),
.B(n_6156),
.Y(n_7818)
);

OAI21x1_ASAP7_75t_L g7819 ( 
.A1(n_7495),
.A2(n_6297),
.B(n_6156),
.Y(n_7819)
);

AOI21xp5_ASAP7_75t_L g7820 ( 
.A1(n_6707),
.A2(n_6242),
.B(n_6267),
.Y(n_7820)
);

INVx3_ASAP7_75t_SL g7821 ( 
.A(n_6835),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_6789),
.Y(n_7822)
);

AND2x4_ASAP7_75t_L g7823 ( 
.A(n_7318),
.B(n_5812),
.Y(n_7823)
);

AOI21x1_ASAP7_75t_L g7824 ( 
.A1(n_7638),
.A2(n_6229),
.B(n_5672),
.Y(n_7824)
);

CKINVDCx20_ASAP7_75t_R g7825 ( 
.A(n_6973),
.Y(n_7825)
);

AND2x2_ASAP7_75t_L g7826 ( 
.A(n_6730),
.B(n_6069),
.Y(n_7826)
);

AND2x2_ASAP7_75t_L g7827 ( 
.A(n_6747),
.B(n_6069),
.Y(n_7827)
);

AO21x2_ASAP7_75t_L g7828 ( 
.A1(n_6994),
.A2(n_5621),
.B(n_5766),
.Y(n_7828)
);

BUFx2_ASAP7_75t_L g7829 ( 
.A(n_7420),
.Y(n_7829)
);

AND2x2_ASAP7_75t_L g7830 ( 
.A(n_6747),
.B(n_6069),
.Y(n_7830)
);

INVx2_ASAP7_75t_L g7831 ( 
.A(n_6734),
.Y(n_7831)
);

OA21x2_ASAP7_75t_L g7832 ( 
.A1(n_7495),
.A2(n_7541),
.B(n_7506),
.Y(n_7832)
);

AOI22xp33_ASAP7_75t_L g7833 ( 
.A1(n_6968),
.A2(n_5778),
.B1(n_5749),
.B2(n_5839),
.Y(n_7833)
);

OAI21x1_ASAP7_75t_L g7834 ( 
.A1(n_7506),
.A2(n_6297),
.B(n_5672),
.Y(n_7834)
);

OAI21x1_ASAP7_75t_L g7835 ( 
.A1(n_7541),
.A2(n_6297),
.B(n_5668),
.Y(n_7835)
);

OAI21x1_ASAP7_75t_L g7836 ( 
.A1(n_7558),
.A2(n_5668),
.B(n_5940),
.Y(n_7836)
);

NAND2xp5_ASAP7_75t_SL g7837 ( 
.A(n_7101),
.B(n_5609),
.Y(n_7837)
);

NAND2xp5_ASAP7_75t_L g7838 ( 
.A(n_6787),
.B(n_5740),
.Y(n_7838)
);

INVx2_ASAP7_75t_L g7839 ( 
.A(n_6742),
.Y(n_7839)
);

NOR2xp33_ASAP7_75t_L g7840 ( 
.A(n_7412),
.B(n_6189),
.Y(n_7840)
);

OA21x2_ASAP7_75t_L g7841 ( 
.A1(n_7558),
.A2(n_7584),
.B(n_7580),
.Y(n_7841)
);

OAI21x1_ASAP7_75t_L g7842 ( 
.A1(n_7580),
.A2(n_5940),
.B(n_5693),
.Y(n_7842)
);

AO21x2_ASAP7_75t_L g7843 ( 
.A1(n_6994),
.A2(n_5766),
.B(n_5581),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_6968),
.A2(n_7401),
.B1(n_7488),
.B2(n_7531),
.Y(n_7844)
);

NAND2x1_ASAP7_75t_L g7845 ( 
.A(n_6751),
.B(n_5812),
.Y(n_7845)
);

INVx1_ASAP7_75t_L g7846 ( 
.A(n_6789),
.Y(n_7846)
);

OAI21x1_ASAP7_75t_L g7847 ( 
.A1(n_7584),
.A2(n_5940),
.B(n_5693),
.Y(n_7847)
);

AND2x2_ASAP7_75t_L g7848 ( 
.A(n_6747),
.B(n_6792),
.Y(n_7848)
);

OAI22xp5_ASAP7_75t_SL g7849 ( 
.A1(n_7101),
.A2(n_6539),
.B1(n_5627),
.B2(n_5789),
.Y(n_7849)
);

INVx4_ASAP7_75t_L g7850 ( 
.A(n_6750),
.Y(n_7850)
);

INVxp67_ASAP7_75t_SL g7851 ( 
.A(n_6870),
.Y(n_7851)
);

OAI21x1_ASAP7_75t_L g7852 ( 
.A1(n_7602),
.A2(n_5751),
.B(n_5615),
.Y(n_7852)
);

INVx2_ASAP7_75t_L g7853 ( 
.A(n_6742),
.Y(n_7853)
);

CKINVDCx20_ASAP7_75t_R g7854 ( 
.A(n_6995),
.Y(n_7854)
);

OAI21xp5_ASAP7_75t_L g7855 ( 
.A1(n_7531),
.A2(n_5567),
.B(n_5854),
.Y(n_7855)
);

AND2x2_ASAP7_75t_L g7856 ( 
.A(n_6792),
.B(n_5675),
.Y(n_7856)
);

INVx2_ASAP7_75t_L g7857 ( 
.A(n_6742),
.Y(n_7857)
);

OAI21x1_ASAP7_75t_L g7858 ( 
.A1(n_7602),
.A2(n_5751),
.B(n_5615),
.Y(n_7858)
);

AND2x2_ASAP7_75t_L g7859 ( 
.A(n_6792),
.B(n_5675),
.Y(n_7859)
);

OAI21x1_ASAP7_75t_L g7860 ( 
.A1(n_7618),
.A2(n_5615),
.B(n_6418),
.Y(n_7860)
);

AO21x2_ASAP7_75t_L g7861 ( 
.A1(n_7013),
.A2(n_5766),
.B(n_6324),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_6789),
.Y(n_7862)
);

CKINVDCx5p33_ASAP7_75t_R g7863 ( 
.A(n_6855),
.Y(n_7863)
);

AND2x2_ASAP7_75t_L g7864 ( 
.A(n_6797),
.B(n_6580),
.Y(n_7864)
);

AOI211xp5_ASAP7_75t_L g7865 ( 
.A1(n_7531),
.A2(n_5872),
.B(n_5849),
.C(n_5792),
.Y(n_7865)
);

AOI21xp5_ASAP7_75t_L g7866 ( 
.A1(n_6707),
.A2(n_6242),
.B(n_6267),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_6802),
.Y(n_7867)
);

OAI21x1_ASAP7_75t_L g7868 ( 
.A1(n_7618),
.A2(n_5615),
.B(n_6418),
.Y(n_7868)
);

OAI21x1_ASAP7_75t_L g7869 ( 
.A1(n_7624),
.A2(n_5615),
.B(n_6418),
.Y(n_7869)
);

BUFx6f_ASAP7_75t_L g7870 ( 
.A(n_7329),
.Y(n_7870)
);

INVxp33_ASAP7_75t_L g7871 ( 
.A(n_6815),
.Y(n_7871)
);

OR2x2_ASAP7_75t_L g7872 ( 
.A(n_6797),
.B(n_6420),
.Y(n_7872)
);

OAI21x1_ASAP7_75t_L g7873 ( 
.A1(n_7642),
.A2(n_7651),
.B(n_7648),
.Y(n_7873)
);

AO31x2_ASAP7_75t_L g7874 ( 
.A1(n_7033),
.A2(n_7387),
.A3(n_7600),
.B(n_7377),
.Y(n_7874)
);

OAI21xp5_ASAP7_75t_L g7875 ( 
.A1(n_7178),
.A2(n_5854),
.B(n_5682),
.Y(n_7875)
);

CKINVDCx20_ASAP7_75t_R g7876 ( 
.A(n_6995),
.Y(n_7876)
);

OR2x6_ASAP7_75t_L g7877 ( 
.A(n_7632),
.B(n_6410),
.Y(n_7877)
);

OAI21x1_ASAP7_75t_L g7878 ( 
.A1(n_7642),
.A2(n_6581),
.B(n_5607),
.Y(n_7878)
);

INVx1_ASAP7_75t_L g7879 ( 
.A(n_6802),
.Y(n_7879)
);

AND2x2_ASAP7_75t_L g7880 ( 
.A(n_6797),
.B(n_6580),
.Y(n_7880)
);

BUFx3_ASAP7_75t_L g7881 ( 
.A(n_6751),
.Y(n_7881)
);

BUFx2_ASAP7_75t_L g7882 ( 
.A(n_7420),
.Y(n_7882)
);

HB1xp67_ASAP7_75t_L g7883 ( 
.A(n_6803),
.Y(n_7883)
);

INVx1_ASAP7_75t_L g7884 ( 
.A(n_6802),
.Y(n_7884)
);

OAI21x1_ASAP7_75t_L g7885 ( 
.A1(n_7648),
.A2(n_6581),
.B(n_5607),
.Y(n_7885)
);

AOI22xp33_ASAP7_75t_L g7886 ( 
.A1(n_7488),
.A2(n_6739),
.B1(n_7412),
.B2(n_7629),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_6810),
.Y(n_7887)
);

BUFx12f_ASAP7_75t_L g7888 ( 
.A(n_6999),
.Y(n_7888)
);

A2O1A1Ixp33_ASAP7_75t_L g7889 ( 
.A1(n_6739),
.A2(n_5782),
.B(n_6450),
.C(n_5622),
.Y(n_7889)
);

OAI22xp5_ASAP7_75t_L g7890 ( 
.A1(n_7418),
.A2(n_6182),
.B1(n_6183),
.B2(n_6149),
.Y(n_7890)
);

INVx1_ASAP7_75t_L g7891 ( 
.A(n_6810),
.Y(n_7891)
);

AO21x2_ASAP7_75t_L g7892 ( 
.A1(n_7013),
.A2(n_5766),
.B(n_5756),
.Y(n_7892)
);

HB1xp67_ASAP7_75t_L g7893 ( 
.A(n_6890),
.Y(n_7893)
);

OAI21x1_ASAP7_75t_L g7894 ( 
.A1(n_7651),
.A2(n_6581),
.B(n_5607),
.Y(n_7894)
);

OAI21x1_ASAP7_75t_L g7895 ( 
.A1(n_7670),
.A2(n_6581),
.B(n_5607),
.Y(n_7895)
);

OAI21xp33_ASAP7_75t_L g7896 ( 
.A1(n_7102),
.A2(n_6450),
.B(n_6149),
.Y(n_7896)
);

INVx1_ASAP7_75t_L g7897 ( 
.A(n_6810),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_6824),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_6824),
.Y(n_7899)
);

NAND2xp5_ASAP7_75t_L g7900 ( 
.A(n_6787),
.B(n_5740),
.Y(n_7900)
);

CKINVDCx20_ASAP7_75t_R g7901 ( 
.A(n_6664),
.Y(n_7901)
);

OAI21x1_ASAP7_75t_L g7902 ( 
.A1(n_7670),
.A2(n_6045),
.B(n_5661),
.Y(n_7902)
);

AND2x4_ASAP7_75t_L g7903 ( 
.A(n_7318),
.B(n_5850),
.Y(n_7903)
);

INVx1_ASAP7_75t_L g7904 ( 
.A(n_6824),
.Y(n_7904)
);

BUFx3_ASAP7_75t_L g7905 ( 
.A(n_6751),
.Y(n_7905)
);

OAI21x1_ASAP7_75t_SL g7906 ( 
.A1(n_6745),
.A2(n_5919),
.B(n_5682),
.Y(n_7906)
);

NOR2xp33_ASAP7_75t_L g7907 ( 
.A(n_6931),
.B(n_6189),
.Y(n_7907)
);

INVx2_ASAP7_75t_SL g7908 ( 
.A(n_6649),
.Y(n_7908)
);

OAI21x1_ASAP7_75t_L g7909 ( 
.A1(n_7676),
.A2(n_6045),
.B(n_5661),
.Y(n_7909)
);

INVx2_ASAP7_75t_L g7910 ( 
.A(n_6742),
.Y(n_7910)
);

AOI22xp5_ASAP7_75t_L g7911 ( 
.A1(n_7488),
.A2(n_5791),
.B1(n_5792),
.B2(n_5609),
.Y(n_7911)
);

O2A1O1Ixp33_ASAP7_75t_SL g7912 ( 
.A1(n_6678),
.A2(n_5703),
.B(n_6618),
.C(n_6573),
.Y(n_7912)
);

INVx1_ASAP7_75t_L g7913 ( 
.A(n_6826),
.Y(n_7913)
);

OAI21x1_ASAP7_75t_L g7914 ( 
.A1(n_7676),
.A2(n_5769),
.B(n_5756),
.Y(n_7914)
);

OAI21x1_ASAP7_75t_L g7915 ( 
.A1(n_7702),
.A2(n_5769),
.B(n_6070),
.Y(n_7915)
);

OAI21x1_ASAP7_75t_L g7916 ( 
.A1(n_7702),
.A2(n_6239),
.B(n_6070),
.Y(n_7916)
);

INVx3_ASAP7_75t_L g7917 ( 
.A(n_6631),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_6826),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_6746),
.Y(n_7919)
);

AND2x2_ASAP7_75t_L g7920 ( 
.A(n_6812),
.B(n_6820),
.Y(n_7920)
);

NAND2x1p5_ASAP7_75t_L g7921 ( 
.A(n_7628),
.B(n_5586),
.Y(n_7921)
);

NAND2xp33_ASAP7_75t_L g7922 ( 
.A(n_7102),
.B(n_6539),
.Y(n_7922)
);

NAND2xp5_ASAP7_75t_L g7923 ( 
.A(n_7639),
.B(n_5781),
.Y(n_7923)
);

INVx1_ASAP7_75t_SL g7924 ( 
.A(n_6650),
.Y(n_7924)
);

OR2x2_ASAP7_75t_L g7925 ( 
.A(n_6812),
.B(n_6429),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_6826),
.Y(n_7926)
);

AOI221xp5_ASAP7_75t_L g7927 ( 
.A1(n_7026),
.A2(n_6318),
.B1(n_6266),
.B2(n_6311),
.C(n_6287),
.Y(n_7927)
);

OAI22xp5_ASAP7_75t_L g7928 ( 
.A1(n_7418),
.A2(n_6182),
.B1(n_5855),
.B2(n_5835),
.Y(n_7928)
);

OR2x2_ASAP7_75t_L g7929 ( 
.A(n_6812),
.B(n_6429),
.Y(n_7929)
);

OAI21xp5_ASAP7_75t_L g7930 ( 
.A1(n_7178),
.A2(n_5538),
.B(n_6515),
.Y(n_7930)
);

OAI21x1_ASAP7_75t_L g7931 ( 
.A1(n_7329),
.A2(n_6347),
.B(n_5748),
.Y(n_7931)
);

OAI22xp5_ASAP7_75t_L g7932 ( 
.A1(n_7418),
.A2(n_5855),
.B1(n_5835),
.B2(n_5877),
.Y(n_7932)
);

AND2x4_ASAP7_75t_L g7933 ( 
.A(n_7318),
.B(n_5850),
.Y(n_7933)
);

NAND2xp5_ASAP7_75t_L g7934 ( 
.A(n_7639),
.B(n_6931),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_6837),
.Y(n_7935)
);

INVx2_ASAP7_75t_L g7936 ( 
.A(n_6746),
.Y(n_7936)
);

NOR2xp33_ASAP7_75t_L g7937 ( 
.A(n_6800),
.B(n_6198),
.Y(n_7937)
);

NAND2xp5_ASAP7_75t_L g7938 ( 
.A(n_7637),
.B(n_5781),
.Y(n_7938)
);

OR2x6_ASAP7_75t_L g7939 ( 
.A(n_7632),
.B(n_7154),
.Y(n_7939)
);

INVx2_ASAP7_75t_L g7940 ( 
.A(n_6746),
.Y(n_7940)
);

BUFx3_ASAP7_75t_L g7941 ( 
.A(n_6751),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_6837),
.Y(n_7942)
);

OAI22xp5_ASAP7_75t_L g7943 ( 
.A1(n_6694),
.A2(n_5877),
.B1(n_5717),
.B2(n_5662),
.Y(n_7943)
);

OAI21x1_ASAP7_75t_L g7944 ( 
.A1(n_7325),
.A2(n_6347),
.B(n_5782),
.Y(n_7944)
);

INVx1_ASAP7_75t_L g7945 ( 
.A(n_6837),
.Y(n_7945)
);

AOI22xp5_ASAP7_75t_L g7946 ( 
.A1(n_7697),
.A2(n_5749),
.B1(n_5872),
.B2(n_5821),
.Y(n_7946)
);

OR2x6_ASAP7_75t_L g7947 ( 
.A(n_7632),
.B(n_6410),
.Y(n_7947)
);

INVx5_ASAP7_75t_L g7948 ( 
.A(n_6751),
.Y(n_7948)
);

INVx2_ASAP7_75t_L g7949 ( 
.A(n_6746),
.Y(n_7949)
);

AOI22xp33_ASAP7_75t_L g7950 ( 
.A1(n_7026),
.A2(n_5821),
.B1(n_5919),
.B2(n_5818),
.Y(n_7950)
);

NAND2xp5_ASAP7_75t_L g7951 ( 
.A(n_7637),
.B(n_5838),
.Y(n_7951)
);

AOI21x1_ASAP7_75t_L g7952 ( 
.A1(n_7638),
.A2(n_6103),
.B(n_6044),
.Y(n_7952)
);

CKINVDCx11_ASAP7_75t_R g7953 ( 
.A(n_6999),
.Y(n_7953)
);

AND2x2_ASAP7_75t_L g7954 ( 
.A(n_6820),
.B(n_6847),
.Y(n_7954)
);

BUFx2_ASAP7_75t_L g7955 ( 
.A(n_7420),
.Y(n_7955)
);

A2O1A1Ixp33_ASAP7_75t_L g7956 ( 
.A1(n_7102),
.A2(n_5622),
.B(n_6515),
.C(n_5803),
.Y(n_7956)
);

OA21x2_ASAP7_75t_L g7957 ( 
.A1(n_7028),
.A2(n_7325),
.B(n_7212),
.Y(n_7957)
);

NOR2xp33_ASAP7_75t_L g7958 ( 
.A(n_6800),
.B(n_6198),
.Y(n_7958)
);

HB1xp67_ASAP7_75t_L g7959 ( 
.A(n_6890),
.Y(n_7959)
);

AOI21xp5_ASAP7_75t_L g7960 ( 
.A1(n_6709),
.A2(n_6242),
.B(n_6267),
.Y(n_7960)
);

AND2x4_ASAP7_75t_L g7961 ( 
.A(n_7318),
.B(n_5850),
.Y(n_7961)
);

INVx2_ASAP7_75t_L g7962 ( 
.A(n_6752),
.Y(n_7962)
);

AOI21xp33_ASAP7_75t_L g7963 ( 
.A1(n_7240),
.A2(n_6534),
.B(n_5714),
.Y(n_7963)
);

AND2x6_ASAP7_75t_L g7964 ( 
.A(n_6632),
.B(n_5230),
.Y(n_7964)
);

OAI21x1_ASAP7_75t_L g7965 ( 
.A1(n_6804),
.A2(n_6285),
.B(n_5840),
.Y(n_7965)
);

OAI21x1_ASAP7_75t_L g7966 ( 
.A1(n_6804),
.A2(n_6285),
.B(n_5840),
.Y(n_7966)
);

BUFx2_ASAP7_75t_L g7967 ( 
.A(n_7420),
.Y(n_7967)
);

OAI21x1_ASAP7_75t_L g7968 ( 
.A1(n_6845),
.A2(n_5837),
.B(n_6429),
.Y(n_7968)
);

INVx2_ASAP7_75t_L g7969 ( 
.A(n_6752),
.Y(n_7969)
);

O2A1O1Ixp33_ASAP7_75t_L g7970 ( 
.A1(n_6636),
.A2(n_6219),
.B(n_5651),
.C(n_5714),
.Y(n_7970)
);

INVx1_ASAP7_75t_L g7971 ( 
.A(n_6848),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_6848),
.Y(n_7972)
);

AO21x1_ASAP7_75t_L g7973 ( 
.A1(n_7600),
.A2(n_5849),
.B(n_6544),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_6848),
.Y(n_7974)
);

OA21x2_ASAP7_75t_L g7975 ( 
.A1(n_7028),
.A2(n_6361),
.B(n_6307),
.Y(n_7975)
);

INVx1_ASAP7_75t_L g7976 ( 
.A(n_6851),
.Y(n_7976)
);

BUFx6f_ASAP7_75t_L g7977 ( 
.A(n_6649),
.Y(n_7977)
);

INVx2_ASAP7_75t_SL g7978 ( 
.A(n_6649),
.Y(n_7978)
);

OAI22xp33_ASAP7_75t_L g7979 ( 
.A1(n_7672),
.A2(n_5863),
.B1(n_5878),
.B2(n_5811),
.Y(n_7979)
);

INVx1_ASAP7_75t_SL g7980 ( 
.A(n_6650),
.Y(n_7980)
);

OR2x2_ASAP7_75t_L g7981 ( 
.A(n_6820),
.B(n_6469),
.Y(n_7981)
);

INVx1_ASAP7_75t_L g7982 ( 
.A(n_6851),
.Y(n_7982)
);

CKINVDCx20_ASAP7_75t_R g7983 ( 
.A(n_6664),
.Y(n_7983)
);

NAND2x1p5_ASAP7_75t_L g7984 ( 
.A(n_7628),
.B(n_6694),
.Y(n_7984)
);

OAI22xp5_ASAP7_75t_L g7985 ( 
.A1(n_6694),
.A2(n_6904),
.B1(n_6899),
.B2(n_6896),
.Y(n_7985)
);

NAND2xp5_ASAP7_75t_SL g7986 ( 
.A(n_7101),
.B(n_5649),
.Y(n_7986)
);

OAI21x1_ASAP7_75t_L g7987 ( 
.A1(n_6845),
.A2(n_5837),
.B(n_6469),
.Y(n_7987)
);

OAI21x1_ASAP7_75t_SL g7988 ( 
.A1(n_6745),
.A2(n_7228),
.B(n_7033),
.Y(n_7988)
);

AOI22xp33_ASAP7_75t_L g7989 ( 
.A1(n_7026),
.A2(n_5818),
.B1(n_5538),
.B2(n_5715),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_6851),
.Y(n_7990)
);

INVx2_ASAP7_75t_L g7991 ( 
.A(n_6752),
.Y(n_7991)
);

BUFx5_ASAP7_75t_L g7992 ( 
.A(n_7079),
.Y(n_7992)
);

OAI21x1_ASAP7_75t_L g7993 ( 
.A1(n_7692),
.A2(n_6469),
.B(n_6125),
.Y(n_7993)
);

OAI21x1_ASAP7_75t_L g7994 ( 
.A1(n_7692),
.A2(n_6125),
.B(n_5733),
.Y(n_7994)
);

XNOR2xp5_ASAP7_75t_L g7995 ( 
.A(n_6764),
.B(n_6169),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_6865),
.Y(n_7996)
);

AO21x2_ASAP7_75t_L g7997 ( 
.A1(n_6662),
.A2(n_5766),
.B(n_6496),
.Y(n_7997)
);

AOI21x1_ASAP7_75t_L g7998 ( 
.A1(n_7692),
.A2(n_7470),
.B(n_6773),
.Y(n_7998)
);

AOI22xp33_ASAP7_75t_L g7999 ( 
.A1(n_7043),
.A2(n_5715),
.B1(n_5879),
.B2(n_6202),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_6865),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7637),
.B(n_5838),
.Y(n_8001)
);

AND2x2_ASAP7_75t_L g8002 ( 
.A(n_6847),
.B(n_6596),
.Y(n_8002)
);

CKINVDCx20_ASAP7_75t_R g8003 ( 
.A(n_6764),
.Y(n_8003)
);

OAI21x1_ASAP7_75t_SL g8004 ( 
.A1(n_6745),
.A2(n_5691),
.B(n_6524),
.Y(n_8004)
);

OA21x2_ASAP7_75t_L g8005 ( 
.A1(n_7049),
.A2(n_6361),
.B(n_6307),
.Y(n_8005)
);

AND2x2_ASAP7_75t_L g8006 ( 
.A(n_6847),
.B(n_6715),
.Y(n_8006)
);

INVx2_ASAP7_75t_L g8007 ( 
.A(n_6752),
.Y(n_8007)
);

AND2x4_ASAP7_75t_L g8008 ( 
.A(n_7121),
.B(n_5850),
.Y(n_8008)
);

OAI21xp5_ASAP7_75t_L g8009 ( 
.A1(n_7665),
.A2(n_7043),
.B(n_7697),
.Y(n_8009)
);

HB1xp67_ASAP7_75t_L g8010 ( 
.A(n_6909),
.Y(n_8010)
);

OAI21x1_ASAP7_75t_L g8011 ( 
.A1(n_7099),
.A2(n_5860),
.B(n_5711),
.Y(n_8011)
);

INVxp33_ASAP7_75t_L g8012 ( 
.A(n_6815),
.Y(n_8012)
);

INVx2_ASAP7_75t_L g8013 ( 
.A(n_6755),
.Y(n_8013)
);

NAND2xp5_ASAP7_75t_L g8014 ( 
.A(n_6828),
.B(n_5935),
.Y(n_8014)
);

OA21x2_ASAP7_75t_L g8015 ( 
.A1(n_7049),
.A2(n_6361),
.B(n_6307),
.Y(n_8015)
);

CKINVDCx11_ASAP7_75t_R g8016 ( 
.A(n_7129),
.Y(n_8016)
);

INVx2_ASAP7_75t_L g8017 ( 
.A(n_6755),
.Y(n_8017)
);

BUFx3_ASAP7_75t_L g8018 ( 
.A(n_6751),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_6865),
.Y(n_8019)
);

AOI22xp33_ASAP7_75t_L g8020 ( 
.A1(n_7043),
.A2(n_5879),
.B1(n_6206),
.B2(n_6202),
.Y(n_8020)
);

INVx2_ASAP7_75t_SL g8021 ( 
.A(n_6649),
.Y(n_8021)
);

INVx3_ASAP7_75t_L g8022 ( 
.A(n_6631),
.Y(n_8022)
);

BUFx2_ASAP7_75t_R g8023 ( 
.A(n_7316),
.Y(n_8023)
);

INVx8_ASAP7_75t_L g8024 ( 
.A(n_6795),
.Y(n_8024)
);

OAI21x1_ASAP7_75t_L g8025 ( 
.A1(n_7099),
.A2(n_5711),
.B(n_5707),
.Y(n_8025)
);

AO21x1_ASAP7_75t_L g8026 ( 
.A1(n_7600),
.A2(n_6544),
.B(n_6534),
.Y(n_8026)
);

A2O1A1Ixp33_ASAP7_75t_SL g8027 ( 
.A1(n_6979),
.A2(n_6451),
.B(n_5690),
.C(n_5732),
.Y(n_8027)
);

OAI22xp5_ASAP7_75t_L g8028 ( 
.A1(n_6694),
.A2(n_5717),
.B1(n_5662),
.B2(n_5574),
.Y(n_8028)
);

OAI21x1_ASAP7_75t_L g8029 ( 
.A1(n_7116),
.A2(n_7192),
.B(n_7214),
.Y(n_8029)
);

INVx1_ASAP7_75t_L g8030 ( 
.A(n_6866),
.Y(n_8030)
);

AND2x2_ASAP7_75t_L g8031 ( 
.A(n_6715),
.B(n_6596),
.Y(n_8031)
);

INVx1_ASAP7_75t_L g8032 ( 
.A(n_6866),
.Y(n_8032)
);

OAI21x1_ASAP7_75t_L g8033 ( 
.A1(n_7116),
.A2(n_7192),
.B(n_7214),
.Y(n_8033)
);

HB1xp67_ASAP7_75t_L g8034 ( 
.A(n_6909),
.Y(n_8034)
);

O2A1O1Ixp33_ASAP7_75t_SL g8035 ( 
.A1(n_6678),
.A2(n_6618),
.B(n_6568),
.C(n_6601),
.Y(n_8035)
);

OA21x2_ASAP7_75t_L g8036 ( 
.A1(n_7212),
.A2(n_6387),
.B(n_6375),
.Y(n_8036)
);

OA21x2_ASAP7_75t_L g8037 ( 
.A1(n_7622),
.A2(n_6387),
.B(n_6375),
.Y(n_8037)
);

INVx3_ASAP7_75t_L g8038 ( 
.A(n_6631),
.Y(n_8038)
);

INVx2_ASAP7_75t_L g8039 ( 
.A(n_6755),
.Y(n_8039)
);

INVx1_ASAP7_75t_L g8040 ( 
.A(n_6866),
.Y(n_8040)
);

OAI21x1_ASAP7_75t_L g8041 ( 
.A1(n_6662),
.A2(n_5722),
.B(n_5713),
.Y(n_8041)
);

OAI21x1_ASAP7_75t_L g8042 ( 
.A1(n_6668),
.A2(n_5722),
.B(n_5713),
.Y(n_8042)
);

BUFx2_ASAP7_75t_R g8043 ( 
.A(n_7316),
.Y(n_8043)
);

BUFx6f_ASAP7_75t_L g8044 ( 
.A(n_6649),
.Y(n_8044)
);

AND2x2_ASAP7_75t_L g8045 ( 
.A(n_6715),
.B(n_6609),
.Y(n_8045)
);

BUFx3_ASAP7_75t_L g8046 ( 
.A(n_6751),
.Y(n_8046)
);

AOI21xp5_ASAP7_75t_L g8047 ( 
.A1(n_6709),
.A2(n_6720),
.B(n_6684),
.Y(n_8047)
);

AND2x4_ASAP7_75t_L g8048 ( 
.A(n_7121),
.B(n_5850),
.Y(n_8048)
);

CKINVDCx5p33_ASAP7_75t_R g8049 ( 
.A(n_7394),
.Y(n_8049)
);

INVx6_ASAP7_75t_L g8050 ( 
.A(n_7331),
.Y(n_8050)
);

INVx2_ASAP7_75t_L g8051 ( 
.A(n_6755),
.Y(n_8051)
);

INVx1_ASAP7_75t_L g8052 ( 
.A(n_6880),
.Y(n_8052)
);

AND2x4_ASAP7_75t_L g8053 ( 
.A(n_7121),
.B(n_5850),
.Y(n_8053)
);

AOI22xp33_ASAP7_75t_L g8054 ( 
.A1(n_7697),
.A2(n_6221),
.B1(n_6230),
.B2(n_6206),
.Y(n_8054)
);

OAI21xp5_ASAP7_75t_L g8055 ( 
.A1(n_7665),
.A2(n_7209),
.B(n_7165),
.Y(n_8055)
);

OAI21xp5_ASAP7_75t_L g8056 ( 
.A1(n_7665),
.A2(n_5651),
.B(n_5691),
.Y(n_8056)
);

AND2x2_ASAP7_75t_L g8057 ( 
.A(n_6715),
.B(n_6609),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_6880),
.Y(n_8058)
);

OR2x6_ASAP7_75t_L g8059 ( 
.A(n_7632),
.B(n_6410),
.Y(n_8059)
);

INVx1_ASAP7_75t_L g8060 ( 
.A(n_6880),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_6882),
.Y(n_8061)
);

O2A1O1Ixp33_ASAP7_75t_L g8062 ( 
.A1(n_6636),
.A2(n_6219),
.B(n_5796),
.C(n_5776),
.Y(n_8062)
);

OAI22xp33_ASAP7_75t_L g8063 ( 
.A1(n_7672),
.A2(n_5863),
.B1(n_5878),
.B2(n_5811),
.Y(n_8063)
);

INVx2_ASAP7_75t_L g8064 ( 
.A(n_6783),
.Y(n_8064)
);

CKINVDCx5p33_ASAP7_75t_R g8065 ( 
.A(n_7394),
.Y(n_8065)
);

AOI22xp5_ASAP7_75t_L g8066 ( 
.A1(n_6920),
.A2(n_6077),
.B1(n_6084),
.B2(n_5705),
.Y(n_8066)
);

CKINVDCx20_ASAP7_75t_R g8067 ( 
.A(n_6788),
.Y(n_8067)
);

AND2x4_ASAP7_75t_L g8068 ( 
.A(n_7121),
.B(n_5850),
.Y(n_8068)
);

INVx4_ASAP7_75t_L g8069 ( 
.A(n_6750),
.Y(n_8069)
);

NAND2x1p5_ASAP7_75t_L g8070 ( 
.A(n_6694),
.B(n_5586),
.Y(n_8070)
);

AOI21xp33_ASAP7_75t_SL g8071 ( 
.A1(n_6697),
.A2(n_5895),
.B(n_6382),
.Y(n_8071)
);

OAI21x1_ASAP7_75t_L g8072 ( 
.A1(n_6656),
.A2(n_6759),
.B(n_6695),
.Y(n_8072)
);

CKINVDCx16_ASAP7_75t_R g8073 ( 
.A(n_6750),
.Y(n_8073)
);

AOI21xp5_ASAP7_75t_L g8074 ( 
.A1(n_6720),
.A2(n_6242),
.B(n_6267),
.Y(n_8074)
);

HB1xp67_ASAP7_75t_L g8075 ( 
.A(n_6974),
.Y(n_8075)
);

OR2x2_ASAP7_75t_L g8076 ( 
.A(n_6818),
.B(n_6624),
.Y(n_8076)
);

OAI21x1_ASAP7_75t_L g8077 ( 
.A1(n_6695),
.A2(n_6759),
.B(n_6956),
.Y(n_8077)
);

AOI21xp5_ASAP7_75t_L g8078 ( 
.A1(n_6677),
.A2(n_6684),
.B(n_6756),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_6882),
.Y(n_8079)
);

INVx1_ASAP7_75t_L g8080 ( 
.A(n_6882),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_6889),
.Y(n_8081)
);

BUFx6f_ASAP7_75t_L g8082 ( 
.A(n_6649),
.Y(n_8082)
);

AND2x4_ASAP7_75t_L g8083 ( 
.A(n_7155),
.B(n_5859),
.Y(n_8083)
);

NOR2xp33_ASAP7_75t_L g8084 ( 
.A(n_7122),
.B(n_6221),
.Y(n_8084)
);

INVx2_ASAP7_75t_SL g8085 ( 
.A(n_6649),
.Y(n_8085)
);

AOI22xp33_ASAP7_75t_L g8086 ( 
.A1(n_6896),
.A2(n_6230),
.B1(n_5690),
.B2(n_5732),
.Y(n_8086)
);

AO31x2_ASAP7_75t_L g8087 ( 
.A1(n_7033),
.A2(n_7387),
.A3(n_7377),
.B(n_7566),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_6889),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_6889),
.Y(n_8089)
);

AOI22xp33_ASAP7_75t_L g8090 ( 
.A1(n_6920),
.A2(n_6169),
.B1(n_5803),
.B2(n_6082),
.Y(n_8090)
);

INVx2_ASAP7_75t_L g8091 ( 
.A(n_6783),
.Y(n_8091)
);

CKINVDCx11_ASAP7_75t_R g8092 ( 
.A(n_7129),
.Y(n_8092)
);

CKINVDCx11_ASAP7_75t_R g8093 ( 
.A(n_6750),
.Y(n_8093)
);

OR2x2_ASAP7_75t_L g8094 ( 
.A(n_6818),
.B(n_5652),
.Y(n_8094)
);

AO21x2_ASAP7_75t_L g8095 ( 
.A1(n_6705),
.A2(n_5712),
.B(n_6318),
.Y(n_8095)
);

INVx1_ASAP7_75t_SL g8096 ( 
.A(n_6650),
.Y(n_8096)
);

AO31x2_ASAP7_75t_L g8097 ( 
.A1(n_7033),
.A2(n_6174),
.A3(n_6194),
.B(n_6141),
.Y(n_8097)
);

OA21x2_ASAP7_75t_L g8098 ( 
.A1(n_7622),
.A2(n_6387),
.B(n_6375),
.Y(n_8098)
);

AND2x4_ASAP7_75t_L g8099 ( 
.A(n_7155),
.B(n_5859),
.Y(n_8099)
);

NAND2x1p5_ASAP7_75t_L g8100 ( 
.A(n_7209),
.B(n_5803),
.Y(n_8100)
);

HB1xp67_ASAP7_75t_L g8101 ( 
.A(n_6974),
.Y(n_8101)
);

INVx1_ASAP7_75t_L g8102 ( 
.A(n_6905),
.Y(n_8102)
);

INVx2_ASAP7_75t_SL g8103 ( 
.A(n_6649),
.Y(n_8103)
);

AND2x2_ASAP7_75t_L g8104 ( 
.A(n_6715),
.B(n_5859),
.Y(n_8104)
);

OAI22xp33_ASAP7_75t_L g8105 ( 
.A1(n_7672),
.A2(n_5649),
.B1(n_5811),
.B2(n_5803),
.Y(n_8105)
);

OAI21x1_ASAP7_75t_L g8106 ( 
.A1(n_6695),
.A2(n_6613),
.B(n_5928),
.Y(n_8106)
);

AOI21x1_ASAP7_75t_L g8107 ( 
.A1(n_7470),
.A2(n_6103),
.B(n_6044),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_6905),
.Y(n_8108)
);

OAI21xp5_ASAP7_75t_L g8109 ( 
.A1(n_7209),
.A2(n_5796),
.B(n_6077),
.Y(n_8109)
);

NOR2x1_ASAP7_75t_SL g8110 ( 
.A(n_7382),
.B(n_5747),
.Y(n_8110)
);

HB1xp67_ASAP7_75t_L g8111 ( 
.A(n_7012),
.Y(n_8111)
);

INVx1_ASAP7_75t_L g8112 ( 
.A(n_6905),
.Y(n_8112)
);

CKINVDCx5p33_ASAP7_75t_R g8113 ( 
.A(n_6740),
.Y(n_8113)
);

BUFx6f_ASAP7_75t_L g8114 ( 
.A(n_6649),
.Y(n_8114)
);

AND2x2_ASAP7_75t_L g8115 ( 
.A(n_6715),
.B(n_5859),
.Y(n_8115)
);

INVxp67_ASAP7_75t_L g8116 ( 
.A(n_6644),
.Y(n_8116)
);

AOI22xp5_ASAP7_75t_L g8117 ( 
.A1(n_6899),
.A2(n_6084),
.B1(n_5705),
.B2(n_6108),
.Y(n_8117)
);

OAI21x1_ASAP7_75t_L g8118 ( 
.A1(n_6695),
.A2(n_6613),
.B(n_5928),
.Y(n_8118)
);

BUFx3_ASAP7_75t_L g8119 ( 
.A(n_6751),
.Y(n_8119)
);

OAI21x1_ASAP7_75t_L g8120 ( 
.A1(n_6759),
.A2(n_6613),
.B(n_5928),
.Y(n_8120)
);

AO31x2_ASAP7_75t_L g8121 ( 
.A1(n_7387),
.A2(n_6174),
.A3(n_6194),
.B(n_6141),
.Y(n_8121)
);

A2O1A1Ixp33_ASAP7_75t_L g8122 ( 
.A1(n_6719),
.A2(n_6082),
.B(n_5803),
.C(n_6108),
.Y(n_8122)
);

HB1xp67_ASAP7_75t_SL g8123 ( 
.A(n_7264),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_6913),
.Y(n_8124)
);

OAI21xp5_ASAP7_75t_L g8125 ( 
.A1(n_7165),
.A2(n_6498),
.B(n_5712),
.Y(n_8125)
);

BUFx4f_ASAP7_75t_L g8126 ( 
.A(n_6835),
.Y(n_8126)
);

OAI21x1_ASAP7_75t_L g8127 ( 
.A1(n_6759),
.A2(n_5928),
.B(n_5924),
.Y(n_8127)
);

AOI22xp33_ASAP7_75t_SL g8128 ( 
.A1(n_7047),
.A2(n_6778),
.B1(n_6819),
.B2(n_6932),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_6913),
.Y(n_8129)
);

OAI221xp5_ASAP7_75t_L g8130 ( 
.A1(n_7144),
.A2(n_6451),
.B1(n_6470),
.B2(n_6426),
.C(n_6431),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_6913),
.Y(n_8131)
);

INVx2_ASAP7_75t_L g8132 ( 
.A(n_6783),
.Y(n_8132)
);

BUFx3_ASAP7_75t_L g8133 ( 
.A(n_6751),
.Y(n_8133)
);

OAI21x1_ASAP7_75t_L g8134 ( 
.A1(n_6759),
.A2(n_5928),
.B(n_5924),
.Y(n_8134)
);

INVx1_ASAP7_75t_SL g8135 ( 
.A(n_6699),
.Y(n_8135)
);

AOI22xp33_ASAP7_75t_SL g8136 ( 
.A1(n_7047),
.A2(n_6082),
.B1(n_6219),
.B2(n_6473),
.Y(n_8136)
);

OAI21x1_ASAP7_75t_L g8137 ( 
.A1(n_6956),
.A2(n_5936),
.B(n_5924),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_6917),
.Y(n_8138)
);

AOI221xp5_ASAP7_75t_L g8139 ( 
.A1(n_6886),
.A2(n_6311),
.B1(n_6313),
.B2(n_6287),
.C(n_6279),
.Y(n_8139)
);

OAI21x1_ASAP7_75t_L g8140 ( 
.A1(n_6956),
.A2(n_5936),
.B(n_5924),
.Y(n_8140)
);

INVx2_ASAP7_75t_L g8141 ( 
.A(n_6783),
.Y(n_8141)
);

OAI21x1_ASAP7_75t_L g8142 ( 
.A1(n_6956),
.A2(n_5992),
.B(n_5936),
.Y(n_8142)
);

NAND2xp5_ASAP7_75t_L g8143 ( 
.A(n_6828),
.B(n_5935),
.Y(n_8143)
);

AND2x2_ASAP7_75t_L g8144 ( 
.A(n_6743),
.B(n_5859),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_6832),
.Y(n_8145)
);

OAI21x1_ASAP7_75t_L g8146 ( 
.A1(n_6956),
.A2(n_5992),
.B(n_5936),
.Y(n_8146)
);

AOI22xp33_ASAP7_75t_L g8147 ( 
.A1(n_7213),
.A2(n_6082),
.B1(n_5689),
.B2(n_6380),
.Y(n_8147)
);

INVx4_ASAP7_75t_L g8148 ( 
.A(n_6795),
.Y(n_8148)
);

OAI21xp5_ASAP7_75t_L g8149 ( 
.A1(n_7144),
.A2(n_6498),
.B(n_5627),
.Y(n_8149)
);

OAI21x1_ASAP7_75t_L g8150 ( 
.A1(n_7292),
.A2(n_5992),
.B(n_5936),
.Y(n_8150)
);

AOI22xp5_ASAP7_75t_SL g8151 ( 
.A1(n_7274),
.A2(n_6129),
.B1(n_6172),
.B2(n_5898),
.Y(n_8151)
);

AO21x1_ASAP7_75t_L g8152 ( 
.A1(n_6778),
.A2(n_5689),
.B(n_6329),
.Y(n_8152)
);

OAI21x1_ASAP7_75t_SL g8153 ( 
.A1(n_7228),
.A2(n_6524),
.B(n_6380),
.Y(n_8153)
);

BUFx2_ASAP7_75t_L g8154 ( 
.A(n_7420),
.Y(n_8154)
);

INVx1_ASAP7_75t_L g8155 ( 
.A(n_6917),
.Y(n_8155)
);

OA21x2_ASAP7_75t_L g8156 ( 
.A1(n_7667),
.A2(n_6391),
.B(n_5972),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_6917),
.Y(n_8157)
);

CKINVDCx5p33_ASAP7_75t_R g8158 ( 
.A(n_6794),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_6919),
.Y(n_8159)
);

OR2x6_ASAP7_75t_L g8160 ( 
.A(n_7632),
.B(n_7154),
.Y(n_8160)
);

OA21x2_ASAP7_75t_L g8161 ( 
.A1(n_7667),
.A2(n_6391),
.B(n_5972),
.Y(n_8161)
);

OR2x6_ASAP7_75t_L g8162 ( 
.A(n_7632),
.B(n_6410),
.Y(n_8162)
);

O2A1O1Ixp33_ASAP7_75t_SL g8163 ( 
.A1(n_6719),
.A2(n_6568),
.B(n_6601),
.C(n_6573),
.Y(n_8163)
);

OAI21xp5_ASAP7_75t_L g8164 ( 
.A1(n_7144),
.A2(n_6933),
.B(n_7137),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_6832),
.Y(n_8165)
);

AO21x2_ASAP7_75t_L g8166 ( 
.A1(n_6705),
.A2(n_6329),
.B(n_5845),
.Y(n_8166)
);

NOR2x1_ASAP7_75t_SL g8167 ( 
.A(n_7386),
.B(n_5747),
.Y(n_8167)
);

OAI21x1_ASAP7_75t_L g8168 ( 
.A1(n_7292),
.A2(n_5999),
.B(n_5992),
.Y(n_8168)
);

AND2x2_ASAP7_75t_L g8169 ( 
.A(n_6743),
.B(n_5859),
.Y(n_8169)
);

HB1xp67_ASAP7_75t_L g8170 ( 
.A(n_7012),
.Y(n_8170)
);

NAND2xp5_ASAP7_75t_L g8171 ( 
.A(n_6828),
.B(n_5954),
.Y(n_8171)
);

AOI22xp5_ASAP7_75t_L g8172 ( 
.A1(n_6904),
.A2(n_5868),
.B1(n_6473),
.B2(n_5767),
.Y(n_8172)
);

OAI21x1_ASAP7_75t_L g8173 ( 
.A1(n_7292),
.A2(n_5999),
.B(n_5992),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_6919),
.Y(n_8174)
);

OAI21x1_ASAP7_75t_L g8175 ( 
.A1(n_7292),
.A2(n_6023),
.B(n_5999),
.Y(n_8175)
);

OAI21x1_ASAP7_75t_L g8176 ( 
.A1(n_7292),
.A2(n_6023),
.B(n_5999),
.Y(n_8176)
);

OAI21x1_ASAP7_75t_L g8177 ( 
.A1(n_7688),
.A2(n_6023),
.B(n_5999),
.Y(n_8177)
);

OAI21x1_ASAP7_75t_L g8178 ( 
.A1(n_7688),
.A2(n_6026),
.B(n_6023),
.Y(n_8178)
);

AOI21xp5_ASAP7_75t_L g8179 ( 
.A1(n_6677),
.A2(n_6242),
.B(n_6267),
.Y(n_8179)
);

INVx2_ASAP7_75t_L g8180 ( 
.A(n_6832),
.Y(n_8180)
);

AOI21xp5_ASAP7_75t_L g8181 ( 
.A1(n_6756),
.A2(n_6242),
.B(n_6267),
.Y(n_8181)
);

OAI21x1_ASAP7_75t_SL g8182 ( 
.A1(n_7228),
.A2(n_6524),
.B(n_5767),
.Y(n_8182)
);

OAI21x1_ASAP7_75t_L g8183 ( 
.A1(n_6891),
.A2(n_6026),
.B(n_6023),
.Y(n_8183)
);

A2O1A1Ixp33_ASAP7_75t_L g8184 ( 
.A1(n_7137),
.A2(n_7345),
.B(n_7063),
.C(n_7105),
.Y(n_8184)
);

NAND2xp5_ASAP7_75t_L g8185 ( 
.A(n_6801),
.B(n_5954),
.Y(n_8185)
);

INVx3_ASAP7_75t_L g8186 ( 
.A(n_6631),
.Y(n_8186)
);

BUFx2_ASAP7_75t_L g8187 ( 
.A(n_7420),
.Y(n_8187)
);

OA21x2_ASAP7_75t_L g8188 ( 
.A1(n_7703),
.A2(n_6391),
.B(n_5972),
.Y(n_8188)
);

BUFx3_ASAP7_75t_L g8189 ( 
.A(n_6751),
.Y(n_8189)
);

NAND2xp5_ASAP7_75t_L g8190 ( 
.A(n_6801),
.B(n_5967),
.Y(n_8190)
);

BUFx6f_ASAP7_75t_L g8191 ( 
.A(n_6649),
.Y(n_8191)
);

OAI22xp33_ASAP7_75t_L g8192 ( 
.A1(n_7345),
.A2(n_5649),
.B1(n_5811),
.B2(n_6082),
.Y(n_8192)
);

AOI21x1_ASAP7_75t_L g8193 ( 
.A1(n_7470),
.A2(n_6103),
.B(n_6129),
.Y(n_8193)
);

AOI22xp33_ASAP7_75t_L g8194 ( 
.A1(n_7213),
.A2(n_5667),
.B1(n_6470),
.B2(n_5699),
.Y(n_8194)
);

AOI22xp5_ASAP7_75t_L g8195 ( 
.A1(n_6819),
.A2(n_5868),
.B1(n_6495),
.B2(n_6313),
.Y(n_8195)
);

OR2x2_ASAP7_75t_L g8196 ( 
.A(n_6818),
.B(n_5652),
.Y(n_8196)
);

BUFx3_ASAP7_75t_L g8197 ( 
.A(n_6751),
.Y(n_8197)
);

OR2x2_ASAP7_75t_L g8198 ( 
.A(n_6818),
.B(n_5658),
.Y(n_8198)
);

AND2x4_ASAP7_75t_L g8199 ( 
.A(n_7155),
.B(n_5859),
.Y(n_8199)
);

AOI22xp33_ASAP7_75t_L g8200 ( 
.A1(n_7213),
.A2(n_5667),
.B1(n_5699),
.B2(n_5686),
.Y(n_8200)
);

CKINVDCx11_ASAP7_75t_R g8201 ( 
.A(n_6795),
.Y(n_8201)
);

NOR2xp33_ASAP7_75t_L g8202 ( 
.A(n_7122),
.B(n_5568),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_6919),
.Y(n_8203)
);

OAI21x1_ASAP7_75t_L g8204 ( 
.A1(n_7200),
.A2(n_6068),
.B(n_6055),
.Y(n_8204)
);

INVx3_ASAP7_75t_L g8205 ( 
.A(n_6631),
.Y(n_8205)
);

AO21x2_ASAP7_75t_L g8206 ( 
.A1(n_7607),
.A2(n_5845),
.B(n_6132),
.Y(n_8206)
);

OAI21x1_ASAP7_75t_L g8207 ( 
.A1(n_7200),
.A2(n_6068),
.B(n_6055),
.Y(n_8207)
);

OR2x6_ASAP7_75t_L g8208 ( 
.A(n_7632),
.B(n_7154),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_6922),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_6922),
.Y(n_8210)
);

OAI21xp5_ASAP7_75t_L g8211 ( 
.A1(n_6933),
.A2(n_6587),
.B(n_6356),
.Y(n_8211)
);

OAI21x1_ASAP7_75t_SL g8212 ( 
.A1(n_7595),
.A2(n_6587),
.B(n_6471),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_6801),
.B(n_5967),
.Y(n_8213)
);

O2A1O1Ixp33_ASAP7_75t_L g8214 ( 
.A1(n_6636),
.A2(n_6219),
.B(n_5776),
.C(n_5848),
.Y(n_8214)
);

INVx4_ASAP7_75t_L g8215 ( 
.A(n_6795),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_6922),
.Y(n_8216)
);

OAI21x1_ASAP7_75t_L g8217 ( 
.A1(n_6774),
.A2(n_6088),
.B(n_6080),
.Y(n_8217)
);

OAI21xp5_ASAP7_75t_L g8218 ( 
.A1(n_6933),
.A2(n_6356),
.B(n_6351),
.Y(n_8218)
);

O2A1O1Ixp33_ASAP7_75t_L g8219 ( 
.A1(n_6636),
.A2(n_5848),
.B(n_6357),
.C(n_6351),
.Y(n_8219)
);

NAND3xp33_ASAP7_75t_L g8220 ( 
.A(n_7227),
.B(n_6370),
.C(n_6357),
.Y(n_8220)
);

OAI21xp5_ASAP7_75t_L g8221 ( 
.A1(n_6886),
.A2(n_6390),
.B(n_6370),
.Y(n_8221)
);

BUFx2_ASAP7_75t_L g8222 ( 
.A(n_7420),
.Y(n_8222)
);

INVxp67_ASAP7_75t_L g8223 ( 
.A(n_6644),
.Y(n_8223)
);

OAI21xp5_ASAP7_75t_L g8224 ( 
.A1(n_7003),
.A2(n_6390),
.B(n_6495),
.Y(n_8224)
);

AOI21xp5_ASAP7_75t_L g8225 ( 
.A1(n_6651),
.A2(n_6267),
.B(n_6410),
.Y(n_8225)
);

HB1xp67_ASAP7_75t_L g8226 ( 
.A(n_7054),
.Y(n_8226)
);

OA21x2_ASAP7_75t_L g8227 ( 
.A1(n_7152),
.A2(n_5996),
.B(n_5962),
.Y(n_8227)
);

INVx2_ASAP7_75t_SL g8228 ( 
.A(n_6686),
.Y(n_8228)
);

AOI21x1_ASAP7_75t_L g8229 ( 
.A1(n_6773),
.A2(n_6979),
.B(n_7655),
.Y(n_8229)
);

BUFx3_ASAP7_75t_L g8230 ( 
.A(n_6817),
.Y(n_8230)
);

CKINVDCx5p33_ASAP7_75t_R g8231 ( 
.A(n_6794),
.Y(n_8231)
);

AOI221xp5_ASAP7_75t_L g8232 ( 
.A1(n_6932),
.A2(n_6778),
.B1(n_6819),
.B2(n_6647),
.C(n_7503),
.Y(n_8232)
);

OAI21x1_ASAP7_75t_L g8233 ( 
.A1(n_6774),
.A2(n_6088),
.B(n_6080),
.Y(n_8233)
);

O2A1O1Ixp5_ASAP7_75t_L g8234 ( 
.A1(n_7063),
.A2(n_7196),
.B(n_7164),
.C(n_7091),
.Y(n_8234)
);

AOI21xp5_ASAP7_75t_SL g8235 ( 
.A1(n_7595),
.A2(n_6518),
.B(n_6507),
.Y(n_8235)
);

INVx2_ASAP7_75t_L g8236 ( 
.A(n_6832),
.Y(n_8236)
);

CKINVDCx8_ASAP7_75t_R g8237 ( 
.A(n_6697),
.Y(n_8237)
);

AOI21x1_ASAP7_75t_L g8238 ( 
.A1(n_6773),
.A2(n_5996),
.B(n_5962),
.Y(n_8238)
);

BUFx2_ASAP7_75t_R g8239 ( 
.A(n_7490),
.Y(n_8239)
);

OAI21x1_ASAP7_75t_L g8240 ( 
.A1(n_6774),
.A2(n_6089),
.B(n_6088),
.Y(n_8240)
);

OAI221xp5_ASAP7_75t_L g8241 ( 
.A1(n_6809),
.A2(n_6426),
.B1(n_6431),
.B2(n_6382),
.C(n_6499),
.Y(n_8241)
);

CKINVDCx11_ASAP7_75t_R g8242 ( 
.A(n_6811),
.Y(n_8242)
);

BUFx3_ASAP7_75t_L g8243 ( 
.A(n_6817),
.Y(n_8243)
);

OAI21x1_ASAP7_75t_L g8244 ( 
.A1(n_6774),
.A2(n_6089),
.B(n_6088),
.Y(n_8244)
);

OAI21x1_ASAP7_75t_L g8245 ( 
.A1(n_6774),
.A2(n_6089),
.B(n_6088),
.Y(n_8245)
);

AOI221xp5_ASAP7_75t_L g8246 ( 
.A1(n_6932),
.A2(n_6385),
.B1(n_6362),
.B2(n_6279),
.C(n_6494),
.Y(n_8246)
);

OAI21x1_ASAP7_75t_L g8247 ( 
.A1(n_6937),
.A2(n_6092),
.B(n_6089),
.Y(n_8247)
);

NAND2x1p5_ASAP7_75t_L g8248 ( 
.A(n_6686),
.B(n_5829),
.Y(n_8248)
);

BUFx3_ASAP7_75t_L g8249 ( 
.A(n_6817),
.Y(n_8249)
);

OAI21x1_ASAP7_75t_L g8250 ( 
.A1(n_6937),
.A2(n_6092),
.B(n_6089),
.Y(n_8250)
);

NOR2xp33_ASAP7_75t_L g8251 ( 
.A(n_7122),
.B(n_5568),
.Y(n_8251)
);

OAI21x1_ASAP7_75t_L g8252 ( 
.A1(n_6937),
.A2(n_6093),
.B(n_6092),
.Y(n_8252)
);

INVx2_ASAP7_75t_L g8253 ( 
.A(n_6836),
.Y(n_8253)
);

NOR2xp67_ASAP7_75t_L g8254 ( 
.A(n_7475),
.B(n_5548),
.Y(n_8254)
);

INVx1_ASAP7_75t_L g8255 ( 
.A(n_6949),
.Y(n_8255)
);

OAI21x1_ASAP7_75t_L g8256 ( 
.A1(n_6937),
.A2(n_6093),
.B(n_6092),
.Y(n_8256)
);

OAI22xp5_ASAP7_75t_L g8257 ( 
.A1(n_6842),
.A2(n_6857),
.B1(n_6674),
.B2(n_7474),
.Y(n_8257)
);

AO21x2_ASAP7_75t_L g8258 ( 
.A1(n_7607),
.A2(n_5845),
.B(n_6133),
.Y(n_8258)
);

NAND2xp5_ASAP7_75t_L g8259 ( 
.A(n_7666),
.B(n_6013),
.Y(n_8259)
);

INVx1_ASAP7_75t_L g8260 ( 
.A(n_6949),
.Y(n_8260)
);

NAND2xp5_ASAP7_75t_L g8261 ( 
.A(n_7666),
.B(n_6013),
.Y(n_8261)
);

OAI21x1_ASAP7_75t_L g8262 ( 
.A1(n_6937),
.A2(n_6093),
.B(n_6092),
.Y(n_8262)
);

OAI22xp5_ASAP7_75t_L g8263 ( 
.A1(n_6842),
.A2(n_5789),
.B1(n_6096),
.B2(n_5574),
.Y(n_8263)
);

AO31x2_ASAP7_75t_L g8264 ( 
.A1(n_7377),
.A2(n_6174),
.A3(n_6194),
.B(n_6141),
.Y(n_8264)
);

INVx1_ASAP7_75t_L g8265 ( 
.A(n_6949),
.Y(n_8265)
);

OAI21x1_ASAP7_75t_L g8266 ( 
.A1(n_6952),
.A2(n_6112),
.B(n_6093),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_6957),
.Y(n_8267)
);

INVx2_ASAP7_75t_L g8268 ( 
.A(n_6836),
.Y(n_8268)
);

INVx1_ASAP7_75t_L g8269 ( 
.A(n_6957),
.Y(n_8269)
);

INVx3_ASAP7_75t_L g8270 ( 
.A(n_6631),
.Y(n_8270)
);

OAI21x1_ASAP7_75t_L g8271 ( 
.A1(n_6952),
.A2(n_6112),
.B(n_6093),
.Y(n_8271)
);

AND2x2_ASAP7_75t_L g8272 ( 
.A(n_6743),
.B(n_5859),
.Y(n_8272)
);

HB1xp67_ASAP7_75t_L g8273 ( 
.A(n_7054),
.Y(n_8273)
);

INVx2_ASAP7_75t_SL g8274 ( 
.A(n_6686),
.Y(n_8274)
);

OAI22xp5_ASAP7_75t_L g8275 ( 
.A1(n_6857),
.A2(n_5789),
.B1(n_6096),
.B2(n_5574),
.Y(n_8275)
);

AO31x2_ASAP7_75t_L g8276 ( 
.A1(n_7566),
.A2(n_6214),
.A3(n_6217),
.B(n_6213),
.Y(n_8276)
);

OAI21xp5_ASAP7_75t_L g8277 ( 
.A1(n_7003),
.A2(n_6499),
.B(n_6494),
.Y(n_8277)
);

BUFx6f_ASAP7_75t_L g8278 ( 
.A(n_6686),
.Y(n_8278)
);

OAI21x1_ASAP7_75t_L g8279 ( 
.A1(n_6952),
.A2(n_6154),
.B(n_6112),
.Y(n_8279)
);

INVxp67_ASAP7_75t_L g8280 ( 
.A(n_6673),
.Y(n_8280)
);

CKINVDCx5p33_ASAP7_75t_R g8281 ( 
.A(n_7493),
.Y(n_8281)
);

BUFx6f_ASAP7_75t_L g8282 ( 
.A(n_6686),
.Y(n_8282)
);

INVx1_ASAP7_75t_L g8283 ( 
.A(n_6957),
.Y(n_8283)
);

OAI22xp5_ASAP7_75t_L g8284 ( 
.A1(n_6674),
.A2(n_7479),
.B1(n_7474),
.B2(n_6841),
.Y(n_8284)
);

NOR2x1_ASAP7_75t_SL g8285 ( 
.A(n_7386),
.B(n_5747),
.Y(n_8285)
);

OAI21x1_ASAP7_75t_L g8286 ( 
.A1(n_6952),
.A2(n_6154),
.B(n_6112),
.Y(n_8286)
);

BUFx2_ASAP7_75t_L g8287 ( 
.A(n_7420),
.Y(n_8287)
);

INVx3_ASAP7_75t_L g8288 ( 
.A(n_6631),
.Y(n_8288)
);

O2A1O1Ixp33_ASAP7_75t_SL g8289 ( 
.A1(n_7408),
.A2(n_6563),
.B(n_6518),
.C(n_6559),
.Y(n_8289)
);

BUFx2_ASAP7_75t_L g8290 ( 
.A(n_7420),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_6985),
.Y(n_8291)
);

OAI221xp5_ASAP7_75t_L g8292 ( 
.A1(n_6809),
.A2(n_6875),
.B1(n_6897),
.B2(n_6841),
.C(n_6813),
.Y(n_8292)
);

NAND2x1p5_ASAP7_75t_L g8293 ( 
.A(n_6686),
.B(n_5831),
.Y(n_8293)
);

AOI22xp5_ASAP7_75t_L g8294 ( 
.A1(n_7227),
.A2(n_6385),
.B1(n_6362),
.B2(n_6535),
.Y(n_8294)
);

INVx2_ASAP7_75t_L g8295 ( 
.A(n_6836),
.Y(n_8295)
);

AOI21xp5_ASAP7_75t_L g8296 ( 
.A1(n_6651),
.A2(n_6410),
.B(n_6453),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_6985),
.Y(n_8297)
);

INVxp67_ASAP7_75t_L g8298 ( 
.A(n_6673),
.Y(n_8298)
);

AOI22xp33_ASAP7_75t_L g8299 ( 
.A1(n_7227),
.A2(n_7115),
.B1(n_7457),
.B2(n_7419),
.Y(n_8299)
);

AO21x1_ASAP7_75t_L g8300 ( 
.A1(n_7091),
.A2(n_5852),
.B(n_5709),
.Y(n_8300)
);

OAI21x1_ASAP7_75t_L g8301 ( 
.A1(n_6952),
.A2(n_6154),
.B(n_6112),
.Y(n_8301)
);

NOR2xp33_ASAP7_75t_L g8302 ( 
.A(n_7356),
.B(n_5591),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_6985),
.Y(n_8303)
);

AOI21x1_ASAP7_75t_L g8304 ( 
.A1(n_7655),
.A2(n_5998),
.B(n_5996),
.Y(n_8304)
);

INVx2_ASAP7_75t_L g8305 ( 
.A(n_6836),
.Y(n_8305)
);

INVx1_ASAP7_75t_L g8306 ( 
.A(n_6988),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_6988),
.Y(n_8307)
);

CKINVDCx20_ASAP7_75t_R g8308 ( 
.A(n_6788),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_6988),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_6992),
.Y(n_8310)
);

INVx2_ASAP7_75t_SL g8311 ( 
.A(n_6686),
.Y(n_8311)
);

AND2x2_ASAP7_75t_L g8312 ( 
.A(n_6743),
.B(n_5869),
.Y(n_8312)
);

AO21x1_ASAP7_75t_L g8313 ( 
.A1(n_7386),
.A2(n_7544),
.B(n_7496),
.Y(n_8313)
);

INVx1_ASAP7_75t_L g8314 ( 
.A(n_6992),
.Y(n_8314)
);

OAI22xp5_ASAP7_75t_L g8315 ( 
.A1(n_7474),
.A2(n_6096),
.B1(n_6563),
.B2(n_6471),
.Y(n_8315)
);

NAND2xp5_ASAP7_75t_L g8316 ( 
.A(n_7077),
.B(n_6022),
.Y(n_8316)
);

OA21x2_ASAP7_75t_L g8317 ( 
.A1(n_7152),
.A2(n_6016),
.B(n_5998),
.Y(n_8317)
);

INVx2_ASAP7_75t_SL g8318 ( 
.A(n_6686),
.Y(n_8318)
);

OAI21xp5_ASAP7_75t_L g8319 ( 
.A1(n_7003),
.A2(n_6535),
.B(n_6548),
.Y(n_8319)
);

OA21x2_ASAP7_75t_L g8320 ( 
.A1(n_7393),
.A2(n_6016),
.B(n_5998),
.Y(n_8320)
);

AOI22xp5_ASAP7_75t_L g8321 ( 
.A1(n_6647),
.A2(n_6873),
.B1(n_6858),
.B2(n_7164),
.Y(n_8321)
);

NOR2xp33_ASAP7_75t_L g8322 ( 
.A(n_7356),
.B(n_5591),
.Y(n_8322)
);

NAND2x1p5_ASAP7_75t_L g8323 ( 
.A(n_6686),
.B(n_5831),
.Y(n_8323)
);

OAI21x1_ASAP7_75t_L g8324 ( 
.A1(n_7433),
.A2(n_6228),
.B(n_6164),
.Y(n_8324)
);

AOI22xp33_ASAP7_75t_L g8325 ( 
.A1(n_7115),
.A2(n_5709),
.B1(n_5686),
.B2(n_6616),
.Y(n_8325)
);

OAI221xp5_ASAP7_75t_L g8326 ( 
.A1(n_6809),
.A2(n_6512),
.B1(n_6525),
.B2(n_6509),
.C(n_5836),
.Y(n_8326)
);

AOI21x1_ASAP7_75t_L g8327 ( 
.A1(n_7646),
.A2(n_6031),
.B(n_6016),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_L g8328 ( 
.A(n_7077),
.B(n_6022),
.Y(n_8328)
);

BUFx6f_ASAP7_75t_L g8329 ( 
.A(n_6686),
.Y(n_8329)
);

NAND3xp33_ASAP7_75t_SL g8330 ( 
.A(n_6636),
.B(n_5669),
.C(n_5620),
.Y(n_8330)
);

INVx3_ASAP7_75t_L g8331 ( 
.A(n_6631),
.Y(n_8331)
);

OAI22xp5_ASAP7_75t_L g8332 ( 
.A1(n_7474),
.A2(n_6507),
.B1(n_6559),
.B2(n_6543),
.Y(n_8332)
);

INVx1_ASAP7_75t_L g8333 ( 
.A(n_6992),
.Y(n_8333)
);

INVx2_ASAP7_75t_SL g8334 ( 
.A(n_6796),
.Y(n_8334)
);

NAND2x1p5_ASAP7_75t_L g8335 ( 
.A(n_6796),
.B(n_6895),
.Y(n_8335)
);

AO32x2_ASAP7_75t_L g8336 ( 
.A1(n_7341),
.A2(n_6620),
.A3(n_6617),
.B1(n_5909),
.B2(n_5921),
.Y(n_8336)
);

NAND2xp5_ASAP7_75t_L g8337 ( 
.A(n_7077),
.B(n_6050),
.Y(n_8337)
);

OAI21xp5_ASAP7_75t_L g8338 ( 
.A1(n_7475),
.A2(n_6548),
.B(n_5847),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_6996),
.Y(n_8339)
);

BUFx6f_ASAP7_75t_L g8340 ( 
.A(n_6796),
.Y(n_8340)
);

INVx1_ASAP7_75t_L g8341 ( 
.A(n_6996),
.Y(n_8341)
);

AND2x2_ASAP7_75t_L g8342 ( 
.A(n_6768),
.B(n_5869),
.Y(n_8342)
);

INVx1_ASAP7_75t_L g8343 ( 
.A(n_6996),
.Y(n_8343)
);

AOI21xp33_ASAP7_75t_L g8344 ( 
.A1(n_7419),
.A2(n_6058),
.B(n_6050),
.Y(n_8344)
);

INVx1_ASAP7_75t_L g8345 ( 
.A(n_6997),
.Y(n_8345)
);

NAND2x1p5_ASAP7_75t_L g8346 ( 
.A(n_6796),
.B(n_6895),
.Y(n_8346)
);

HB1xp67_ASAP7_75t_L g8347 ( 
.A(n_7064),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_6997),
.Y(n_8348)
);

OAI21x1_ASAP7_75t_L g8349 ( 
.A1(n_7433),
.A2(n_6228),
.B(n_6164),
.Y(n_8349)
);

OAI21x1_ASAP7_75t_L g8350 ( 
.A1(n_7433),
.A2(n_6259),
.B(n_6228),
.Y(n_8350)
);

CKINVDCx8_ASAP7_75t_R g8351 ( 
.A(n_6726),
.Y(n_8351)
);

AO21x2_ASAP7_75t_L g8352 ( 
.A1(n_7607),
.A2(n_5845),
.B(n_6133),
.Y(n_8352)
);

INVx2_ASAP7_75t_SL g8353 ( 
.A(n_6796),
.Y(n_8353)
);

INVx5_ASAP7_75t_L g8354 ( 
.A(n_6817),
.Y(n_8354)
);

AOI222xp33_ASAP7_75t_L g8355 ( 
.A1(n_6858),
.A2(n_6186),
.B1(n_6126),
.B2(n_6246),
.C1(n_6130),
.C2(n_6109),
.Y(n_8355)
);

OAI21x1_ASAP7_75t_L g8356 ( 
.A1(n_7433),
.A2(n_6259),
.B(n_6228),
.Y(n_8356)
);

INVx2_ASAP7_75t_SL g8357 ( 
.A(n_6796),
.Y(n_8357)
);

NOR3xp33_ASAP7_75t_SL g8358 ( 
.A(n_6622),
.B(n_6671),
.C(n_6814),
.Y(n_8358)
);

OA21x2_ASAP7_75t_L g8359 ( 
.A1(n_7223),
.A2(n_6214),
.B(n_6213),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_6997),
.Y(n_8360)
);

NAND2xp5_ASAP7_75t_L g8361 ( 
.A(n_7090),
.B(n_7098),
.Y(n_8361)
);

INVx6_ASAP7_75t_L g8362 ( 
.A(n_7331),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_7016),
.Y(n_8363)
);

AOI22xp33_ASAP7_75t_L g8364 ( 
.A1(n_7419),
.A2(n_7457),
.B1(n_7409),
.B2(n_7005),
.Y(n_8364)
);

AOI221xp5_ASAP7_75t_L g8365 ( 
.A1(n_6647),
.A2(n_6035),
.B1(n_6081),
.B2(n_6072),
.C(n_6066),
.Y(n_8365)
);

NAND2x1p5_ASAP7_75t_L g8366 ( 
.A(n_6796),
.B(n_5831),
.Y(n_8366)
);

HB1xp67_ASAP7_75t_L g8367 ( 
.A(n_7064),
.Y(n_8367)
);

BUFx8_ASAP7_75t_L g8368 ( 
.A(n_6811),
.Y(n_8368)
);

OA21x2_ASAP7_75t_L g8369 ( 
.A1(n_6850),
.A2(n_6031),
.B(n_6213),
.Y(n_8369)
);

AOI21xp5_ASAP7_75t_L g8370 ( 
.A1(n_6651),
.A2(n_6467),
.B(n_6453),
.Y(n_8370)
);

INVx3_ASAP7_75t_L g8371 ( 
.A(n_6663),
.Y(n_8371)
);

OAI21x1_ASAP7_75t_L g8372 ( 
.A1(n_7433),
.A2(n_7546),
.B(n_7440),
.Y(n_8372)
);

OAI21x1_ASAP7_75t_L g8373 ( 
.A1(n_7440),
.A2(n_6280),
.B(n_6259),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_7016),
.Y(n_8374)
);

AND2x2_ASAP7_75t_L g8375 ( 
.A(n_6768),
.B(n_5869),
.Y(n_8375)
);

HB1xp67_ASAP7_75t_L g8376 ( 
.A(n_7080),
.Y(n_8376)
);

AND2x2_ASAP7_75t_L g8377 ( 
.A(n_6768),
.B(n_5869),
.Y(n_8377)
);

NOR2xp33_ASAP7_75t_L g8378 ( 
.A(n_7356),
.B(n_5620),
.Y(n_8378)
);

OAI21x1_ASAP7_75t_L g8379 ( 
.A1(n_7440),
.A2(n_6280),
.B(n_6259),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7016),
.Y(n_8380)
);

OAI21x1_ASAP7_75t_L g8381 ( 
.A1(n_7440),
.A2(n_6280),
.B(n_6259),
.Y(n_8381)
);

AOI22xp33_ASAP7_75t_L g8382 ( 
.A1(n_7457),
.A2(n_6616),
.B1(n_5760),
.B2(n_6130),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_7025),
.Y(n_8383)
);

INVx3_ASAP7_75t_L g8384 ( 
.A(n_6663),
.Y(n_8384)
);

AOI22xp33_ASAP7_75t_L g8385 ( 
.A1(n_7409),
.A2(n_6616),
.B1(n_5760),
.B2(n_6130),
.Y(n_8385)
);

INVx8_ASAP7_75t_L g8386 ( 
.A(n_6811),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7025),
.Y(n_8387)
);

INVx2_ASAP7_75t_L g8388 ( 
.A(n_6843),
.Y(n_8388)
);

OAI21x1_ASAP7_75t_L g8389 ( 
.A1(n_7440),
.A2(n_6315),
.B(n_6280),
.Y(n_8389)
);

INVx2_ASAP7_75t_SL g8390 ( 
.A(n_6796),
.Y(n_8390)
);

AND2x2_ASAP7_75t_L g8391 ( 
.A(n_6768),
.B(n_5869),
.Y(n_8391)
);

HB1xp67_ASAP7_75t_L g8392 ( 
.A(n_7080),
.Y(n_8392)
);

AND2x2_ASAP7_75t_L g8393 ( 
.A(n_6799),
.B(n_5869),
.Y(n_8393)
);

OAI22xp5_ASAP7_75t_L g8394 ( 
.A1(n_7479),
.A2(n_5895),
.B1(n_6120),
.B2(n_6102),
.Y(n_8394)
);

AND2x2_ASAP7_75t_L g8395 ( 
.A(n_6799),
.B(n_5869),
.Y(n_8395)
);

AND2x4_ASAP7_75t_L g8396 ( 
.A(n_7155),
.B(n_5869),
.Y(n_8396)
);

AOI221xp5_ASAP7_75t_L g8397 ( 
.A1(n_7503),
.A2(n_6858),
.B1(n_6873),
.B2(n_7271),
.C(n_7538),
.Y(n_8397)
);

AOI21xp5_ASAP7_75t_L g8398 ( 
.A1(n_6879),
.A2(n_6467),
.B(n_6453),
.Y(n_8398)
);

OR2x6_ASAP7_75t_L g8399 ( 
.A(n_7154),
.B(n_6527),
.Y(n_8399)
);

INVx5_ASAP7_75t_L g8400 ( 
.A(n_6817),
.Y(n_8400)
);

NAND2xp33_ASAP7_75t_R g8401 ( 
.A(n_7339),
.B(n_6590),
.Y(n_8401)
);

NOR2xp33_ASAP7_75t_L g8402 ( 
.A(n_7066),
.B(n_7219),
.Y(n_8402)
);

INVx2_ASAP7_75t_SL g8403 ( 
.A(n_6796),
.Y(n_8403)
);

BUFx2_ASAP7_75t_SL g8404 ( 
.A(n_6823),
.Y(n_8404)
);

OA21x2_ASAP7_75t_L g8405 ( 
.A1(n_7223),
.A2(n_6217),
.B(n_6214),
.Y(n_8405)
);

AOI22xp33_ASAP7_75t_L g8406 ( 
.A1(n_7409),
.A2(n_5760),
.B1(n_6186),
.B2(n_6126),
.Y(n_8406)
);

AOI221xp5_ASAP7_75t_L g8407 ( 
.A1(n_7503),
.A2(n_6619),
.B1(n_6066),
.B2(n_6081),
.C(n_6072),
.Y(n_8407)
);

INVx2_ASAP7_75t_SL g8408 ( 
.A(n_6796),
.Y(n_8408)
);

NAND2xp5_ASAP7_75t_L g8409 ( 
.A(n_7090),
.B(n_7098),
.Y(n_8409)
);

INVx1_ASAP7_75t_L g8410 ( 
.A(n_7025),
.Y(n_8410)
);

OAI21x1_ASAP7_75t_L g8411 ( 
.A1(n_7546),
.A2(n_6315),
.B(n_6280),
.Y(n_8411)
);

INVx2_ASAP7_75t_L g8412 ( 
.A(n_6843),
.Y(n_8412)
);

NAND2xp5_ASAP7_75t_L g8413 ( 
.A(n_7090),
.B(n_6058),
.Y(n_8413)
);

OAI22xp5_ASAP7_75t_L g8414 ( 
.A1(n_7479),
.A2(n_6120),
.B1(n_6207),
.B2(n_6102),
.Y(n_8414)
);

BUFx5_ASAP7_75t_L g8415 ( 
.A(n_7079),
.Y(n_8415)
);

AO21x1_ASAP7_75t_L g8416 ( 
.A1(n_7496),
.A2(n_5852),
.B(n_6135),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_7031),
.Y(n_8417)
);

INVx1_ASAP7_75t_SL g8418 ( 
.A(n_6699),
.Y(n_8418)
);

OAI21x1_ASAP7_75t_L g8419 ( 
.A1(n_7546),
.A2(n_6325),
.B(n_6315),
.Y(n_8419)
);

O2A1O1Ixp33_ASAP7_75t_SL g8420 ( 
.A1(n_7408),
.A2(n_5680),
.B(n_5737),
.C(n_5669),
.Y(n_8420)
);

INVx3_ASAP7_75t_L g8421 ( 
.A(n_6663),
.Y(n_8421)
);

OAI21x1_ASAP7_75t_L g8422 ( 
.A1(n_7546),
.A2(n_6325),
.B(n_6315),
.Y(n_8422)
);

INVx3_ASAP7_75t_L g8423 ( 
.A(n_6663),
.Y(n_8423)
);

BUFx3_ASAP7_75t_L g8424 ( 
.A(n_6817),
.Y(n_8424)
);

OAI21x1_ASAP7_75t_L g8425 ( 
.A1(n_7546),
.A2(n_6325),
.B(n_6315),
.Y(n_8425)
);

NAND3xp33_ASAP7_75t_L g8426 ( 
.A(n_6722),
.B(n_6512),
.C(n_6509),
.Y(n_8426)
);

O2A1O1Ixp33_ASAP7_75t_SL g8427 ( 
.A1(n_7454),
.A2(n_5737),
.B(n_5680),
.C(n_6355),
.Y(n_8427)
);

AOI21xp5_ASAP7_75t_L g8428 ( 
.A1(n_6879),
.A2(n_6467),
.B(n_6453),
.Y(n_8428)
);

INVx8_ASAP7_75t_L g8429 ( 
.A(n_6811),
.Y(n_8429)
);

OR2x2_ASAP7_75t_L g8430 ( 
.A(n_6624),
.B(n_5658),
.Y(n_8430)
);

OAI21x1_ASAP7_75t_SL g8431 ( 
.A1(n_7640),
.A2(n_5628),
.B(n_5610),
.Y(n_8431)
);

INVx1_ASAP7_75t_L g8432 ( 
.A(n_7031),
.Y(n_8432)
);

OAI21xp5_ASAP7_75t_L g8433 ( 
.A1(n_7475),
.A2(n_5847),
.B(n_5774),
.Y(n_8433)
);

INVx2_ASAP7_75t_SL g8434 ( 
.A(n_6895),
.Y(n_8434)
);

INVx1_ASAP7_75t_SL g8435 ( 
.A(n_6699),
.Y(n_8435)
);

AND2x4_ASAP7_75t_L g8436 ( 
.A(n_7184),
.B(n_5880),
.Y(n_8436)
);

OA21x2_ASAP7_75t_L g8437 ( 
.A1(n_6758),
.A2(n_6222),
.B(n_6217),
.Y(n_8437)
);

A2O1A1Ixp33_ASAP7_75t_L g8438 ( 
.A1(n_7345),
.A2(n_6363),
.B(n_6394),
.C(n_6355),
.Y(n_8438)
);

INVx1_ASAP7_75t_SL g8439 ( 
.A(n_7092),
.Y(n_8439)
);

OR2x2_ASAP7_75t_L g8440 ( 
.A(n_6624),
.B(n_6584),
.Y(n_8440)
);

OR2x6_ASAP7_75t_L g8441 ( 
.A(n_7154),
.B(n_5735),
.Y(n_8441)
);

BUFx3_ASAP7_75t_L g8442 ( 
.A(n_6817),
.Y(n_8442)
);

INVx2_ASAP7_75t_L g8443 ( 
.A(n_6843),
.Y(n_8443)
);

BUFx2_ASAP7_75t_R g8444 ( 
.A(n_7490),
.Y(n_8444)
);

INVx1_ASAP7_75t_L g8445 ( 
.A(n_7031),
.Y(n_8445)
);

CKINVDCx5p33_ASAP7_75t_R g8446 ( 
.A(n_7493),
.Y(n_8446)
);

AOI21xp5_ASAP7_75t_L g8447 ( 
.A1(n_6665),
.A2(n_6467),
.B(n_6453),
.Y(n_8447)
);

INVx2_ASAP7_75t_L g8448 ( 
.A(n_6843),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_7038),
.Y(n_8449)
);

INVx1_ASAP7_75t_L g8450 ( 
.A(n_7038),
.Y(n_8450)
);

AND2x2_ASAP7_75t_L g8451 ( 
.A(n_6799),
.B(n_5880),
.Y(n_8451)
);

OAI22xp5_ASAP7_75t_L g8452 ( 
.A1(n_7479),
.A2(n_6120),
.B1(n_6207),
.B2(n_6102),
.Y(n_8452)
);

AOI22xp33_ASAP7_75t_L g8453 ( 
.A1(n_7005),
.A2(n_6186),
.B1(n_6246),
.B2(n_6126),
.Y(n_8453)
);

AO21x2_ASAP7_75t_L g8454 ( 
.A1(n_6758),
.A2(n_6147),
.B(n_6143),
.Y(n_8454)
);

INVx2_ASAP7_75t_L g8455 ( 
.A(n_6860),
.Y(n_8455)
);

OAI21x1_ASAP7_75t_L g8456 ( 
.A1(n_7681),
.A2(n_6327),
.B(n_6325),
.Y(n_8456)
);

BUFx2_ASAP7_75t_L g8457 ( 
.A(n_7420),
.Y(n_8457)
);

O2A1O1Ixp33_ASAP7_75t_L g8458 ( 
.A1(n_7060),
.A2(n_5706),
.B(n_6086),
.C(n_6035),
.Y(n_8458)
);

AOI21xp5_ASAP7_75t_SL g8459 ( 
.A1(n_7640),
.A2(n_5960),
.B(n_5891),
.Y(n_8459)
);

INVx1_ASAP7_75t_L g8460 ( 
.A(n_7038),
.Y(n_8460)
);

NOR2xp33_ASAP7_75t_L g8461 ( 
.A(n_7066),
.B(n_6215),
.Y(n_8461)
);

NOR2xp33_ASAP7_75t_L g8462 ( 
.A(n_7219),
.B(n_6215),
.Y(n_8462)
);

INVx3_ASAP7_75t_L g8463 ( 
.A(n_6663),
.Y(n_8463)
);

HB1xp67_ASAP7_75t_L g8464 ( 
.A(n_7096),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7044),
.Y(n_8465)
);

OAI21x1_ASAP7_75t_L g8466 ( 
.A1(n_7681),
.A2(n_6327),
.B(n_6325),
.Y(n_8466)
);

NAND3xp33_ASAP7_75t_L g8467 ( 
.A(n_6722),
.B(n_6525),
.C(n_5642),
.Y(n_8467)
);

BUFx2_ASAP7_75t_L g8468 ( 
.A(n_7079),
.Y(n_8468)
);

AOI21x1_ASAP7_75t_L g8469 ( 
.A1(n_7646),
.A2(n_6031),
.B(n_6222),
.Y(n_8469)
);

INVx1_ASAP7_75t_L g8470 ( 
.A(n_7044),
.Y(n_8470)
);

OAI22xp5_ASAP7_75t_L g8471 ( 
.A1(n_6813),
.A2(n_6207),
.B1(n_5556),
.B2(n_5563),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_6860),
.Y(n_8472)
);

O2A1O1Ixp33_ASAP7_75t_L g8473 ( 
.A1(n_7060),
.A2(n_5706),
.B(n_6105),
.C(n_6086),
.Y(n_8473)
);

NAND2xp5_ASAP7_75t_L g8474 ( 
.A(n_7098),
.B(n_6397),
.Y(n_8474)
);

OAI21x1_ASAP7_75t_L g8475 ( 
.A1(n_7681),
.A2(n_6386),
.B(n_6327),
.Y(n_8475)
);

AOI21xp5_ASAP7_75t_L g8476 ( 
.A1(n_6665),
.A2(n_6467),
.B(n_6453),
.Y(n_8476)
);

AND2x2_ASAP7_75t_L g8477 ( 
.A(n_6799),
.B(n_5880),
.Y(n_8477)
);

AND2x4_ASAP7_75t_L g8478 ( 
.A(n_7184),
.B(n_5880),
.Y(n_8478)
);

AND2x4_ASAP7_75t_L g8479 ( 
.A(n_7184),
.B(n_5880),
.Y(n_8479)
);

INVx2_ASAP7_75t_L g8480 ( 
.A(n_6860),
.Y(n_8480)
);

INVx4_ASAP7_75t_L g8481 ( 
.A(n_6993),
.Y(n_8481)
);

OAI21x1_ASAP7_75t_L g8482 ( 
.A1(n_7681),
.A2(n_6386),
.B(n_6327),
.Y(n_8482)
);

BUFx6f_ASAP7_75t_L g8483 ( 
.A(n_6895),
.Y(n_8483)
);

NAND2xp5_ASAP7_75t_L g8484 ( 
.A(n_7687),
.B(n_6397),
.Y(n_8484)
);

OAI21xp5_ASAP7_75t_L g8485 ( 
.A1(n_7594),
.A2(n_5774),
.B(n_5772),
.Y(n_8485)
);

AND2x2_ASAP7_75t_L g8486 ( 
.A(n_6834),
.B(n_5880),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7044),
.Y(n_8487)
);

OA21x2_ASAP7_75t_L g8488 ( 
.A1(n_7172),
.A2(n_6223),
.B(n_6222),
.Y(n_8488)
);

NAND2xp5_ASAP7_75t_L g8489 ( 
.A(n_7687),
.B(n_6446),
.Y(n_8489)
);

AND2x4_ASAP7_75t_L g8490 ( 
.A(n_7184),
.B(n_7289),
.Y(n_8490)
);

INVx1_ASAP7_75t_SL g8491 ( 
.A(n_7092),
.Y(n_8491)
);

OAI21x1_ASAP7_75t_L g8492 ( 
.A1(n_7681),
.A2(n_6386),
.B(n_6327),
.Y(n_8492)
);

OAI21x1_ASAP7_75t_L g8493 ( 
.A1(n_7695),
.A2(n_6436),
.B(n_6386),
.Y(n_8493)
);

BUFx6f_ASAP7_75t_L g8494 ( 
.A(n_6895),
.Y(n_8494)
);

NAND2xp5_ASAP7_75t_L g8495 ( 
.A(n_7687),
.B(n_6446),
.Y(n_8495)
);

INVx2_ASAP7_75t_SL g8496 ( 
.A(n_6895),
.Y(n_8496)
);

NOR2xp33_ASAP7_75t_L g8497 ( 
.A(n_7235),
.B(n_6502),
.Y(n_8497)
);

OAI21x1_ASAP7_75t_L g8498 ( 
.A1(n_7695),
.A2(n_6436),
.B(n_6386),
.Y(n_8498)
);

OAI21xp5_ASAP7_75t_L g8499 ( 
.A1(n_7594),
.A2(n_5772),
.B(n_5637),
.Y(n_8499)
);

INVx2_ASAP7_75t_L g8500 ( 
.A(n_6860),
.Y(n_8500)
);

AO21x2_ASAP7_75t_L g8501 ( 
.A1(n_7172),
.A2(n_6147),
.B(n_6143),
.Y(n_8501)
);

OAI21x1_ASAP7_75t_L g8502 ( 
.A1(n_7695),
.A2(n_6437),
.B(n_6436),
.Y(n_8502)
);

AND2x2_ASAP7_75t_L g8503 ( 
.A(n_6834),
.B(n_5880),
.Y(n_8503)
);

INVxp67_ASAP7_75t_L g8504 ( 
.A(n_6736),
.Y(n_8504)
);

OAI22xp5_ASAP7_75t_L g8505 ( 
.A1(n_7649),
.A2(n_5556),
.B1(n_5563),
.B2(n_5535),
.Y(n_8505)
);

OA21x2_ASAP7_75t_L g8506 ( 
.A1(n_7172),
.A2(n_6232),
.B(n_6223),
.Y(n_8506)
);

AO22x2_ASAP7_75t_L g8507 ( 
.A1(n_7625),
.A2(n_5548),
.B1(n_5588),
.B2(n_5554),
.Y(n_8507)
);

OAI22x1_ASAP7_75t_L g8508 ( 
.A1(n_6875),
.A2(n_5636),
.B1(n_5856),
.B2(n_5592),
.Y(n_8508)
);

AND2x2_ASAP7_75t_L g8509 ( 
.A(n_6834),
.B(n_5880),
.Y(n_8509)
);

INVx1_ASAP7_75t_L g8510 ( 
.A(n_7046),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_6864),
.Y(n_8511)
);

AOI22xp33_ASAP7_75t_SL g8512 ( 
.A1(n_7047),
.A2(n_5790),
.B1(n_5820),
.B2(n_5677),
.Y(n_8512)
);

NAND2xp5_ASAP7_75t_L g8513 ( 
.A(n_7689),
.B(n_6502),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_7046),
.Y(n_8514)
);

OAI21x1_ASAP7_75t_L g8515 ( 
.A1(n_7695),
.A2(n_6437),
.B(n_6436),
.Y(n_8515)
);

O2A1O1Ixp33_ASAP7_75t_L g8516 ( 
.A1(n_7060),
.A2(n_5706),
.B(n_6105),
.C(n_6098),
.Y(n_8516)
);

OAI21xp5_ASAP7_75t_L g8517 ( 
.A1(n_7594),
.A2(n_5637),
.B(n_5630),
.Y(n_8517)
);

INVxp67_ASAP7_75t_SL g8518 ( 
.A(n_6643),
.Y(n_8518)
);

NAND2xp5_ASAP7_75t_L g8519 ( 
.A(n_7689),
.B(n_6558),
.Y(n_8519)
);

AND2x4_ASAP7_75t_L g8520 ( 
.A(n_7289),
.B(n_7322),
.Y(n_8520)
);

NOR2xp33_ASAP7_75t_L g8521 ( 
.A(n_7235),
.B(n_7234),
.Y(n_8521)
);

AO21x2_ASAP7_75t_L g8522 ( 
.A1(n_7482),
.A2(n_6173),
.B(n_6158),
.Y(n_8522)
);

OAI21x1_ASAP7_75t_L g8523 ( 
.A1(n_7695),
.A2(n_6437),
.B(n_6436),
.Y(n_8523)
);

BUFx2_ASAP7_75t_L g8524 ( 
.A(n_7079),
.Y(n_8524)
);

INVx1_ASAP7_75t_L g8525 ( 
.A(n_7046),
.Y(n_8525)
);

BUFx6f_ASAP7_75t_L g8526 ( 
.A(n_6895),
.Y(n_8526)
);

NOR2xp33_ASAP7_75t_L g8527 ( 
.A(n_7234),
.B(n_6558),
.Y(n_8527)
);

AND2x4_ASAP7_75t_L g8528 ( 
.A(n_7289),
.B(n_5893),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_7050),
.Y(n_8529)
);

BUFx6f_ASAP7_75t_L g8530 ( 
.A(n_6895),
.Y(n_8530)
);

INVx4_ASAP7_75t_L g8531 ( 
.A(n_6993),
.Y(n_8531)
);

NAND2xp5_ASAP7_75t_L g8532 ( 
.A(n_7689),
.B(n_7698),
.Y(n_8532)
);

NAND3xp33_ASAP7_75t_L g8533 ( 
.A(n_7271),
.B(n_5642),
.C(n_5640),
.Y(n_8533)
);

AOI21x1_ASAP7_75t_L g8534 ( 
.A1(n_7544),
.A2(n_6232),
.B(n_6223),
.Y(n_8534)
);

AO32x2_ASAP7_75t_L g8535 ( 
.A1(n_7341),
.A2(n_6620),
.A3(n_6617),
.B1(n_5909),
.B2(n_5921),
.Y(n_8535)
);

OA21x2_ASAP7_75t_L g8536 ( 
.A1(n_7482),
.A2(n_6240),
.B(n_6232),
.Y(n_8536)
);

BUFx8_ASAP7_75t_L g8537 ( 
.A(n_6993),
.Y(n_8537)
);

NOR2xp67_ASAP7_75t_L g8538 ( 
.A(n_7156),
.B(n_5548),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_7050),
.Y(n_8539)
);

HB1xp67_ASAP7_75t_L g8540 ( 
.A(n_7096),
.Y(n_8540)
);

NOR2xp33_ASAP7_75t_L g8541 ( 
.A(n_7010),
.B(n_6155),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_7050),
.Y(n_8542)
);

AOI221xp5_ASAP7_75t_L g8543 ( 
.A1(n_6873),
.A2(n_7562),
.B1(n_7538),
.B2(n_6874),
.C(n_6862),
.Y(n_8543)
);

AOI22xp5_ASAP7_75t_L g8544 ( 
.A1(n_7196),
.A2(n_6394),
.B1(n_6363),
.B2(n_6561),
.Y(n_8544)
);

AOI22xp33_ASAP7_75t_L g8545 ( 
.A1(n_6861),
.A2(n_6320),
.B1(n_6403),
.B2(n_6246),
.Y(n_8545)
);

CKINVDCx5p33_ASAP7_75t_R g8546 ( 
.A(n_6671),
.Y(n_8546)
);

AND2x2_ASAP7_75t_L g8547 ( 
.A(n_6834),
.B(n_5893),
.Y(n_8547)
);

INVx2_ASAP7_75t_L g8548 ( 
.A(n_6864),
.Y(n_8548)
);

BUFx2_ASAP7_75t_L g8549 ( 
.A(n_7079),
.Y(n_8549)
);

OA21x2_ASAP7_75t_L g8550 ( 
.A1(n_7482),
.A2(n_7512),
.B(n_7381),
.Y(n_8550)
);

AO21x1_ASAP7_75t_L g8551 ( 
.A1(n_7579),
.A2(n_7633),
.B(n_7598),
.Y(n_8551)
);

NAND2xp5_ASAP7_75t_L g8552 ( 
.A(n_7698),
.B(n_6584),
.Y(n_8552)
);

O2A1O1Ixp33_ASAP7_75t_SL g8553 ( 
.A1(n_7454),
.A2(n_6574),
.B(n_6561),
.C(n_6611),
.Y(n_8553)
);

NOR2xp33_ASAP7_75t_L g8554 ( 
.A(n_7010),
.B(n_6155),
.Y(n_8554)
);

INVx2_ASAP7_75t_L g8555 ( 
.A(n_6864),
.Y(n_8555)
);

NAND2xp5_ASAP7_75t_L g8556 ( 
.A(n_7698),
.B(n_6603),
.Y(n_8556)
);

OAI21x1_ASAP7_75t_L g8557 ( 
.A1(n_7250),
.A2(n_6472),
.B(n_6441),
.Y(n_8557)
);

INVx2_ASAP7_75t_SL g8558 ( 
.A(n_6895),
.Y(n_8558)
);

BUFx6f_ASAP7_75t_L g8559 ( 
.A(n_6895),
.Y(n_8559)
);

AND2x4_ASAP7_75t_L g8560 ( 
.A(n_7289),
.B(n_5893),
.Y(n_8560)
);

OAI21x1_ASAP7_75t_L g8561 ( 
.A1(n_7250),
.A2(n_6480),
.B(n_6472),
.Y(n_8561)
);

AOI22xp33_ASAP7_75t_L g8562 ( 
.A1(n_6861),
.A2(n_6403),
.B1(n_6425),
.B2(n_6320),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_7051),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_7051),
.Y(n_8564)
);

OR2x6_ASAP7_75t_L g8565 ( 
.A(n_7154),
.B(n_5827),
.Y(n_8565)
);

OAI21x1_ASAP7_75t_L g8566 ( 
.A1(n_7250),
.A2(n_6480),
.B(n_6472),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7051),
.Y(n_8567)
);

BUFx6f_ASAP7_75t_L g8568 ( 
.A(n_6908),
.Y(n_8568)
);

NAND2x1p5_ASAP7_75t_L g8569 ( 
.A(n_6908),
.B(n_5831),
.Y(n_8569)
);

INVx1_ASAP7_75t_L g8570 ( 
.A(n_7053),
.Y(n_8570)
);

OAI21x1_ASAP7_75t_L g8571 ( 
.A1(n_6725),
.A2(n_6484),
.B(n_6480),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_7053),
.Y(n_8572)
);

CKINVDCx20_ASAP7_75t_R g8573 ( 
.A(n_6839),
.Y(n_8573)
);

NAND2xp5_ASAP7_75t_L g8574 ( 
.A(n_6672),
.B(n_6603),
.Y(n_8574)
);

OA21x2_ASAP7_75t_L g8575 ( 
.A1(n_7381),
.A2(n_6256),
.B(n_6240),
.Y(n_8575)
);

OAI22xp5_ASAP7_75t_L g8576 ( 
.A1(n_7649),
.A2(n_5563),
.B1(n_5589),
.B2(n_5556),
.Y(n_8576)
);

INVx2_ASAP7_75t_L g8577 ( 
.A(n_6864),
.Y(n_8577)
);

OAI21x1_ASAP7_75t_L g8578 ( 
.A1(n_6725),
.A2(n_6484),
.B(n_6480),
.Y(n_8578)
);

INVx1_ASAP7_75t_L g8579 ( 
.A(n_7053),
.Y(n_8579)
);

BUFx3_ASAP7_75t_L g8580 ( 
.A(n_6817),
.Y(n_8580)
);

INVx3_ASAP7_75t_L g8581 ( 
.A(n_6663),
.Y(n_8581)
);

INVx2_ASAP7_75t_L g8582 ( 
.A(n_6871),
.Y(n_8582)
);

OAI21x1_ASAP7_75t_L g8583 ( 
.A1(n_6725),
.A2(n_6805),
.B(n_7517),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_7065),
.Y(n_8584)
);

NAND2x1p5_ASAP7_75t_L g8585 ( 
.A(n_6908),
.B(n_5831),
.Y(n_8585)
);

BUFx2_ASAP7_75t_SL g8586 ( 
.A(n_6823),
.Y(n_8586)
);

OAI21x1_ASAP7_75t_SL g8587 ( 
.A1(n_7105),
.A2(n_5628),
.B(n_5610),
.Y(n_8587)
);

BUFx2_ASAP7_75t_L g8588 ( 
.A(n_7079),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_6871),
.Y(n_8589)
);

AO21x2_ASAP7_75t_L g8590 ( 
.A1(n_7270),
.A2(n_6173),
.B(n_6158),
.Y(n_8590)
);

OAI21x1_ASAP7_75t_L g8591 ( 
.A1(n_6805),
.A2(n_6484),
.B(n_6480),
.Y(n_8591)
);

AND2x4_ASAP7_75t_L g8592 ( 
.A(n_7322),
.B(n_5893),
.Y(n_8592)
);

INVx5_ASAP7_75t_L g8593 ( 
.A(n_6817),
.Y(n_8593)
);

OR2x2_ASAP7_75t_L g8594 ( 
.A(n_7191),
.B(n_7201),
.Y(n_8594)
);

BUFx6f_ASAP7_75t_L g8595 ( 
.A(n_6908),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_7065),
.Y(n_8596)
);

OAI21x1_ASAP7_75t_L g8597 ( 
.A1(n_6805),
.A2(n_6485),
.B(n_6484),
.Y(n_8597)
);

OAI21x1_ASAP7_75t_SL g8598 ( 
.A1(n_7105),
.A2(n_5628),
.B(n_5610),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_7065),
.Y(n_8599)
);

INVx1_ASAP7_75t_L g8600 ( 
.A(n_7068),
.Y(n_8600)
);

OAI21x1_ASAP7_75t_L g8601 ( 
.A1(n_7517),
.A2(n_6485),
.B(n_6484),
.Y(n_8601)
);

INVx2_ASAP7_75t_L g8602 ( 
.A(n_6871),
.Y(n_8602)
);

BUFx3_ASAP7_75t_L g8603 ( 
.A(n_6817),
.Y(n_8603)
);

AO21x2_ASAP7_75t_L g8604 ( 
.A1(n_7270),
.A2(n_6184),
.B(n_6177),
.Y(n_8604)
);

NAND2xp5_ASAP7_75t_L g8605 ( 
.A(n_6672),
.B(n_6611),
.Y(n_8605)
);

BUFx6f_ASAP7_75t_L g8606 ( 
.A(n_6908),
.Y(n_8606)
);

INVx2_ASAP7_75t_L g8607 ( 
.A(n_6871),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_7068),
.Y(n_8608)
);

AO21x2_ASAP7_75t_L g8609 ( 
.A1(n_7388),
.A2(n_6184),
.B(n_6177),
.Y(n_8609)
);

O2A1O1Ixp33_ASAP7_75t_L g8610 ( 
.A1(n_7060),
.A2(n_5706),
.B(n_6111),
.C(n_6098),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_7068),
.Y(n_8611)
);

NOR2x1_ASAP7_75t_R g8612 ( 
.A(n_6993),
.B(n_6320),
.Y(n_8612)
);

OAI21x1_ASAP7_75t_L g8613 ( 
.A1(n_7022),
.A2(n_7626),
.B(n_7311),
.Y(n_8613)
);

NAND2xp5_ASAP7_75t_SL g8614 ( 
.A(n_6840),
.B(n_5893),
.Y(n_8614)
);

BUFx2_ASAP7_75t_L g8615 ( 
.A(n_7079),
.Y(n_8615)
);

OAI22xp5_ASAP7_75t_L g8616 ( 
.A1(n_6960),
.A2(n_5589),
.B1(n_5601),
.B2(n_5563),
.Y(n_8616)
);

AOI21xp5_ASAP7_75t_L g8617 ( 
.A1(n_6665),
.A2(n_6467),
.B(n_6453),
.Y(n_8617)
);

INVx1_ASAP7_75t_L g8618 ( 
.A(n_7072),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_7072),
.Y(n_8619)
);

INVx1_ASAP7_75t_L g8620 ( 
.A(n_7072),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_7074),
.Y(n_8621)
);

AOI21xp5_ASAP7_75t_L g8622 ( 
.A1(n_6782),
.A2(n_6555),
.B(n_6467),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_6893),
.Y(n_8623)
);

AO21x2_ASAP7_75t_L g8624 ( 
.A1(n_7388),
.A2(n_6204),
.B(n_6191),
.Y(n_8624)
);

OAI21x1_ASAP7_75t_L g8625 ( 
.A1(n_7022),
.A2(n_6549),
.B(n_5900),
.Y(n_8625)
);

AND2x2_ASAP7_75t_L g8626 ( 
.A(n_6876),
.B(n_5893),
.Y(n_8626)
);

INVx1_ASAP7_75t_L g8627 ( 
.A(n_7074),
.Y(n_8627)
);

AOI22xp33_ASAP7_75t_L g8628 ( 
.A1(n_6958),
.A2(n_6425),
.B1(n_6520),
.B2(n_6403),
.Y(n_8628)
);

O2A1O1Ixp33_ASAP7_75t_SL g8629 ( 
.A1(n_7274),
.A2(n_7391),
.B(n_6977),
.C(n_7045),
.Y(n_8629)
);

BUFx3_ASAP7_75t_L g8630 ( 
.A(n_6817),
.Y(n_8630)
);

NOR2xp33_ASAP7_75t_L g8631 ( 
.A(n_7056),
.B(n_7069),
.Y(n_8631)
);

NAND2x1p5_ASAP7_75t_L g8632 ( 
.A(n_6908),
.B(n_6972),
.Y(n_8632)
);

NAND3xp33_ASAP7_75t_L g8633 ( 
.A(n_6862),
.B(n_5655),
.C(n_5640),
.Y(n_8633)
);

OAI22xp5_ASAP7_75t_L g8634 ( 
.A1(n_6960),
.A2(n_5601),
.B1(n_5589),
.B2(n_5677),
.Y(n_8634)
);

BUFx2_ASAP7_75t_L g8635 ( 
.A(n_7079),
.Y(n_8635)
);

AO31x2_ASAP7_75t_L g8636 ( 
.A1(n_7566),
.A2(n_6256),
.A3(n_6265),
.B(n_6240),
.Y(n_8636)
);

BUFx3_ASAP7_75t_L g8637 ( 
.A(n_6817),
.Y(n_8637)
);

BUFx2_ASAP7_75t_L g8638 ( 
.A(n_7079),
.Y(n_8638)
);

O2A1O1Ixp33_ASAP7_75t_L g8639 ( 
.A1(n_7060),
.A2(n_6111),
.B(n_6139),
.C(n_6136),
.Y(n_8639)
);

INVx1_ASAP7_75t_L g8640 ( 
.A(n_7074),
.Y(n_8640)
);

OAI21x1_ASAP7_75t_SL g8641 ( 
.A1(n_7395),
.A2(n_5653),
.B(n_5984),
.Y(n_8641)
);

AOI21xp33_ASAP7_75t_L g8642 ( 
.A1(n_7018),
.A2(n_5655),
.B(n_5626),
.Y(n_8642)
);

CKINVDCx5p33_ASAP7_75t_R g8643 ( 
.A(n_7514),
.Y(n_8643)
);

INVx1_ASAP7_75t_L g8644 ( 
.A(n_7082),
.Y(n_8644)
);

AOI21xp5_ASAP7_75t_L g8645 ( 
.A1(n_6782),
.A2(n_6555),
.B(n_6265),
.Y(n_8645)
);

OA21x2_ASAP7_75t_L g8646 ( 
.A1(n_7512),
.A2(n_6265),
.B(n_6256),
.Y(n_8646)
);

INVx2_ASAP7_75t_L g8647 ( 
.A(n_6893),
.Y(n_8647)
);

BUFx12f_ASAP7_75t_L g8648 ( 
.A(n_7186),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_7082),
.Y(n_8649)
);

AND2x2_ASAP7_75t_SL g8650 ( 
.A(n_6980),
.B(n_6392),
.Y(n_8650)
);

INVx2_ASAP7_75t_L g8651 ( 
.A(n_6893),
.Y(n_8651)
);

NOR2x1_ASAP7_75t_SL g8652 ( 
.A(n_6642),
.B(n_5747),
.Y(n_8652)
);

A2O1A1Ixp33_ASAP7_75t_L g8653 ( 
.A1(n_6977),
.A2(n_5790),
.B(n_5820),
.C(n_5677),
.Y(n_8653)
);

AOI21xp5_ASAP7_75t_L g8654 ( 
.A1(n_6716),
.A2(n_6555),
.B(n_6691),
.Y(n_8654)
);

OAI21x1_ASAP7_75t_L g8655 ( 
.A1(n_7022),
.A2(n_6549),
.B(n_6612),
.Y(n_8655)
);

INVx2_ASAP7_75t_L g8656 ( 
.A(n_6893),
.Y(n_8656)
);

OAI21xp5_ASAP7_75t_L g8657 ( 
.A1(n_6875),
.A2(n_5630),
.B(n_5618),
.Y(n_8657)
);

NOR2x1_ASAP7_75t_SL g8658 ( 
.A(n_6642),
.B(n_5747),
.Y(n_8658)
);

AND2x2_ASAP7_75t_L g8659 ( 
.A(n_6876),
.B(n_6877),
.Y(n_8659)
);

HB1xp67_ASAP7_75t_L g8660 ( 
.A(n_7120),
.Y(n_8660)
);

NAND2x1p5_ASAP7_75t_L g8661 ( 
.A(n_6908),
.B(n_5831),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_7082),
.Y(n_8662)
);

AOI22xp5_ASAP7_75t_L g8663 ( 
.A1(n_7146),
.A2(n_5547),
.B1(n_6057),
.B2(n_6136),
.Y(n_8663)
);

NAND2xp5_ASAP7_75t_L g8664 ( 
.A(n_6672),
.B(n_6615),
.Y(n_8664)
);

OAI21x1_ASAP7_75t_L g8665 ( 
.A1(n_7626),
.A2(n_7311),
.B(n_7597),
.Y(n_8665)
);

NOR2xp67_ASAP7_75t_L g8666 ( 
.A(n_7156),
.B(n_5554),
.Y(n_8666)
);

NOR2xp33_ASAP7_75t_L g8667 ( 
.A(n_7056),
.B(n_6139),
.Y(n_8667)
);

INVx2_ASAP7_75t_L g8668 ( 
.A(n_6898),
.Y(n_8668)
);

NOR2xp33_ASAP7_75t_L g8669 ( 
.A(n_7069),
.B(n_6276),
.Y(n_8669)
);

OAI22xp33_ASAP7_75t_L g8670 ( 
.A1(n_6897),
.A2(n_6057),
.B1(n_6606),
.B2(n_5790),
.Y(n_8670)
);

AOI22xp33_ASAP7_75t_L g8671 ( 
.A1(n_6958),
.A2(n_6520),
.B1(n_6551),
.B2(n_6425),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_6898),
.Y(n_8672)
);

A2O1A1Ixp33_ASAP7_75t_L g8673 ( 
.A1(n_7002),
.A2(n_5790),
.B(n_5820),
.C(n_5677),
.Y(n_8673)
);

BUFx6f_ASAP7_75t_L g8674 ( 
.A(n_6908),
.Y(n_8674)
);

INVx2_ASAP7_75t_L g8675 ( 
.A(n_6898),
.Y(n_8675)
);

INVx2_ASAP7_75t_SL g8676 ( 
.A(n_6908),
.Y(n_8676)
);

AO21x2_ASAP7_75t_L g8677 ( 
.A1(n_7578),
.A2(n_6204),
.B(n_6191),
.Y(n_8677)
);

NAND2xp5_ASAP7_75t_L g8678 ( 
.A(n_6675),
.B(n_6615),
.Y(n_8678)
);

CKINVDCx5p33_ASAP7_75t_R g8679 ( 
.A(n_7514),
.Y(n_8679)
);

INVx1_ASAP7_75t_L g8680 ( 
.A(n_7083),
.Y(n_8680)
);

NAND2x1p5_ASAP7_75t_L g8681 ( 
.A(n_6908),
.B(n_5831),
.Y(n_8681)
);

NAND2xp5_ASAP7_75t_SL g8682 ( 
.A(n_6840),
.B(n_5893),
.Y(n_8682)
);

INVx2_ASAP7_75t_L g8683 ( 
.A(n_6898),
.Y(n_8683)
);

NOR2x1_ASAP7_75t_R g8684 ( 
.A(n_7078),
.B(n_6520),
.Y(n_8684)
);

AOI21xp5_ASAP7_75t_L g8685 ( 
.A1(n_6716),
.A2(n_6555),
.B(n_6124),
.Y(n_8685)
);

O2A1O1Ixp33_ASAP7_75t_L g8686 ( 
.A1(n_7432),
.A2(n_6144),
.B(n_6163),
.C(n_6142),
.Y(n_8686)
);

INVx1_ASAP7_75t_L g8687 ( 
.A(n_7083),
.Y(n_8687)
);

OAI21xp5_ASAP7_75t_L g8688 ( 
.A1(n_7432),
.A2(n_5618),
.B(n_5626),
.Y(n_8688)
);

INVx3_ASAP7_75t_L g8689 ( 
.A(n_6663),
.Y(n_8689)
);

O2A1O1Ixp33_ASAP7_75t_SL g8690 ( 
.A1(n_7391),
.A2(n_5636),
.B(n_5856),
.C(n_5592),
.Y(n_8690)
);

AOI22xp33_ASAP7_75t_SL g8691 ( 
.A1(n_7052),
.A2(n_5823),
.B1(n_5858),
.B2(n_5820),
.Y(n_8691)
);

CKINVDCx20_ASAP7_75t_R g8692 ( 
.A(n_6839),
.Y(n_8692)
);

INVx1_ASAP7_75t_L g8693 ( 
.A(n_7083),
.Y(n_8693)
);

INVx1_ASAP7_75t_L g8694 ( 
.A(n_7084),
.Y(n_8694)
);

NAND2xp5_ASAP7_75t_L g8695 ( 
.A(n_6675),
.B(n_6396),
.Y(n_8695)
);

BUFx3_ASAP7_75t_L g8696 ( 
.A(n_7079),
.Y(n_8696)
);

NAND2x1p5_ASAP7_75t_L g8697 ( 
.A(n_6972),
.B(n_7117),
.Y(n_8697)
);

OAI22xp33_ASAP7_75t_L g8698 ( 
.A1(n_6897),
.A2(n_7349),
.B1(n_7373),
.B2(n_7359),
.Y(n_8698)
);

AOI221xp5_ASAP7_75t_L g8699 ( 
.A1(n_7538),
.A2(n_6619),
.B1(n_6163),
.B2(n_6179),
.C(n_6144),
.Y(n_8699)
);

AND2x4_ASAP7_75t_L g8700 ( 
.A(n_7322),
.B(n_5893),
.Y(n_8700)
);

INVxp67_ASAP7_75t_SL g8701 ( 
.A(n_6643),
.Y(n_8701)
);

INVx1_ASAP7_75t_L g8702 ( 
.A(n_7084),
.Y(n_8702)
);

INVx1_ASAP7_75t_SL g8703 ( 
.A(n_7092),
.Y(n_8703)
);

INVx2_ASAP7_75t_L g8704 ( 
.A(n_6900),
.Y(n_8704)
);

INVx1_ASAP7_75t_L g8705 ( 
.A(n_7084),
.Y(n_8705)
);

OAI21xp5_ASAP7_75t_L g8706 ( 
.A1(n_7477),
.A2(n_5618),
.B(n_5606),
.Y(n_8706)
);

OAI21xp5_ASAP7_75t_L g8707 ( 
.A1(n_7477),
.A2(n_5606),
.B(n_5595),
.Y(n_8707)
);

OAI22xp33_ASAP7_75t_L g8708 ( 
.A1(n_7349),
.A2(n_6057),
.B1(n_6606),
.B2(n_5823),
.Y(n_8708)
);

INVx1_ASAP7_75t_L g8709 ( 
.A(n_7095),
.Y(n_8709)
);

NAND2xp5_ASAP7_75t_L g8710 ( 
.A(n_6675),
.B(n_6396),
.Y(n_8710)
);

INVx3_ASAP7_75t_SL g8711 ( 
.A(n_6835),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_7095),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_7095),
.Y(n_8713)
);

NAND2xp5_ASAP7_75t_L g8714 ( 
.A(n_6679),
.B(n_6443),
.Y(n_8714)
);

AND2x2_ASAP7_75t_L g8715 ( 
.A(n_6876),
.B(n_5922),
.Y(n_8715)
);

BUFx2_ASAP7_75t_SL g8716 ( 
.A(n_6823),
.Y(n_8716)
);

AND2x4_ASAP7_75t_L g8717 ( 
.A(n_7322),
.B(n_5922),
.Y(n_8717)
);

INVx2_ASAP7_75t_L g8718 ( 
.A(n_6900),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_7112),
.Y(n_8719)
);

AND2x2_ASAP7_75t_L g8720 ( 
.A(n_6876),
.B(n_5922),
.Y(n_8720)
);

HB1xp67_ASAP7_75t_L g8721 ( 
.A(n_7120),
.Y(n_8721)
);

AND2x4_ASAP7_75t_L g8722 ( 
.A(n_7348),
.B(n_5922),
.Y(n_8722)
);

CKINVDCx5p33_ASAP7_75t_R g8723 ( 
.A(n_7216),
.Y(n_8723)
);

OA21x2_ASAP7_75t_L g8724 ( 
.A1(n_7536),
.A2(n_6210),
.B(n_6208),
.Y(n_8724)
);

AND2x2_ASAP7_75t_L g8725 ( 
.A(n_6877),
.B(n_5922),
.Y(n_8725)
);

INVx2_ASAP7_75t_SL g8726 ( 
.A(n_6972),
.Y(n_8726)
);

NAND2xp5_ASAP7_75t_L g8727 ( 
.A(n_6679),
.B(n_6443),
.Y(n_8727)
);

AO21x2_ASAP7_75t_L g8728 ( 
.A1(n_7578),
.A2(n_6210),
.B(n_6208),
.Y(n_8728)
);

AOI221xp5_ASAP7_75t_L g8729 ( 
.A1(n_7562),
.A2(n_6181),
.B1(n_6195),
.B2(n_6179),
.C(n_6142),
.Y(n_8729)
);

AO21x2_ASAP7_75t_L g8730 ( 
.A1(n_7076),
.A2(n_6234),
.B(n_6212),
.Y(n_8730)
);

AND2x4_ASAP7_75t_L g8731 ( 
.A(n_7348),
.B(n_5922),
.Y(n_8731)
);

BUFx2_ASAP7_75t_L g8732 ( 
.A(n_7079),
.Y(n_8732)
);

INVx2_ASAP7_75t_L g8733 ( 
.A(n_6900),
.Y(n_8733)
);

AO21x2_ASAP7_75t_L g8734 ( 
.A1(n_7076),
.A2(n_6234),
.B(n_6212),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_7112),
.Y(n_8735)
);

OAI21xp5_ASAP7_75t_L g8736 ( 
.A1(n_6840),
.A2(n_5606),
.B(n_5595),
.Y(n_8736)
);

AO31x2_ASAP7_75t_L g8737 ( 
.A1(n_7585),
.A2(n_7204),
.A3(n_7162),
.B(n_7604),
.Y(n_8737)
);

INVx5_ASAP7_75t_L g8738 ( 
.A(n_6663),
.Y(n_8738)
);

AO21x2_ASAP7_75t_L g8739 ( 
.A1(n_7076),
.A2(n_7334),
.B(n_6691),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_7112),
.Y(n_8740)
);

OAI21xp5_ASAP7_75t_L g8741 ( 
.A1(n_7097),
.A2(n_5606),
.B(n_5595),
.Y(n_8741)
);

AO22x2_ASAP7_75t_L g8742 ( 
.A1(n_7625),
.A2(n_5588),
.B1(n_5554),
.B2(n_5783),
.Y(n_8742)
);

INVx3_ASAP7_75t_L g8743 ( 
.A(n_6663),
.Y(n_8743)
);

OAI22xp5_ASAP7_75t_L g8744 ( 
.A1(n_6780),
.A2(n_6859),
.B1(n_7484),
.B2(n_6728),
.Y(n_8744)
);

INVx1_ASAP7_75t_L g8745 ( 
.A(n_7114),
.Y(n_8745)
);

AOI21xp5_ASAP7_75t_L g8746 ( 
.A1(n_6716),
.A2(n_6555),
.B(n_6124),
.Y(n_8746)
);

INVx1_ASAP7_75t_L g8747 ( 
.A(n_7114),
.Y(n_8747)
);

AND2x2_ASAP7_75t_L g8748 ( 
.A(n_6877),
.B(n_5922),
.Y(n_8748)
);

OAI21x1_ASAP7_75t_SL g8749 ( 
.A1(n_7395),
.A2(n_5653),
.B(n_5984),
.Y(n_8749)
);

OAI21x1_ASAP7_75t_L g8750 ( 
.A1(n_6635),
.A2(n_6703),
.B(n_6645),
.Y(n_8750)
);

OA21x2_ASAP7_75t_L g8751 ( 
.A1(n_7536),
.A2(n_6193),
.B(n_5923),
.Y(n_8751)
);

OR2x6_ASAP7_75t_L g8752 ( 
.A(n_7154),
.B(n_5827),
.Y(n_8752)
);

OR2x6_ASAP7_75t_L g8753 ( 
.A(n_7154),
.B(n_5827),
.Y(n_8753)
);

OAI22xp33_ASAP7_75t_L g8754 ( 
.A1(n_7349),
.A2(n_6057),
.B1(n_6606),
.B2(n_5858),
.Y(n_8754)
);

AND2x4_ASAP7_75t_L g8755 ( 
.A(n_7348),
.B(n_5922),
.Y(n_8755)
);

AO21x2_ASAP7_75t_L g8756 ( 
.A1(n_7076),
.A2(n_6269),
.B(n_6260),
.Y(n_8756)
);

AOI21xp5_ASAP7_75t_L g8757 ( 
.A1(n_6691),
.A2(n_6555),
.B(n_6124),
.Y(n_8757)
);

BUFx2_ASAP7_75t_L g8758 ( 
.A(n_7079),
.Y(n_8758)
);

BUFx3_ASAP7_75t_L g8759 ( 
.A(n_7278),
.Y(n_8759)
);

INVx1_ASAP7_75t_L g8760 ( 
.A(n_7114),
.Y(n_8760)
);

INVx4_ASAP7_75t_L g8761 ( 
.A(n_7078),
.Y(n_8761)
);

OAI22xp5_ASAP7_75t_L g8762 ( 
.A1(n_6780),
.A2(n_5601),
.B1(n_5589),
.B2(n_5823),
.Y(n_8762)
);

OR2x2_ASAP7_75t_L g8763 ( 
.A(n_7191),
.B(n_6593),
.Y(n_8763)
);

BUFx2_ASAP7_75t_L g8764 ( 
.A(n_7278),
.Y(n_8764)
);

BUFx2_ASAP7_75t_R g8765 ( 
.A(n_6814),
.Y(n_8765)
);

OAI22xp5_ASAP7_75t_L g8766 ( 
.A1(n_6859),
.A2(n_5601),
.B1(n_5858),
.B2(n_5823),
.Y(n_8766)
);

AOI22xp5_ASAP7_75t_L g8767 ( 
.A1(n_7146),
.A2(n_5547),
.B1(n_6195),
.B2(n_6181),
.Y(n_8767)
);

AOI22xp33_ASAP7_75t_L g8768 ( 
.A1(n_7170),
.A2(n_6728),
.B1(n_7319),
.B2(n_7149),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_L g8769 ( 
.A(n_6679),
.B(n_6488),
.Y(n_8769)
);

AO21x2_ASAP7_75t_L g8770 ( 
.A1(n_7076),
.A2(n_6269),
.B(n_6260),
.Y(n_8770)
);

NOR2xp33_ASAP7_75t_SL g8771 ( 
.A(n_7264),
.B(n_5557),
.Y(n_8771)
);

AOI22xp5_ASAP7_75t_L g8772 ( 
.A1(n_7146),
.A2(n_5547),
.B1(n_6276),
.B2(n_6243),
.Y(n_8772)
);

INVx2_ASAP7_75t_L g8773 ( 
.A(n_6900),
.Y(n_8773)
);

OR2x2_ASAP7_75t_L g8774 ( 
.A(n_7191),
.B(n_6593),
.Y(n_8774)
);

NAND2xp5_ASAP7_75t_L g8775 ( 
.A(n_6777),
.B(n_6488),
.Y(n_8775)
);

NOR2xp33_ASAP7_75t_L g8776 ( 
.A(n_7100),
.B(n_6349),
.Y(n_8776)
);

AOI22xp5_ASAP7_75t_L g8777 ( 
.A1(n_7150),
.A2(n_5547),
.B1(n_6295),
.B2(n_6243),
.Y(n_8777)
);

INVx1_ASAP7_75t_SL g8778 ( 
.A(n_7123),
.Y(n_8778)
);

AND2x2_ASAP7_75t_L g8779 ( 
.A(n_6877),
.B(n_5930),
.Y(n_8779)
);

INVx2_ASAP7_75t_L g8780 ( 
.A(n_6903),
.Y(n_8780)
);

AOI221xp5_ASAP7_75t_L g8781 ( 
.A1(n_7562),
.A2(n_6312),
.B1(n_6319),
.B2(n_6299),
.C(n_6295),
.Y(n_8781)
);

AND2x2_ASAP7_75t_L g8782 ( 
.A(n_6888),
.B(n_5930),
.Y(n_8782)
);

INVx1_ASAP7_75t_L g8783 ( 
.A(n_7119),
.Y(n_8783)
);

AOI22xp5_ASAP7_75t_L g8784 ( 
.A1(n_7150),
.A2(n_5547),
.B1(n_6312),
.B2(n_6299),
.Y(n_8784)
);

AOI21xp5_ASAP7_75t_L g8785 ( 
.A1(n_7677),
.A2(n_6555),
.B(n_6124),
.Y(n_8785)
);

HB1xp67_ASAP7_75t_L g8786 ( 
.A(n_6736),
.Y(n_8786)
);

OA21x2_ASAP7_75t_L g8787 ( 
.A1(n_7210),
.A2(n_6193),
.B(n_5923),
.Y(n_8787)
);

CKINVDCx20_ASAP7_75t_R g8788 ( 
.A(n_6938),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_7119),
.Y(n_8789)
);

AO31x2_ASAP7_75t_L g8790 ( 
.A1(n_7204),
.A2(n_6061),
.A3(n_6062),
.B(n_6042),
.Y(n_8790)
);

OAI22xp5_ASAP7_75t_L g8791 ( 
.A1(n_7484),
.A2(n_5858),
.B1(n_6333),
.B2(n_6319),
.Y(n_8791)
);

OAI21x1_ASAP7_75t_L g8792 ( 
.A1(n_6635),
.A2(n_6703),
.B(n_6645),
.Y(n_8792)
);

AOI22xp33_ASAP7_75t_L g8793 ( 
.A1(n_7170),
.A2(n_6551),
.B1(n_6583),
.B2(n_6606),
.Y(n_8793)
);

AOI21xp5_ASAP7_75t_L g8794 ( 
.A1(n_7677),
.A2(n_6124),
.B(n_5831),
.Y(n_8794)
);

NAND2xp5_ASAP7_75t_L g8795 ( 
.A(n_6777),
.B(n_6598),
.Y(n_8795)
);

HB1xp67_ASAP7_75t_L g8796 ( 
.A(n_6852),
.Y(n_8796)
);

NAND2x1p5_ASAP7_75t_L g8797 ( 
.A(n_6972),
.B(n_5831),
.Y(n_8797)
);

NOR2xp33_ASAP7_75t_SL g8798 ( 
.A(n_7293),
.B(n_5670),
.Y(n_8798)
);

INVx2_ASAP7_75t_L g8799 ( 
.A(n_6903),
.Y(n_8799)
);

AND2x4_ASAP7_75t_L g8800 ( 
.A(n_7348),
.B(n_5930),
.Y(n_8800)
);

NOR2xp67_ASAP7_75t_L g8801 ( 
.A(n_7168),
.B(n_5588),
.Y(n_8801)
);

OAI21x1_ASAP7_75t_SL g8802 ( 
.A1(n_7395),
.A2(n_5653),
.B(n_5984),
.Y(n_8802)
);

NAND2xp5_ASAP7_75t_L g8803 ( 
.A(n_6777),
.B(n_6598),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_7119),
.Y(n_8804)
);

INVx5_ASAP7_75t_L g8805 ( 
.A(n_6670),
.Y(n_8805)
);

CKINVDCx6p67_ASAP7_75t_R g8806 ( 
.A(n_7078),
.Y(n_8806)
);

OAI22xp5_ASAP7_75t_L g8807 ( 
.A1(n_7089),
.A2(n_6333),
.B1(n_6349),
.B2(n_6335),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_7126),
.Y(n_8808)
);

AO31x2_ASAP7_75t_L g8809 ( 
.A1(n_7204),
.A2(n_6073),
.A3(n_6075),
.B(n_6061),
.Y(n_8809)
);

AND2x4_ASAP7_75t_L g8810 ( 
.A(n_7353),
.B(n_5930),
.Y(n_8810)
);

INVx2_ASAP7_75t_L g8811 ( 
.A(n_6903),
.Y(n_8811)
);

NAND2xp5_ASAP7_75t_L g8812 ( 
.A(n_6790),
.B(n_6530),
.Y(n_8812)
);

OA21x2_ASAP7_75t_L g8813 ( 
.A1(n_7210),
.A2(n_6289),
.B(n_6283),
.Y(n_8813)
);

NAND2x1p5_ASAP7_75t_L g8814 ( 
.A(n_6972),
.B(n_6124),
.Y(n_8814)
);

NAND2xp5_ASAP7_75t_L g8815 ( 
.A(n_6790),
.B(n_6831),
.Y(n_8815)
);

AOI21xp5_ASAP7_75t_L g8816 ( 
.A1(n_7097),
.A2(n_6257),
.B(n_6124),
.Y(n_8816)
);

OA21x2_ASAP7_75t_L g8817 ( 
.A1(n_7210),
.A2(n_6289),
.B(n_6283),
.Y(n_8817)
);

CKINVDCx20_ASAP7_75t_R g8818 ( 
.A(n_6938),
.Y(n_8818)
);

INVx1_ASAP7_75t_L g8819 ( 
.A(n_7126),
.Y(n_8819)
);

INVx6_ASAP7_75t_L g8820 ( 
.A(n_7331),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_7126),
.Y(n_8821)
);

BUFx2_ASAP7_75t_R g8822 ( 
.A(n_6867),
.Y(n_8822)
);

AND2x4_ASAP7_75t_L g8823 ( 
.A(n_7353),
.B(n_5930),
.Y(n_8823)
);

INVx2_ASAP7_75t_L g8824 ( 
.A(n_6903),
.Y(n_8824)
);

O2A1O1Ixp33_ASAP7_75t_SL g8825 ( 
.A1(n_7008),
.A2(n_6369),
.B(n_6371),
.C(n_6335),
.Y(n_8825)
);

AOI21x1_ASAP7_75t_L g8826 ( 
.A1(n_7579),
.A2(n_5747),
.B(n_5799),
.Y(n_8826)
);

OAI21xp5_ASAP7_75t_L g8827 ( 
.A1(n_7113),
.A2(n_5606),
.B(n_5595),
.Y(n_8827)
);

INVx1_ASAP7_75t_L g8828 ( 
.A(n_7138),
.Y(n_8828)
);

AND2x2_ASAP7_75t_L g8829 ( 
.A(n_6888),
.B(n_5930),
.Y(n_8829)
);

AOI22xp5_ASAP7_75t_L g8830 ( 
.A1(n_7150),
.A2(n_5547),
.B1(n_6371),
.B2(n_6369),
.Y(n_8830)
);

INVx1_ASAP7_75t_L g8831 ( 
.A(n_7138),
.Y(n_8831)
);

INVx1_ASAP7_75t_SL g8832 ( 
.A(n_7123),
.Y(n_8832)
);

NAND2xp33_ASAP7_75t_L g8833 ( 
.A(n_6726),
.B(n_4865),
.Y(n_8833)
);

OAI22xp5_ASAP7_75t_SL g8834 ( 
.A1(n_7008),
.A2(n_7045),
.B1(n_6987),
.B2(n_7078),
.Y(n_8834)
);

AND2x4_ASAP7_75t_L g8835 ( 
.A(n_7353),
.B(n_5930),
.Y(n_8835)
);

OAI22xp33_ASAP7_75t_L g8836 ( 
.A1(n_7373),
.A2(n_6388),
.B1(n_6399),
.B2(n_6389),
.Y(n_8836)
);

INVx4_ASAP7_75t_L g8837 ( 
.A(n_7259),
.Y(n_8837)
);

OAI21xp5_ASAP7_75t_L g8838 ( 
.A1(n_7113),
.A2(n_5595),
.B(n_5550),
.Y(n_8838)
);

AOI22xp5_ASAP7_75t_L g8839 ( 
.A1(n_7162),
.A2(n_5547),
.B1(n_6389),
.B2(n_6388),
.Y(n_8839)
);

AOI221xp5_ASAP7_75t_L g8840 ( 
.A1(n_6874),
.A2(n_6408),
.B1(n_6413),
.B2(n_6405),
.C(n_6399),
.Y(n_8840)
);

AND2x6_ASAP7_75t_L g8841 ( 
.A(n_6632),
.B(n_5230),
.Y(n_8841)
);

CKINVDCx5p33_ASAP7_75t_R g8842 ( 
.A(n_7216),
.Y(n_8842)
);

A2O1A1Ixp33_ASAP7_75t_L g8843 ( 
.A1(n_7002),
.A2(n_6249),
.B(n_6532),
.C(n_6241),
.Y(n_8843)
);

INVx3_ASAP7_75t_L g8844 ( 
.A(n_6670),
.Y(n_8844)
);

OR2x2_ASAP7_75t_L g8845 ( 
.A(n_7201),
.B(n_7215),
.Y(n_8845)
);

CKINVDCx5p33_ASAP7_75t_R g8846 ( 
.A(n_7246),
.Y(n_8846)
);

CKINVDCx16_ASAP7_75t_R g8847 ( 
.A(n_7259),
.Y(n_8847)
);

INVx1_ASAP7_75t_L g8848 ( 
.A(n_7138),
.Y(n_8848)
);

AND2x2_ASAP7_75t_L g8849 ( 
.A(n_6888),
.B(n_5930),
.Y(n_8849)
);

AND2x2_ASAP7_75t_L g8850 ( 
.A(n_6888),
.B(n_5949),
.Y(n_8850)
);

BUFx6f_ASAP7_75t_L g8851 ( 
.A(n_6972),
.Y(n_8851)
);

OR2x6_ASAP7_75t_L g8852 ( 
.A(n_7483),
.B(n_5827),
.Y(n_8852)
);

INVx1_ASAP7_75t_L g8853 ( 
.A(n_7163),
.Y(n_8853)
);

CKINVDCx20_ASAP7_75t_R g8854 ( 
.A(n_7678),
.Y(n_8854)
);

INVx1_ASAP7_75t_L g8855 ( 
.A(n_7163),
.Y(n_8855)
);

AND2x2_ASAP7_75t_L g8856 ( 
.A(n_6901),
.B(n_5949),
.Y(n_8856)
);

AOI22xp33_ASAP7_75t_L g8857 ( 
.A1(n_7170),
.A2(n_6551),
.B1(n_6583),
.B2(n_5836),
.Y(n_8857)
);

INVx2_ASAP7_75t_L g8858 ( 
.A(n_6926),
.Y(n_8858)
);

BUFx3_ASAP7_75t_L g8859 ( 
.A(n_7278),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_7163),
.Y(n_8860)
);

INVx2_ASAP7_75t_L g8861 ( 
.A(n_6926),
.Y(n_8861)
);

BUFx2_ASAP7_75t_L g8862 ( 
.A(n_7278),
.Y(n_8862)
);

CKINVDCx5p33_ASAP7_75t_R g8863 ( 
.A(n_7246),
.Y(n_8863)
);

AND2x2_ASAP7_75t_L g8864 ( 
.A(n_6901),
.B(n_6918),
.Y(n_8864)
);

AOI21xp5_ASAP7_75t_L g8865 ( 
.A1(n_6655),
.A2(n_6257),
.B(n_6124),
.Y(n_8865)
);

AOI222xp33_ASAP7_75t_L g8866 ( 
.A1(n_7315),
.A2(n_6583),
.B1(n_6405),
.B2(n_6413),
.C1(n_6438),
.C2(n_6415),
.Y(n_8866)
);

BUFx6f_ASAP7_75t_L g8867 ( 
.A(n_6972),
.Y(n_8867)
);

AO21x2_ASAP7_75t_L g8868 ( 
.A1(n_7076),
.A2(n_7334),
.B(n_7598),
.Y(n_8868)
);

OAI22xp5_ASAP7_75t_L g8869 ( 
.A1(n_7089),
.A2(n_6415),
.B1(n_6438),
.B2(n_6408),
.Y(n_8869)
);

AND2x6_ASAP7_75t_L g8870 ( 
.A(n_6632),
.B(n_5268),
.Y(n_8870)
);

INVx1_ASAP7_75t_L g8871 ( 
.A(n_7179),
.Y(n_8871)
);

AO31x2_ASAP7_75t_L g8872 ( 
.A1(n_7162),
.A2(n_7604),
.A3(n_7341),
.B(n_7340),
.Y(n_8872)
);

NOR2x1_ASAP7_75t_SL g8873 ( 
.A(n_6642),
.B(n_5949),
.Y(n_8873)
);

AND2x2_ASAP7_75t_L g8874 ( 
.A(n_6901),
.B(n_5949),
.Y(n_8874)
);

CKINVDCx20_ASAP7_75t_R g8875 ( 
.A(n_7678),
.Y(n_8875)
);

NOR2xp33_ASAP7_75t_L g8876 ( 
.A(n_7100),
.B(n_6452),
.Y(n_8876)
);

HB1xp67_ASAP7_75t_L g8877 ( 
.A(n_6852),
.Y(n_8877)
);

A2O1A1Ixp33_ASAP7_75t_L g8878 ( 
.A1(n_7130),
.A2(n_6249),
.B(n_6532),
.C(n_6241),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_7179),
.Y(n_8879)
);

AOI22xp33_ASAP7_75t_L g8880 ( 
.A1(n_7319),
.A2(n_5550),
.B1(n_5547),
.B2(n_5794),
.Y(n_8880)
);

INVx2_ASAP7_75t_L g8881 ( 
.A(n_6926),
.Y(n_8881)
);

INVx2_ASAP7_75t_L g8882 ( 
.A(n_6926),
.Y(n_8882)
);

INVx1_ASAP7_75t_L g8883 ( 
.A(n_7179),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_7188),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_7188),
.Y(n_8885)
);

INVx1_ASAP7_75t_L g8886 ( 
.A(n_7188),
.Y(n_8886)
);

INVxp67_ASAP7_75t_L g8887 ( 
.A(n_6831),
.Y(n_8887)
);

NOR2xp33_ASAP7_75t_R g8888 ( 
.A(n_6867),
.B(n_5670),
.Y(n_8888)
);

INVx2_ASAP7_75t_L g8889 ( 
.A(n_6930),
.Y(n_8889)
);

INVx1_ASAP7_75t_L g8890 ( 
.A(n_7189),
.Y(n_8890)
);

CKINVDCx5p33_ASAP7_75t_R g8891 ( 
.A(n_7252),
.Y(n_8891)
);

A2O1A1Ixp33_ASAP7_75t_L g8892 ( 
.A1(n_7130),
.A2(n_6249),
.B(n_6532),
.C(n_6241),
.Y(n_8892)
);

NOR2xp33_ASAP7_75t_L g8893 ( 
.A(n_7582),
.B(n_6516),
.Y(n_8893)
);

OAI21x1_ASAP7_75t_SL g8894 ( 
.A1(n_7131),
.A2(n_7444),
.B(n_7125),
.Y(n_8894)
);

BUFx2_ASAP7_75t_L g8895 ( 
.A(n_7278),
.Y(n_8895)
);

OA21x2_ASAP7_75t_L g8896 ( 
.A1(n_7509),
.A2(n_6300),
.B(n_6291),
.Y(n_8896)
);

CKINVDCx5p33_ASAP7_75t_R g8897 ( 
.A(n_7252),
.Y(n_8897)
);

CKINVDCx6p67_ASAP7_75t_R g8898 ( 
.A(n_7259),
.Y(n_8898)
);

OAI22xp33_ASAP7_75t_L g8899 ( 
.A1(n_7373),
.A2(n_6460),
.B1(n_6463),
.B2(n_6452),
.Y(n_8899)
);

INVx1_ASAP7_75t_L g8900 ( 
.A(n_7189),
.Y(n_8900)
);

NAND2xp5_ASAP7_75t_L g8901 ( 
.A(n_6790),
.B(n_6530),
.Y(n_8901)
);

INVx1_ASAP7_75t_L g8902 ( 
.A(n_7189),
.Y(n_8902)
);

INVx2_ASAP7_75t_R g8903 ( 
.A(n_6972),
.Y(n_8903)
);

OAI22xp5_ASAP7_75t_L g8904 ( 
.A1(n_7315),
.A2(n_6463),
.B1(n_6477),
.B2(n_6460),
.Y(n_8904)
);

INVx2_ASAP7_75t_L g8905 ( 
.A(n_6930),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_6831),
.B(n_6572),
.Y(n_8906)
);

AOI21xp5_ASAP7_75t_L g8907 ( 
.A1(n_6655),
.A2(n_6257),
.B(n_6124),
.Y(n_8907)
);

INVx1_ASAP7_75t_L g8908 ( 
.A(n_7195),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_7195),
.Y(n_8909)
);

INVx2_ASAP7_75t_L g8910 ( 
.A(n_6930),
.Y(n_8910)
);

OAI22xp5_ASAP7_75t_L g8911 ( 
.A1(n_6883),
.A2(n_6483),
.B1(n_6487),
.B2(n_6477),
.Y(n_8911)
);

CKINVDCx6p67_ASAP7_75t_R g8912 ( 
.A(n_7259),
.Y(n_8912)
);

INVx2_ASAP7_75t_SL g8913 ( 
.A(n_6972),
.Y(n_8913)
);

INVx2_ASAP7_75t_L g8914 ( 
.A(n_6930),
.Y(n_8914)
);

AND2x2_ASAP7_75t_L g8915 ( 
.A(n_6901),
.B(n_5949),
.Y(n_8915)
);

AND2x2_ASAP7_75t_L g8916 ( 
.A(n_6918),
.B(n_5949),
.Y(n_8916)
);

NAND2xp5_ASAP7_75t_L g8917 ( 
.A(n_6838),
.B(n_6572),
.Y(n_8917)
);

NOR2x1_ASAP7_75t_SL g8918 ( 
.A(n_7458),
.B(n_5949),
.Y(n_8918)
);

INVx3_ASAP7_75t_SL g8919 ( 
.A(n_6835),
.Y(n_8919)
);

INVx2_ASAP7_75t_L g8920 ( 
.A(n_6935),
.Y(n_8920)
);

OAI21xp5_ASAP7_75t_L g8921 ( 
.A1(n_6753),
.A2(n_5550),
.B(n_5794),
.Y(n_8921)
);

OR2x6_ASAP7_75t_L g8922 ( 
.A(n_7483),
.B(n_5827),
.Y(n_8922)
);

OA21x2_ASAP7_75t_L g8923 ( 
.A1(n_7509),
.A2(n_6300),
.B(n_6291),
.Y(n_8923)
);

INVx2_ASAP7_75t_L g8924 ( 
.A(n_6935),
.Y(n_8924)
);

OR2x2_ASAP7_75t_L g8925 ( 
.A(n_7201),
.B(n_6593),
.Y(n_8925)
);

CKINVDCx5p33_ASAP7_75t_R g8926 ( 
.A(n_7436),
.Y(n_8926)
);

NOR2xp33_ASAP7_75t_L g8927 ( 
.A(n_7582),
.B(n_7606),
.Y(n_8927)
);

OAI22xp5_ASAP7_75t_L g8928 ( 
.A1(n_6883),
.A2(n_6487),
.B1(n_6489),
.B2(n_6483),
.Y(n_8928)
);

OAI222xp33_ASAP7_75t_L g8929 ( 
.A1(n_7052),
.A2(n_6489),
.B1(n_6492),
.B2(n_6565),
.C1(n_6554),
.C2(n_6516),
.Y(n_8929)
);

INVx2_ASAP7_75t_L g8930 ( 
.A(n_6935),
.Y(n_8930)
);

OR2x6_ASAP7_75t_L g8931 ( 
.A(n_7483),
.B(n_5830),
.Y(n_8931)
);

INVx1_ASAP7_75t_L g8932 ( 
.A(n_7195),
.Y(n_8932)
);

BUFx3_ASAP7_75t_L g8933 ( 
.A(n_7278),
.Y(n_8933)
);

AOI22xp33_ASAP7_75t_L g8934 ( 
.A1(n_7149),
.A2(n_5550),
.B1(n_5813),
.B2(n_5726),
.Y(n_8934)
);

NAND2x1p5_ASAP7_75t_L g8935 ( 
.A(n_6972),
.B(n_6257),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_7197),
.Y(n_8936)
);

A2O1A1Ixp33_ASAP7_75t_L g8937 ( 
.A1(n_7683),
.A2(n_6249),
.B(n_6532),
.C(n_6241),
.Y(n_8937)
);

NOR2xp33_ASAP7_75t_L g8938 ( 
.A(n_7606),
.B(n_6492),
.Y(n_8938)
);

BUFx6f_ASAP7_75t_L g8939 ( 
.A(n_7117),
.Y(n_8939)
);

BUFx3_ASAP7_75t_L g8940 ( 
.A(n_7278),
.Y(n_8940)
);

AOI21xp5_ASAP7_75t_L g8941 ( 
.A1(n_6669),
.A2(n_6273),
.B(n_6257),
.Y(n_8941)
);

AOI21xp5_ASAP7_75t_L g8942 ( 
.A1(n_6669),
.A2(n_7249),
.B(n_7180),
.Y(n_8942)
);

INVx3_ASAP7_75t_L g8943 ( 
.A(n_6670),
.Y(n_8943)
);

AOI22xp33_ASAP7_75t_SL g8944 ( 
.A1(n_7052),
.A2(n_5670),
.B1(n_6024),
.B2(n_5834),
.Y(n_8944)
);

NOR2xp67_ASAP7_75t_L g8945 ( 
.A(n_7168),
.B(n_5783),
.Y(n_8945)
);

INVx2_ASAP7_75t_L g8946 ( 
.A(n_6935),
.Y(n_8946)
);

OAI22xp5_ASAP7_75t_L g8947 ( 
.A1(n_6921),
.A2(n_6565),
.B1(n_6566),
.B2(n_6554),
.Y(n_8947)
);

BUFx6f_ASAP7_75t_L g8948 ( 
.A(n_7117),
.Y(n_8948)
);

INVx1_ASAP7_75t_L g8949 ( 
.A(n_7197),
.Y(n_8949)
);

AND2x4_ASAP7_75t_L g8950 ( 
.A(n_7353),
.B(n_5949),
.Y(n_8950)
);

INVx1_ASAP7_75t_L g8951 ( 
.A(n_7197),
.Y(n_8951)
);

OA21x2_ASAP7_75t_L g8952 ( 
.A1(n_7520),
.A2(n_6302),
.B(n_6301),
.Y(n_8952)
);

INVx5_ASAP7_75t_L g8953 ( 
.A(n_6670),
.Y(n_8953)
);

OA21x2_ASAP7_75t_L g8954 ( 
.A1(n_7520),
.A2(n_6302),
.B(n_6301),
.Y(n_8954)
);

AND2x2_ASAP7_75t_L g8955 ( 
.A(n_6918),
.B(n_5963),
.Y(n_8955)
);

INVx2_ASAP7_75t_L g8956 ( 
.A(n_6940),
.Y(n_8956)
);

CKINVDCx16_ASAP7_75t_R g8957 ( 
.A(n_7346),
.Y(n_8957)
);

NOR2xp33_ASAP7_75t_L g8958 ( 
.A(n_6729),
.B(n_6577),
.Y(n_8958)
);

OR2x6_ASAP7_75t_L g8959 ( 
.A(n_7483),
.B(n_7226),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_7202),
.Y(n_8960)
);

OA21x2_ASAP7_75t_L g8961 ( 
.A1(n_7633),
.A2(n_6698),
.B(n_6685),
.Y(n_8961)
);

OR2x6_ASAP7_75t_L g8962 ( 
.A(n_7483),
.B(n_7226),
.Y(n_8962)
);

INVx2_ASAP7_75t_SL g8963 ( 
.A(n_7117),
.Y(n_8963)
);

AO21x2_ASAP7_75t_L g8964 ( 
.A1(n_7334),
.A2(n_6330),
.B(n_6316),
.Y(n_8964)
);

CKINVDCx5p33_ASAP7_75t_R g8965 ( 
.A(n_7436),
.Y(n_8965)
);

OAI22xp5_ASAP7_75t_L g8966 ( 
.A1(n_6921),
.A2(n_6577),
.B1(n_6566),
.B2(n_5726),
.Y(n_8966)
);

INVx2_ASAP7_75t_L g8967 ( 
.A(n_6940),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_7202),
.Y(n_8968)
);

AOI22xp33_ASAP7_75t_L g8969 ( 
.A1(n_7006),
.A2(n_5550),
.B1(n_5813),
.B2(n_5731),
.Y(n_8969)
);

AND2x2_ASAP7_75t_L g8970 ( 
.A(n_6918),
.B(n_5963),
.Y(n_8970)
);

INVx1_ASAP7_75t_L g8971 ( 
.A(n_7202),
.Y(n_8971)
);

O2A1O1Ixp33_ASAP7_75t_L g8972 ( 
.A1(n_7402),
.A2(n_7148),
.B(n_7018),
.C(n_7683),
.Y(n_8972)
);

NAND2x1p5_ASAP7_75t_L g8973 ( 
.A(n_7117),
.B(n_6257),
.Y(n_8973)
);

BUFx12f_ASAP7_75t_L g8974 ( 
.A(n_7186),
.Y(n_8974)
);

AND2x6_ASAP7_75t_L g8975 ( 
.A(n_6632),
.B(n_5314),
.Y(n_8975)
);

CKINVDCx11_ASAP7_75t_R g8976 ( 
.A(n_7346),
.Y(n_8976)
);

NOR2xp33_ASAP7_75t_SL g8977 ( 
.A(n_7293),
.B(n_5670),
.Y(n_8977)
);

AND2x4_ASAP7_75t_L g8978 ( 
.A(n_7384),
.B(n_5963),
.Y(n_8978)
);

NOR2x1_ASAP7_75t_SL g8979 ( 
.A(n_7458),
.B(n_5963),
.Y(n_8979)
);

OAI21xp5_ASAP7_75t_L g8980 ( 
.A1(n_6753),
.A2(n_5731),
.B(n_5725),
.Y(n_8980)
);

BUFx12f_ASAP7_75t_L g8981 ( 
.A(n_7355),
.Y(n_8981)
);

INVx2_ASAP7_75t_L g8982 ( 
.A(n_6940),
.Y(n_8982)
);

NOR2x1_ASAP7_75t_L g8983 ( 
.A(n_7449),
.B(n_6562),
.Y(n_8983)
);

OAI222xp33_ASAP7_75t_L g8984 ( 
.A1(n_7279),
.A2(n_5867),
.B1(n_5865),
.B2(n_5763),
.C1(n_5750),
.C2(n_5764),
.Y(n_8984)
);

OAI21x1_ASAP7_75t_L g8985 ( 
.A1(n_6766),
.A2(n_6849),
.B(n_6846),
.Y(n_8985)
);

O2A1O1Ixp33_ASAP7_75t_L g8986 ( 
.A1(n_7402),
.A2(n_5750),
.B(n_5762),
.C(n_5725),
.Y(n_8986)
);

INVx1_ASAP7_75t_L g8987 ( 
.A(n_7203),
.Y(n_8987)
);

INVx6_ASAP7_75t_L g8988 ( 
.A(n_7331),
.Y(n_8988)
);

NOR3xp33_ASAP7_75t_SL g8989 ( 
.A(n_6991),
.B(n_5763),
.C(n_5762),
.Y(n_8989)
);

OAI21x1_ASAP7_75t_L g8990 ( 
.A1(n_6766),
.A2(n_6849),
.B(n_6846),
.Y(n_8990)
);

NAND2x1_ASAP7_75t_L g8991 ( 
.A(n_7278),
.B(n_5963),
.Y(n_8991)
);

CKINVDCx16_ASAP7_75t_R g8992 ( 
.A(n_7346),
.Y(n_8992)
);

OAI22xp5_ASAP7_75t_L g8993 ( 
.A1(n_6954),
.A2(n_5764),
.B1(n_5865),
.B2(n_6241),
.Y(n_8993)
);

OAI22xp5_ASAP7_75t_L g8994 ( 
.A1(n_6954),
.A2(n_6249),
.B1(n_6576),
.B2(n_6532),
.Y(n_8994)
);

INVx1_ASAP7_75t_SL g8995 ( 
.A(n_7123),
.Y(n_8995)
);

INVxp67_ASAP7_75t_L g8996 ( 
.A(n_6838),
.Y(n_8996)
);

A2O1A1Ixp33_ASAP7_75t_L g8997 ( 
.A1(n_7352),
.A2(n_6604),
.B(n_6576),
.C(n_6014),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_7203),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_7203),
.Y(n_8999)
);

A2O1A1Ixp33_ASAP7_75t_L g9000 ( 
.A1(n_7352),
.A2(n_6604),
.B(n_6576),
.C(n_6014),
.Y(n_9000)
);

OA21x2_ASAP7_75t_L g9001 ( 
.A1(n_6685),
.A2(n_6330),
.B(n_6316),
.Y(n_9001)
);

OAI222xp33_ASAP7_75t_L g9002 ( 
.A1(n_7279),
.A2(n_7148),
.B1(n_7194),
.B2(n_6753),
.C1(n_7229),
.C2(n_6660),
.Y(n_9002)
);

AOI21xp5_ASAP7_75t_L g9003 ( 
.A1(n_7180),
.A2(n_6273),
.B(n_6257),
.Y(n_9003)
);

INVx3_ASAP7_75t_L g9004 ( 
.A(n_6670),
.Y(n_9004)
);

INVx1_ASAP7_75t_L g9005 ( 
.A(n_7211),
.Y(n_9005)
);

NAND2x1p5_ASAP7_75t_L g9006 ( 
.A(n_7117),
.B(n_6257),
.Y(n_9006)
);

AND2x2_ASAP7_75t_L g9007 ( 
.A(n_6964),
.B(n_5963),
.Y(n_9007)
);

BUFx6f_ASAP7_75t_L g9008 ( 
.A(n_7117),
.Y(n_9008)
);

BUFx12f_ASAP7_75t_L g9009 ( 
.A(n_7355),
.Y(n_9009)
);

BUFx2_ASAP7_75t_SL g9010 ( 
.A(n_6823),
.Y(n_9010)
);

NAND2xp5_ASAP7_75t_L g9011 ( 
.A(n_6838),
.B(n_6586),
.Y(n_9011)
);

NAND2xp5_ASAP7_75t_L g9012 ( 
.A(n_6863),
.B(n_6586),
.Y(n_9012)
);

INVx1_ASAP7_75t_L g9013 ( 
.A(n_7211),
.Y(n_9013)
);

INVx2_ASAP7_75t_L g9014 ( 
.A(n_6940),
.Y(n_9014)
);

NAND2xp5_ASAP7_75t_L g9015 ( 
.A(n_6863),
.B(n_6605),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_7211),
.Y(n_9016)
);

NAND2x1_ASAP7_75t_L g9017 ( 
.A(n_7278),
.B(n_5963),
.Y(n_9017)
);

AND2x4_ASAP7_75t_L g9018 ( 
.A(n_7384),
.B(n_5963),
.Y(n_9018)
);

AO21x2_ASAP7_75t_L g9019 ( 
.A1(n_7334),
.A2(n_6338),
.B(n_6331),
.Y(n_9019)
);

OAI21xp5_ASAP7_75t_L g9020 ( 
.A1(n_6660),
.A2(n_5857),
.B(n_5867),
.Y(n_9020)
);

INVx1_ASAP7_75t_L g9021 ( 
.A(n_7217),
.Y(n_9021)
);

AOI22xp5_ASAP7_75t_L g9022 ( 
.A1(n_7093),
.A2(n_5739),
.B1(n_5742),
.B2(n_5719),
.Y(n_9022)
);

INVx1_ASAP7_75t_L g9023 ( 
.A(n_7217),
.Y(n_9023)
);

BUFx3_ASAP7_75t_L g9024 ( 
.A(n_7278),
.Y(n_9024)
);

AOI221xp5_ASAP7_75t_L g9025 ( 
.A1(n_6874),
.A2(n_5857),
.B1(n_6605),
.B2(n_5716),
.C(n_5728),
.Y(n_9025)
);

AO21x2_ASAP7_75t_L g9026 ( 
.A1(n_7334),
.A2(n_6338),
.B(n_6331),
.Y(n_9026)
);

AND2x4_ASAP7_75t_L g9027 ( 
.A(n_7384),
.B(n_6014),
.Y(n_9027)
);

AOI222xp33_ASAP7_75t_L g9028 ( 
.A1(n_7281),
.A2(n_5670),
.B1(n_6024),
.B2(n_5834),
.C1(n_6604),
.C2(n_6576),
.Y(n_9028)
);

AOI22xp33_ASAP7_75t_L g9029 ( 
.A1(n_7006),
.A2(n_5867),
.B1(n_5809),
.B2(n_5808),
.Y(n_9029)
);

INVx2_ASAP7_75t_L g9030 ( 
.A(n_6945),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_7217),
.Y(n_9031)
);

AOI22xp33_ASAP7_75t_L g9032 ( 
.A1(n_8009),
.A2(n_6980),
.B1(n_7625),
.B2(n_7616),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_7708),
.Y(n_9033)
);

AND2x2_ASAP7_75t_L g9034 ( 
.A(n_8031),
.B(n_6685),
.Y(n_9034)
);

AO21x1_ASAP7_75t_L g9035 ( 
.A1(n_7742),
.A2(n_7131),
.B(n_7024),
.Y(n_9035)
);

HB1xp67_ASAP7_75t_L g9036 ( 
.A(n_8796),
.Y(n_9036)
);

CKINVDCx11_ASAP7_75t_R g9037 ( 
.A(n_8237),
.Y(n_9037)
);

INVx2_ASAP7_75t_SL g9038 ( 
.A(n_7771),
.Y(n_9038)
);

AOI22xp33_ASAP7_75t_L g9039 ( 
.A1(n_8009),
.A2(n_7844),
.B1(n_7742),
.B2(n_7806),
.Y(n_9039)
);

INVx2_ASAP7_75t_L g9040 ( 
.A(n_8724),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_7708),
.Y(n_9041)
);

INVx4_ASAP7_75t_L g9042 ( 
.A(n_7888),
.Y(n_9042)
);

AND2x2_ASAP7_75t_L g9043 ( 
.A(n_8031),
.B(n_6698),
.Y(n_9043)
);

HB1xp67_ASAP7_75t_L g9044 ( 
.A(n_8796),
.Y(n_9044)
);

NOR2xp33_ASAP7_75t_L g9045 ( 
.A(n_8073),
.B(n_7153),
.Y(n_9045)
);

INVx4_ASAP7_75t_L g9046 ( 
.A(n_7888),
.Y(n_9046)
);

HB1xp67_ASAP7_75t_L g9047 ( 
.A(n_8877),
.Y(n_9047)
);

NAND2x1p5_ASAP7_75t_L g9048 ( 
.A(n_8983),
.B(n_7449),
.Y(n_9048)
);

AND2x2_ASAP7_75t_L g9049 ( 
.A(n_8031),
.B(n_6698),
.Y(n_9049)
);

INVx2_ASAP7_75t_L g9050 ( 
.A(n_8724),
.Y(n_9050)
);

AOI22xp33_ASAP7_75t_L g9051 ( 
.A1(n_7844),
.A2(n_6980),
.B1(n_7625),
.B2(n_7616),
.Y(n_9051)
);

INVx1_ASAP7_75t_L g9052 ( 
.A(n_7709),
.Y(n_9052)
);

OAI21x1_ASAP7_75t_L g9053 ( 
.A1(n_7873),
.A2(n_7561),
.B(n_7449),
.Y(n_9053)
);

INVx2_ASAP7_75t_L g9054 ( 
.A(n_8724),
.Y(n_9054)
);

INVx4_ASAP7_75t_L g9055 ( 
.A(n_7888),
.Y(n_9055)
);

AOI22xp33_ASAP7_75t_SL g9056 ( 
.A1(n_7806),
.A2(n_6980),
.B1(n_7616),
.B2(n_7093),
.Y(n_9056)
);

CKINVDCx6p67_ASAP7_75t_R g9057 ( 
.A(n_7953),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_7709),
.Y(n_9058)
);

INVx1_ASAP7_75t_L g9059 ( 
.A(n_7716),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_7716),
.Y(n_9060)
);

INVx1_ASAP7_75t_L g9061 ( 
.A(n_7721),
.Y(n_9061)
);

AOI22xp33_ASAP7_75t_L g9062 ( 
.A1(n_7886),
.A2(n_6980),
.B1(n_7625),
.B2(n_7183),
.Y(n_9062)
);

INVx2_ASAP7_75t_L g9063 ( 
.A(n_8724),
.Y(n_9063)
);

INVx1_ASAP7_75t_L g9064 ( 
.A(n_7721),
.Y(n_9064)
);

INVx1_ASAP7_75t_L g9065 ( 
.A(n_7723),
.Y(n_9065)
);

AND2x4_ASAP7_75t_L g9066 ( 
.A(n_8696),
.B(n_8759),
.Y(n_9066)
);

INVxp33_ASAP7_75t_L g9067 ( 
.A(n_8123),
.Y(n_9067)
);

HB1xp67_ASAP7_75t_L g9068 ( 
.A(n_8877),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_7723),
.Y(n_9069)
);

AOI21x1_ASAP7_75t_L g9070 ( 
.A1(n_7998),
.A2(n_7486),
.B(n_7247),
.Y(n_9070)
);

INVx1_ASAP7_75t_L g9071 ( 
.A(n_7725),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_7725),
.Y(n_9072)
);

AOI22xp33_ASAP7_75t_L g9073 ( 
.A1(n_7886),
.A2(n_7183),
.B1(n_7185),
.B2(n_7367),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_7727),
.Y(n_9074)
);

INVx1_ASAP7_75t_L g9075 ( 
.A(n_7727),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_7729),
.Y(n_9076)
);

AOI22xp33_ASAP7_75t_L g9077 ( 
.A1(n_7985),
.A2(n_7185),
.B1(n_7367),
.B2(n_7358),
.Y(n_9077)
);

INVx2_ASAP7_75t_L g9078 ( 
.A(n_8724),
.Y(n_9078)
);

INVx2_ASAP7_75t_L g9079 ( 
.A(n_8724),
.Y(n_9079)
);

INVx4_ASAP7_75t_L g9080 ( 
.A(n_8648),
.Y(n_9080)
);

INVx3_ASAP7_75t_L g9081 ( 
.A(n_7771),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_7729),
.Y(n_9082)
);

INVx2_ASAP7_75t_L g9083 ( 
.A(n_9001),
.Y(n_9083)
);

INVx2_ASAP7_75t_L g9084 ( 
.A(n_9001),
.Y(n_9084)
);

INVx1_ASAP7_75t_L g9085 ( 
.A(n_7735),
.Y(n_9085)
);

NOR2xp33_ASAP7_75t_L g9086 ( 
.A(n_8073),
.B(n_8847),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_7735),
.Y(n_9087)
);

HB1xp67_ASAP7_75t_L g9088 ( 
.A(n_8786),
.Y(n_9088)
);

INVx2_ASAP7_75t_L g9089 ( 
.A(n_9001),
.Y(n_9089)
);

HB1xp67_ASAP7_75t_L g9090 ( 
.A(n_8786),
.Y(n_9090)
);

AOI22xp33_ASAP7_75t_L g9091 ( 
.A1(n_7985),
.A2(n_7358),
.B1(n_7443),
.B2(n_7379),
.Y(n_9091)
);

AOI22xp33_ASAP7_75t_L g9092 ( 
.A1(n_7803),
.A2(n_7379),
.B1(n_7443),
.B2(n_7238),
.Y(n_9092)
);

INVx1_ASAP7_75t_L g9093 ( 
.A(n_7740),
.Y(n_9093)
);

OAI21x1_ASAP7_75t_L g9094 ( 
.A1(n_9003),
.A2(n_7565),
.B(n_7561),
.Y(n_9094)
);

INVx3_ASAP7_75t_L g9095 ( 
.A(n_7771),
.Y(n_9095)
);

INVx2_ASAP7_75t_L g9096 ( 
.A(n_9001),
.Y(n_9096)
);

NAND2x1p5_ASAP7_75t_L g9097 ( 
.A(n_8983),
.B(n_7561),
.Y(n_9097)
);

BUFx6f_ASAP7_75t_L g9098 ( 
.A(n_8648),
.Y(n_9098)
);

CKINVDCx11_ASAP7_75t_R g9099 ( 
.A(n_8237),
.Y(n_9099)
);

BUFx6f_ASAP7_75t_L g9100 ( 
.A(n_8648),
.Y(n_9100)
);

INVx1_ASAP7_75t_L g9101 ( 
.A(n_7740),
.Y(n_9101)
);

HB1xp67_ASAP7_75t_L g9102 ( 
.A(n_7758),
.Y(n_9102)
);

AOI22xp33_ASAP7_75t_L g9103 ( 
.A1(n_7803),
.A2(n_7238),
.B1(n_7093),
.B2(n_7194),
.Y(n_9103)
);

OAI21xp5_ASAP7_75t_L g9104 ( 
.A1(n_7756),
.A2(n_7194),
.B(n_7229),
.Y(n_9104)
);

BUFx10_ASAP7_75t_L g9105 ( 
.A(n_8643),
.Y(n_9105)
);

NAND2x1p5_ASAP7_75t_L g9106 ( 
.A(n_8151),
.B(n_7565),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_7750),
.Y(n_9107)
);

NAND2xp5_ASAP7_75t_L g9108 ( 
.A(n_8887),
.B(n_6863),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_7750),
.Y(n_9109)
);

INVx6_ASAP7_75t_L g9110 ( 
.A(n_8368),
.Y(n_9110)
);

INVx1_ASAP7_75t_L g9111 ( 
.A(n_7757),
.Y(n_9111)
);

NAND2xp5_ASAP7_75t_L g9112 ( 
.A(n_8887),
.B(n_6884),
.Y(n_9112)
);

INVx1_ASAP7_75t_L g9113 ( 
.A(n_7757),
.Y(n_9113)
);

AND2x4_ASAP7_75t_SL g9114 ( 
.A(n_8806),
.B(n_7153),
.Y(n_9114)
);

OAI21xp5_ASAP7_75t_L g9115 ( 
.A1(n_8055),
.A2(n_7229),
.B(n_7279),
.Y(n_9115)
);

INVx1_ASAP7_75t_L g9116 ( 
.A(n_7760),
.Y(n_9116)
);

BUFx2_ASAP7_75t_L g9117 ( 
.A(n_7786),
.Y(n_9117)
);

AOI22xp33_ASAP7_75t_L g9118 ( 
.A1(n_8055),
.A2(n_6660),
.B1(n_7125),
.B2(n_7547),
.Y(n_9118)
);

INVxp67_ASAP7_75t_L g9119 ( 
.A(n_8521),
.Y(n_9119)
);

NAND2xp5_ASAP7_75t_L g9120 ( 
.A(n_8996),
.B(n_6884),
.Y(n_9120)
);

NOR2xp33_ASAP7_75t_L g9121 ( 
.A(n_8847),
.B(n_7153),
.Y(n_9121)
);

INVx2_ASAP7_75t_L g9122 ( 
.A(n_9001),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_9001),
.Y(n_9123)
);

INVx1_ASAP7_75t_L g9124 ( 
.A(n_7760),
.Y(n_9124)
);

AND2x2_ASAP7_75t_L g9125 ( 
.A(n_8045),
.B(n_6944),
.Y(n_9125)
);

OA21x2_ASAP7_75t_L g9126 ( 
.A1(n_7873),
.A2(n_7486),
.B(n_7247),
.Y(n_9126)
);

AOI22xp33_ASAP7_75t_SL g9127 ( 
.A1(n_8056),
.A2(n_7547),
.B1(n_7351),
.B2(n_7346),
.Y(n_9127)
);

OAI21x1_ASAP7_75t_L g9128 ( 
.A1(n_9003),
.A2(n_7565),
.B(n_7444),
.Y(n_9128)
);

INVx1_ASAP7_75t_L g9129 ( 
.A(n_7763),
.Y(n_9129)
);

BUFx6f_ASAP7_75t_L g9130 ( 
.A(n_8974),
.Y(n_9130)
);

BUFx3_ASAP7_75t_L g9131 ( 
.A(n_8974),
.Y(n_9131)
);

AND2x4_ASAP7_75t_L g9132 ( 
.A(n_8696),
.B(n_8759),
.Y(n_9132)
);

HB1xp67_ASAP7_75t_L g9133 ( 
.A(n_7758),
.Y(n_9133)
);

AO21x2_ASAP7_75t_L g9134 ( 
.A1(n_7705),
.A2(n_7486),
.B(n_7247),
.Y(n_9134)
);

BUFx2_ASAP7_75t_R g9135 ( 
.A(n_8237),
.Y(n_9135)
);

BUFx8_ASAP7_75t_SL g9136 ( 
.A(n_8974),
.Y(n_9136)
);

OAI22xp33_ASAP7_75t_L g9137 ( 
.A1(n_7769),
.A2(n_7352),
.B1(n_7359),
.B2(n_6808),
.Y(n_9137)
);

INVx1_ASAP7_75t_L g9138 ( 
.A(n_7763),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_7784),
.Y(n_9139)
);

CKINVDCx5p33_ASAP7_75t_R g9140 ( 
.A(n_8016),
.Y(n_9140)
);

INVx3_ASAP7_75t_L g9141 ( 
.A(n_7771),
.Y(n_9141)
);

OR2x2_ASAP7_75t_L g9142 ( 
.A(n_8815),
.B(n_7030),
.Y(n_9142)
);

NAND2xp5_ASAP7_75t_L g9143 ( 
.A(n_8996),
.B(n_6884),
.Y(n_9143)
);

INVx1_ASAP7_75t_SL g9144 ( 
.A(n_7817),
.Y(n_9144)
);

BUFx2_ASAP7_75t_L g9145 ( 
.A(n_7786),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_8625),
.Y(n_9146)
);

INVx3_ASAP7_75t_L g9147 ( 
.A(n_7771),
.Y(n_9147)
);

INVx2_ASAP7_75t_L g9148 ( 
.A(n_8625),
.Y(n_9148)
);

AOI22xp33_ASAP7_75t_SL g9149 ( 
.A1(n_8056),
.A2(n_7547),
.B1(n_7351),
.B2(n_7125),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_7784),
.Y(n_9150)
);

INVx1_ASAP7_75t_L g9151 ( 
.A(n_7793),
.Y(n_9151)
);

INVx2_ASAP7_75t_L g9152 ( 
.A(n_8625),
.Y(n_9152)
);

INVx1_ASAP7_75t_L g9153 ( 
.A(n_7793),
.Y(n_9153)
);

AOI21x1_ASAP7_75t_L g9154 ( 
.A1(n_7998),
.A2(n_7619),
.B(n_7511),
.Y(n_9154)
);

NAND2xp5_ASAP7_75t_L g9155 ( 
.A(n_7736),
.B(n_7159),
.Y(n_9155)
);

BUFx3_ASAP7_75t_L g9156 ( 
.A(n_8981),
.Y(n_9156)
);

INVx6_ASAP7_75t_L g9157 ( 
.A(n_8368),
.Y(n_9157)
);

NAND2xp5_ASAP7_75t_L g9158 ( 
.A(n_7736),
.B(n_7159),
.Y(n_9158)
);

BUFx2_ASAP7_75t_L g9159 ( 
.A(n_7786),
.Y(n_9159)
);

INVx2_ASAP7_75t_SL g9160 ( 
.A(n_7771),
.Y(n_9160)
);

CKINVDCx20_ASAP7_75t_R g9161 ( 
.A(n_8854),
.Y(n_9161)
);

AO21x1_ASAP7_75t_L g9162 ( 
.A1(n_7713),
.A2(n_7024),
.B(n_6729),
.Y(n_9162)
);

AND2x4_ASAP7_75t_L g9163 ( 
.A(n_8696),
.B(n_6944),
.Y(n_9163)
);

HB1xp67_ASAP7_75t_L g9164 ( 
.A(n_7787),
.Y(n_9164)
);

INVx3_ASAP7_75t_L g9165 ( 
.A(n_7977),
.Y(n_9165)
);

AND2x2_ASAP7_75t_L g9166 ( 
.A(n_8045),
.B(n_6944),
.Y(n_9166)
);

BUFx6f_ASAP7_75t_L g9167 ( 
.A(n_8981),
.Y(n_9167)
);

INVx1_ASAP7_75t_L g9168 ( 
.A(n_7802),
.Y(n_9168)
);

INVx1_ASAP7_75t_L g9169 ( 
.A(n_7802),
.Y(n_9169)
);

NAND2xp5_ASAP7_75t_L g9170 ( 
.A(n_7770),
.B(n_7193),
.Y(n_9170)
);

AOI22xp33_ASAP7_75t_L g9171 ( 
.A1(n_7855),
.A2(n_7547),
.B1(n_7650),
.B2(n_7634),
.Y(n_9171)
);

NAND2xp5_ASAP7_75t_L g9172 ( 
.A(n_7770),
.B(n_7193),
.Y(n_9172)
);

INVx6_ASAP7_75t_L g9173 ( 
.A(n_8368),
.Y(n_9173)
);

AND2x4_ASAP7_75t_L g9174 ( 
.A(n_8696),
.B(n_6944),
.Y(n_9174)
);

INVx2_ASAP7_75t_L g9175 ( 
.A(n_8655),
.Y(n_9175)
);

INVx1_ASAP7_75t_L g9176 ( 
.A(n_7804),
.Y(n_9176)
);

INVx1_ASAP7_75t_L g9177 ( 
.A(n_7804),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_7822),
.Y(n_9178)
);

INVx2_ASAP7_75t_L g9179 ( 
.A(n_8655),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_8655),
.Y(n_9180)
);

HB1xp67_ASAP7_75t_L g9181 ( 
.A(n_7787),
.Y(n_9181)
);

BUFx6f_ASAP7_75t_L g9182 ( 
.A(n_8981),
.Y(n_9182)
);

INVx1_ASAP7_75t_L g9183 ( 
.A(n_7822),
.Y(n_9183)
);

INVx1_ASAP7_75t_L g9184 ( 
.A(n_7846),
.Y(n_9184)
);

INVx1_ASAP7_75t_L g9185 ( 
.A(n_7846),
.Y(n_9185)
);

OAI21xp5_ASAP7_75t_L g9186 ( 
.A1(n_8220),
.A2(n_7309),
.B(n_7359),
.Y(n_9186)
);

INVx1_ASAP7_75t_L g9187 ( 
.A(n_7862),
.Y(n_9187)
);

INVx6_ASAP7_75t_L g9188 ( 
.A(n_8368),
.Y(n_9188)
);

INVx2_ASAP7_75t_L g9189 ( 
.A(n_8730),
.Y(n_9189)
);

INVx6_ASAP7_75t_L g9190 ( 
.A(n_8368),
.Y(n_9190)
);

INVx1_ASAP7_75t_L g9191 ( 
.A(n_7862),
.Y(n_9191)
);

AOI22xp33_ASAP7_75t_L g9192 ( 
.A1(n_7855),
.A2(n_7547),
.B1(n_7650),
.B2(n_7634),
.Y(n_9192)
);

OAI22xp33_ASAP7_75t_L g9193 ( 
.A1(n_7769),
.A2(n_6808),
.B1(n_6714),
.B2(n_7309),
.Y(n_9193)
);

AOI21x1_ASAP7_75t_L g9194 ( 
.A1(n_7998),
.A2(n_7619),
.B(n_7511),
.Y(n_9194)
);

INVx2_ASAP7_75t_L g9195 ( 
.A(n_8730),
.Y(n_9195)
);

OAI21x1_ASAP7_75t_L g9196 ( 
.A1(n_8229),
.A2(n_6856),
.B(n_6849),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_7867),
.Y(n_9197)
);

AND2x4_ASAP7_75t_L g9198 ( 
.A(n_8759),
.B(n_6946),
.Y(n_9198)
);

OAI22xp33_ASAP7_75t_L g9199 ( 
.A1(n_7911),
.A2(n_6808),
.B1(n_6714),
.B2(n_7309),
.Y(n_9199)
);

HB1xp67_ASAP7_75t_L g9200 ( 
.A(n_7811),
.Y(n_9200)
);

AOI22xp33_ASAP7_75t_L g9201 ( 
.A1(n_7783),
.A2(n_7650),
.B1(n_7634),
.B2(n_7518),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_7867),
.Y(n_9202)
);

OR2x6_ASAP7_75t_L g9203 ( 
.A(n_8235),
.B(n_7458),
.Y(n_9203)
);

OAI21x1_ASAP7_75t_L g9204 ( 
.A1(n_8229),
.A2(n_6856),
.B(n_6849),
.Y(n_9204)
);

AO22x1_ASAP7_75t_L g9205 ( 
.A1(n_7713),
.A2(n_6925),
.B1(n_6878),
.B2(n_6991),
.Y(n_9205)
);

OAI22xp5_ASAP7_75t_L g9206 ( 
.A1(n_7790),
.A2(n_7577),
.B1(n_7539),
.B2(n_7545),
.Y(n_9206)
);

NAND2x1p5_ASAP7_75t_L g9207 ( 
.A(n_8151),
.B(n_7117),
.Y(n_9207)
);

INVx1_ASAP7_75t_L g9208 ( 
.A(n_7879),
.Y(n_9208)
);

INVx2_ASAP7_75t_L g9209 ( 
.A(n_8730),
.Y(n_9209)
);

BUFx4f_ASAP7_75t_SL g9210 ( 
.A(n_8854),
.Y(n_9210)
);

CKINVDCx6p67_ASAP7_75t_R g9211 ( 
.A(n_7953),
.Y(n_9211)
);

BUFx6f_ASAP7_75t_L g9212 ( 
.A(n_9009),
.Y(n_9212)
);

INVx1_ASAP7_75t_L g9213 ( 
.A(n_7879),
.Y(n_9213)
);

HB1xp67_ASAP7_75t_L g9214 ( 
.A(n_7811),
.Y(n_9214)
);

INVx2_ASAP7_75t_L g9215 ( 
.A(n_8730),
.Y(n_9215)
);

INVx6_ASAP7_75t_L g9216 ( 
.A(n_8537),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_7884),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_7884),
.Y(n_9218)
);

AND2x4_ASAP7_75t_L g9219 ( 
.A(n_8759),
.B(n_6946),
.Y(n_9219)
);

INVx1_ASAP7_75t_L g9220 ( 
.A(n_7887),
.Y(n_9220)
);

AND2x2_ASAP7_75t_L g9221 ( 
.A(n_8045),
.B(n_6946),
.Y(n_9221)
);

INVx2_ASAP7_75t_L g9222 ( 
.A(n_8730),
.Y(n_9222)
);

CKINVDCx5p33_ASAP7_75t_R g9223 ( 
.A(n_8016),
.Y(n_9223)
);

HB1xp67_ASAP7_75t_L g9224 ( 
.A(n_7883),
.Y(n_9224)
);

INVx1_ASAP7_75t_L g9225 ( 
.A(n_7887),
.Y(n_9225)
);

OAI21x1_ASAP7_75t_L g9226 ( 
.A1(n_8229),
.A2(n_6868),
.B(n_6856),
.Y(n_9226)
);

BUFx4_ASAP7_75t_SL g9227 ( 
.A(n_8875),
.Y(n_9227)
);

OA21x2_ASAP7_75t_L g9228 ( 
.A1(n_7873),
.A2(n_7619),
.B(n_7511),
.Y(n_9228)
);

AO21x1_ASAP7_75t_SL g9229 ( 
.A1(n_7875),
.A2(n_7577),
.B(n_6714),
.Y(n_9229)
);

AO21x2_ASAP7_75t_L g9230 ( 
.A1(n_7705),
.A2(n_7334),
.B(n_6639),
.Y(n_9230)
);

AO21x1_ASAP7_75t_L g9231 ( 
.A1(n_7762),
.A2(n_7448),
.B(n_7413),
.Y(n_9231)
);

BUFx2_ASAP7_75t_L g9232 ( 
.A(n_7786),
.Y(n_9232)
);

INVx1_ASAP7_75t_L g9233 ( 
.A(n_7891),
.Y(n_9233)
);

AOI22xp33_ASAP7_75t_SL g9234 ( 
.A1(n_8650),
.A2(n_7351),
.B1(n_7127),
.B2(n_7220),
.Y(n_9234)
);

OAI22xp33_ASAP7_75t_SL g9235 ( 
.A1(n_8284),
.A2(n_7288),
.B1(n_7297),
.B2(n_7061),
.Y(n_9235)
);

AOI21x1_ASAP7_75t_L g9236 ( 
.A1(n_8107),
.A2(n_6637),
.B(n_6626),
.Y(n_9236)
);

INVx2_ASAP7_75t_L g9237 ( 
.A(n_8734),
.Y(n_9237)
);

AND2x2_ASAP7_75t_L g9238 ( 
.A(n_8057),
.B(n_6946),
.Y(n_9238)
);

INVx1_ASAP7_75t_L g9239 ( 
.A(n_7891),
.Y(n_9239)
);

AOI22xp33_ASAP7_75t_L g9240 ( 
.A1(n_7783),
.A2(n_7650),
.B1(n_7634),
.B2(n_7518),
.Y(n_9240)
);

AOI21xp5_ASAP7_75t_L g9241 ( 
.A1(n_8078),
.A2(n_7430),
.B(n_7413),
.Y(n_9241)
);

AOI22xp33_ASAP7_75t_L g9242 ( 
.A1(n_8182),
.A2(n_7634),
.B1(n_7650),
.B2(n_7127),
.Y(n_9242)
);

INVx1_ASAP7_75t_L g9243 ( 
.A(n_7897),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_7897),
.Y(n_9244)
);

AOI22xp33_ASAP7_75t_L g9245 ( 
.A1(n_8182),
.A2(n_7634),
.B1(n_7650),
.B2(n_7127),
.Y(n_9245)
);

HB1xp67_ASAP7_75t_L g9246 ( 
.A(n_7883),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_7898),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_7898),
.Y(n_9248)
);

INVx1_ASAP7_75t_SL g9249 ( 
.A(n_7817),
.Y(n_9249)
);

AOI22xp33_ASAP7_75t_SL g9250 ( 
.A1(n_8650),
.A2(n_7714),
.B1(n_8257),
.B2(n_8182),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_7899),
.Y(n_9251)
);

OAI21xp5_ASAP7_75t_SL g9252 ( 
.A1(n_7746),
.A2(n_7424),
.B(n_7151),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_7899),
.Y(n_9253)
);

BUFx12f_ASAP7_75t_L g9254 ( 
.A(n_8093),
.Y(n_9254)
);

INVx1_ASAP7_75t_SL g9255 ( 
.A(n_7924),
.Y(n_9255)
);

INVx2_ASAP7_75t_L g9256 ( 
.A(n_8734),
.Y(n_9256)
);

INVx2_ASAP7_75t_L g9257 ( 
.A(n_8734),
.Y(n_9257)
);

AOI22xp33_ASAP7_75t_SL g9258 ( 
.A1(n_8650),
.A2(n_7351),
.B1(n_7220),
.B2(n_7249),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_7904),
.Y(n_9259)
);

HB1xp67_ASAP7_75t_L g9260 ( 
.A(n_7893),
.Y(n_9260)
);

OAI22xp5_ASAP7_75t_L g9261 ( 
.A1(n_7790),
.A2(n_7539),
.B1(n_7545),
.B2(n_7455),
.Y(n_9261)
);

AOI22xp33_ASAP7_75t_SL g9262 ( 
.A1(n_8650),
.A2(n_7180),
.B1(n_7674),
.B2(n_7249),
.Y(n_9262)
);

INVx6_ASAP7_75t_L g9263 ( 
.A(n_8537),
.Y(n_9263)
);

INVx2_ASAP7_75t_L g9264 ( 
.A(n_8734),
.Y(n_9264)
);

AOI22xp33_ASAP7_75t_L g9265 ( 
.A1(n_8054),
.A2(n_7448),
.B1(n_7550),
.B2(n_7029),
.Y(n_9265)
);

AND2x2_ASAP7_75t_L g9266 ( 
.A(n_8057),
.B(n_6953),
.Y(n_9266)
);

AOI22xp33_ASAP7_75t_L g9267 ( 
.A1(n_8054),
.A2(n_7550),
.B1(n_7029),
.B2(n_7704),
.Y(n_9267)
);

AOI21x1_ASAP7_75t_L g9268 ( 
.A1(n_8107),
.A2(n_6637),
.B(n_6626),
.Y(n_9268)
);

INVx2_ASAP7_75t_L g9269 ( 
.A(n_8734),
.Y(n_9269)
);

OAI21x1_ASAP7_75t_L g9270 ( 
.A1(n_8335),
.A2(n_6868),
.B(n_6856),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_7904),
.Y(n_9271)
);

INVx1_ASAP7_75t_L g9272 ( 
.A(n_7913),
.Y(n_9272)
);

BUFx2_ASAP7_75t_L g9273 ( 
.A(n_7786),
.Y(n_9273)
);

NOR2xp33_ASAP7_75t_L g9274 ( 
.A(n_8957),
.B(n_7153),
.Y(n_9274)
);

AOI21x1_ASAP7_75t_L g9275 ( 
.A1(n_8107),
.A2(n_6637),
.B(n_6626),
.Y(n_9275)
);

CKINVDCx20_ASAP7_75t_R g9276 ( 
.A(n_8875),
.Y(n_9276)
);

OAI21x1_ASAP7_75t_L g9277 ( 
.A1(n_8335),
.A2(n_8632),
.B(n_8346),
.Y(n_9277)
);

INVx3_ASAP7_75t_L g9278 ( 
.A(n_7977),
.Y(n_9278)
);

OAI22xp5_ASAP7_75t_L g9279 ( 
.A1(n_7798),
.A2(n_7539),
.B1(n_7545),
.B2(n_7455),
.Y(n_9279)
);

INVx2_ASAP7_75t_L g9280 ( 
.A(n_8756),
.Y(n_9280)
);

INVx4_ASAP7_75t_L g9281 ( 
.A(n_9009),
.Y(n_9281)
);

CKINVDCx5p33_ASAP7_75t_R g9282 ( 
.A(n_8092),
.Y(n_9282)
);

INVx2_ASAP7_75t_SL g9283 ( 
.A(n_8050),
.Y(n_9283)
);

INVx2_ASAP7_75t_L g9284 ( 
.A(n_8756),
.Y(n_9284)
);

INVx4_ASAP7_75t_L g9285 ( 
.A(n_9009),
.Y(n_9285)
);

INVx2_ASAP7_75t_L g9286 ( 
.A(n_8756),
.Y(n_9286)
);

OAI21x1_ASAP7_75t_L g9287 ( 
.A1(n_8335),
.A2(n_6868),
.B(n_6856),
.Y(n_9287)
);

BUFx6f_ASAP7_75t_L g9288 ( 
.A(n_8093),
.Y(n_9288)
);

AND2x2_ASAP7_75t_L g9289 ( 
.A(n_8057),
.B(n_6953),
.Y(n_9289)
);

INVx4_ASAP7_75t_L g9290 ( 
.A(n_8806),
.Y(n_9290)
);

AND2x2_ASAP7_75t_L g9291 ( 
.A(n_8659),
.B(n_6953),
.Y(n_9291)
);

INVx2_ASAP7_75t_L g9292 ( 
.A(n_8756),
.Y(n_9292)
);

INVx1_ASAP7_75t_L g9293 ( 
.A(n_7913),
.Y(n_9293)
);

INVx1_ASAP7_75t_L g9294 ( 
.A(n_7918),
.Y(n_9294)
);

INVx5_ASAP7_75t_L g9295 ( 
.A(n_7977),
.Y(n_9295)
);

CKINVDCx6p67_ASAP7_75t_R g9296 ( 
.A(n_8201),
.Y(n_9296)
);

AND2x4_ASAP7_75t_L g9297 ( 
.A(n_8859),
.B(n_6953),
.Y(n_9297)
);

INVx2_ASAP7_75t_L g9298 ( 
.A(n_8756),
.Y(n_9298)
);

INVx1_ASAP7_75t_L g9299 ( 
.A(n_7918),
.Y(n_9299)
);

INVx2_ASAP7_75t_L g9300 ( 
.A(n_8770),
.Y(n_9300)
);

INVx1_ASAP7_75t_L g9301 ( 
.A(n_7926),
.Y(n_9301)
);

INVx6_ASAP7_75t_L g9302 ( 
.A(n_8537),
.Y(n_9302)
);

BUFx5_ASAP7_75t_L g9303 ( 
.A(n_7964),
.Y(n_9303)
);

INVx2_ASAP7_75t_L g9304 ( 
.A(n_8770),
.Y(n_9304)
);

OAI21x1_ASAP7_75t_L g9305 ( 
.A1(n_8865),
.A2(n_7446),
.B(n_6910),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_7926),
.Y(n_9306)
);

AOI22xp33_ASAP7_75t_L g9307 ( 
.A1(n_8128),
.A2(n_7550),
.B1(n_7704),
.B2(n_7177),
.Y(n_9307)
);

AOI22xp33_ASAP7_75t_SL g9308 ( 
.A1(n_7714),
.A2(n_7674),
.B1(n_7323),
.B2(n_7636),
.Y(n_9308)
);

OAI22xp5_ASAP7_75t_SL g9309 ( 
.A1(n_8128),
.A2(n_8364),
.B1(n_7849),
.B2(n_8834),
.Y(n_9309)
);

CKINVDCx16_ASAP7_75t_R g9310 ( 
.A(n_8123),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_7935),
.Y(n_9311)
);

INVx2_ASAP7_75t_L g9312 ( 
.A(n_8770),
.Y(n_9312)
);

INVx6_ASAP7_75t_L g9313 ( 
.A(n_8537),
.Y(n_9313)
);

AOI22xp33_ASAP7_75t_L g9314 ( 
.A1(n_8153),
.A2(n_7177),
.B1(n_7173),
.B2(n_7041),
.Y(n_9314)
);

NAND2xp5_ASAP7_75t_L g9315 ( 
.A(n_7775),
.B(n_6914),
.Y(n_9315)
);

INVx1_ASAP7_75t_L g9316 ( 
.A(n_7935),
.Y(n_9316)
);

OAI21x1_ASAP7_75t_L g9317 ( 
.A1(n_8865),
.A2(n_7446),
.B(n_6910),
.Y(n_9317)
);

AND2x2_ASAP7_75t_L g9318 ( 
.A(n_8659),
.B(n_6962),
.Y(n_9318)
);

INVx2_ASAP7_75t_L g9319 ( 
.A(n_8770),
.Y(n_9319)
);

INVx1_ASAP7_75t_L g9320 ( 
.A(n_7942),
.Y(n_9320)
);

INVx2_ASAP7_75t_L g9321 ( 
.A(n_8770),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_7942),
.Y(n_9322)
);

INVx1_ASAP7_75t_L g9323 ( 
.A(n_7945),
.Y(n_9323)
);

NAND2xp5_ASAP7_75t_L g9324 ( 
.A(n_7775),
.B(n_6914),
.Y(n_9324)
);

NAND2x1p5_ASAP7_75t_L g9325 ( 
.A(n_7759),
.B(n_7117),
.Y(n_9325)
);

AOI22xp33_ASAP7_75t_SL g9326 ( 
.A1(n_8257),
.A2(n_7674),
.B1(n_7323),
.B2(n_7636),
.Y(n_9326)
);

INVx1_ASAP7_75t_L g9327 ( 
.A(n_7945),
.Y(n_9327)
);

NAND2xp33_ASAP7_75t_SL g9328 ( 
.A(n_8888),
.B(n_7525),
.Y(n_9328)
);

OAI22xp5_ASAP7_75t_L g9329 ( 
.A1(n_7798),
.A2(n_7061),
.B1(n_7297),
.B2(n_7288),
.Y(n_9329)
);

OAI21x1_ASAP7_75t_L g9330 ( 
.A1(n_8335),
.A2(n_6868),
.B(n_6856),
.Y(n_9330)
);

INVx1_ASAP7_75t_L g9331 ( 
.A(n_7971),
.Y(n_9331)
);

INVx2_ASAP7_75t_L g9332 ( 
.A(n_7786),
.Y(n_9332)
);

HB1xp67_ASAP7_75t_L g9333 ( 
.A(n_7893),
.Y(n_9333)
);

AOI22xp33_ASAP7_75t_L g9334 ( 
.A1(n_8153),
.A2(n_7173),
.B1(n_7041),
.B2(n_7226),
.Y(n_9334)
);

INVx4_ASAP7_75t_L g9335 ( 
.A(n_8806),
.Y(n_9335)
);

HB1xp67_ASAP7_75t_L g9336 ( 
.A(n_7959),
.Y(n_9336)
);

INVx2_ASAP7_75t_L g9337 ( 
.A(n_7786),
.Y(n_9337)
);

BUFx8_ASAP7_75t_L g9338 ( 
.A(n_8023),
.Y(n_9338)
);

INVx1_ASAP7_75t_L g9339 ( 
.A(n_7971),
.Y(n_9339)
);

AOI22xp33_ASAP7_75t_SL g9340 ( 
.A1(n_8220),
.A2(n_7323),
.B1(n_7636),
.B2(n_7620),
.Y(n_9340)
);

AND2x2_ASAP7_75t_L g9341 ( 
.A(n_8659),
.B(n_6962),
.Y(n_9341)
);

BUFx2_ASAP7_75t_L g9342 ( 
.A(n_7786),
.Y(n_9342)
);

CKINVDCx20_ASAP7_75t_R g9343 ( 
.A(n_7730),
.Y(n_9343)
);

INVx2_ASAP7_75t_L g9344 ( 
.A(n_9026),
.Y(n_9344)
);

AO21x2_ASAP7_75t_L g9345 ( 
.A1(n_7851),
.A2(n_6639),
.B(n_6629),
.Y(n_9345)
);

INVx1_ASAP7_75t_L g9346 ( 
.A(n_7972),
.Y(n_9346)
);

OAI22x1_ASAP7_75t_L g9347 ( 
.A1(n_8321),
.A2(n_6925),
.B1(n_6878),
.B2(n_7617),
.Y(n_9347)
);

AOI22xp33_ASAP7_75t_L g9348 ( 
.A1(n_8153),
.A2(n_7738),
.B1(n_8397),
.B2(n_7922),
.Y(n_9348)
);

NAND2xp5_ASAP7_75t_L g9349 ( 
.A(n_7801),
.B(n_8299),
.Y(n_9349)
);

AO21x1_ASAP7_75t_L g9350 ( 
.A1(n_7762),
.A2(n_7143),
.B(n_7088),
.Y(n_9350)
);

OA21x2_ASAP7_75t_L g9351 ( 
.A1(n_7819),
.A2(n_6712),
.B(n_6628),
.Y(n_9351)
);

AO21x2_ASAP7_75t_L g9352 ( 
.A1(n_7851),
.A2(n_6639),
.B(n_6629),
.Y(n_9352)
);

CKINVDCx5p33_ASAP7_75t_R g9353 ( 
.A(n_8092),
.Y(n_9353)
);

NAND2xp5_ASAP7_75t_L g9354 ( 
.A(n_7801),
.B(n_8299),
.Y(n_9354)
);

AOI22xp33_ASAP7_75t_L g9355 ( 
.A1(n_7738),
.A2(n_7226),
.B1(n_7307),
.B2(n_7263),
.Y(n_9355)
);

AOI22xp33_ASAP7_75t_SL g9356 ( 
.A1(n_7922),
.A2(n_7668),
.B1(n_7685),
.B2(n_7620),
.Y(n_9356)
);

AOI22xp33_ASAP7_75t_L g9357 ( 
.A1(n_8397),
.A2(n_7226),
.B1(n_7307),
.B2(n_7263),
.Y(n_9357)
);

AOI22xp33_ASAP7_75t_L g9358 ( 
.A1(n_8364),
.A2(n_8292),
.B1(n_7799),
.B2(n_7896),
.Y(n_9358)
);

INVx11_ASAP7_75t_L g9359 ( 
.A(n_8537),
.Y(n_9359)
);

OAI22xp5_ASAP7_75t_L g9360 ( 
.A1(n_7748),
.A2(n_7061),
.B1(n_7297),
.B2(n_7288),
.Y(n_9360)
);

CKINVDCx5p33_ASAP7_75t_R g9361 ( 
.A(n_7730),
.Y(n_9361)
);

AND2x4_ASAP7_75t_L g9362 ( 
.A(n_8859),
.B(n_6962),
.Y(n_9362)
);

INVx3_ASAP7_75t_L g9363 ( 
.A(n_7977),
.Y(n_9363)
);

OAI22xp33_ASAP7_75t_L g9364 ( 
.A1(n_7911),
.A2(n_7424),
.B1(n_6779),
.B2(n_7554),
.Y(n_9364)
);

INVx4_ASAP7_75t_L g9365 ( 
.A(n_8898),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_7972),
.Y(n_9366)
);

INVx1_ASAP7_75t_L g9367 ( 
.A(n_7974),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_7974),
.Y(n_9368)
);

AOI22xp33_ASAP7_75t_L g9369 ( 
.A1(n_8292),
.A2(n_7226),
.B1(n_7307),
.B2(n_7266),
.Y(n_9369)
);

INVxp67_ASAP7_75t_SL g9370 ( 
.A(n_8254),
.Y(n_9370)
);

INVx2_ASAP7_75t_L g9371 ( 
.A(n_9026),
.Y(n_9371)
);

INVx1_ASAP7_75t_L g9372 ( 
.A(n_7976),
.Y(n_9372)
);

OA21x2_ASAP7_75t_L g9373 ( 
.A1(n_7819),
.A2(n_6712),
.B(n_6628),
.Y(n_9373)
);

NOR2xp67_ASAP7_75t_SL g9374 ( 
.A(n_8351),
.B(n_7500),
.Y(n_9374)
);

OAI22xp33_ASAP7_75t_R g9375 ( 
.A1(n_7754),
.A2(n_7814),
.B1(n_8631),
.B2(n_7840),
.Y(n_9375)
);

INVx1_ASAP7_75t_L g9376 ( 
.A(n_7976),
.Y(n_9376)
);

AOI22xp33_ASAP7_75t_L g9377 ( 
.A1(n_7799),
.A2(n_7226),
.B1(n_7307),
.B2(n_7266),
.Y(n_9377)
);

INVx3_ASAP7_75t_L g9378 ( 
.A(n_7977),
.Y(n_9378)
);

INVx1_ASAP7_75t_L g9379 ( 
.A(n_7982),
.Y(n_9379)
);

BUFx2_ASAP7_75t_SL g9380 ( 
.A(n_8351),
.Y(n_9380)
);

AOI22xp33_ASAP7_75t_SL g9381 ( 
.A1(n_8028),
.A2(n_7668),
.B1(n_7685),
.B2(n_7620),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_7982),
.Y(n_9382)
);

NAND2xp5_ASAP7_75t_L g9383 ( 
.A(n_7934),
.B(n_6915),
.Y(n_9383)
);

HB1xp67_ASAP7_75t_L g9384 ( 
.A(n_7959),
.Y(n_9384)
);

INVx1_ASAP7_75t_L g9385 ( 
.A(n_7990),
.Y(n_9385)
);

BUFx2_ASAP7_75t_R g9386 ( 
.A(n_8351),
.Y(n_9386)
);

BUFx6f_ASAP7_75t_L g9387 ( 
.A(n_8201),
.Y(n_9387)
);

AOI21x1_ASAP7_75t_L g9388 ( 
.A1(n_7986),
.A2(n_6641),
.B(n_6638),
.Y(n_9388)
);

CKINVDCx20_ASAP7_75t_R g9389 ( 
.A(n_7825),
.Y(n_9389)
);

AOI22xp33_ASAP7_75t_L g9390 ( 
.A1(n_7896),
.A2(n_7226),
.B1(n_7307),
.B2(n_7256),
.Y(n_9390)
);

INVxp67_ASAP7_75t_L g9391 ( 
.A(n_8521),
.Y(n_9391)
);

CKINVDCx20_ASAP7_75t_R g9392 ( 
.A(n_7825),
.Y(n_9392)
);

CKINVDCx20_ASAP7_75t_R g9393 ( 
.A(n_7854),
.Y(n_9393)
);

AND2x2_ASAP7_75t_L g9394 ( 
.A(n_8864),
.B(n_6962),
.Y(n_9394)
);

INVx2_ASAP7_75t_SL g9395 ( 
.A(n_8050),
.Y(n_9395)
);

INVx2_ASAP7_75t_SL g9396 ( 
.A(n_8050),
.Y(n_9396)
);

INVx1_ASAP7_75t_L g9397 ( 
.A(n_7990),
.Y(n_9397)
);

INVx2_ASAP7_75t_L g9398 ( 
.A(n_8964),
.Y(n_9398)
);

INVx2_ASAP7_75t_L g9399 ( 
.A(n_8964),
.Y(n_9399)
);

AND2x2_ASAP7_75t_L g9400 ( 
.A(n_8864),
.B(n_6966),
.Y(n_9400)
);

INVx2_ASAP7_75t_L g9401 ( 
.A(n_8964),
.Y(n_9401)
);

AOI22xp33_ASAP7_75t_SL g9402 ( 
.A1(n_8028),
.A2(n_7685),
.B1(n_7668),
.B2(n_7571),
.Y(n_9402)
);

AO21x1_ASAP7_75t_SL g9403 ( 
.A1(n_7875),
.A2(n_6779),
.B(n_6793),
.Y(n_9403)
);

INVx1_ASAP7_75t_L g9404 ( 
.A(n_7996),
.Y(n_9404)
);

AOI22xp33_ASAP7_75t_L g9405 ( 
.A1(n_7833),
.A2(n_7710),
.B1(n_7837),
.B2(n_7728),
.Y(n_9405)
);

BUFx2_ASAP7_75t_R g9406 ( 
.A(n_8679),
.Y(n_9406)
);

INVx1_ASAP7_75t_L g9407 ( 
.A(n_7996),
.Y(n_9407)
);

INVx1_ASAP7_75t_L g9408 ( 
.A(n_8000),
.Y(n_9408)
);

NAND2xp5_ASAP7_75t_L g9409 ( 
.A(n_7934),
.B(n_6915),
.Y(n_9409)
);

INVx6_ASAP7_75t_L g9410 ( 
.A(n_7850),
.Y(n_9410)
);

INVx2_ASAP7_75t_L g9411 ( 
.A(n_9026),
.Y(n_9411)
);

INVx2_ASAP7_75t_L g9412 ( 
.A(n_9026),
.Y(n_9412)
);

HB1xp67_ASAP7_75t_L g9413 ( 
.A(n_8010),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_8000),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8019),
.Y(n_9415)
);

NAND2xp5_ASAP7_75t_L g9416 ( 
.A(n_7838),
.B(n_7399),
.Y(n_9416)
);

INVx1_ASAP7_75t_L g9417 ( 
.A(n_8019),
.Y(n_9417)
);

OAI21xp5_ASAP7_75t_L g9418 ( 
.A1(n_7748),
.A2(n_7299),
.B(n_7621),
.Y(n_9418)
);

OAI21x1_ASAP7_75t_L g9419 ( 
.A1(n_8907),
.A2(n_7446),
.B(n_6872),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_8030),
.Y(n_9420)
);

INVx1_ASAP7_75t_L g9421 ( 
.A(n_8030),
.Y(n_9421)
);

HB1xp67_ASAP7_75t_L g9422 ( 
.A(n_8010),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8032),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_8032),
.Y(n_9424)
);

AO21x2_ASAP7_75t_L g9425 ( 
.A1(n_7819),
.A2(n_6629),
.B(n_6628),
.Y(n_9425)
);

OA21x2_ASAP7_75t_L g9426 ( 
.A1(n_8029),
.A2(n_6822),
.B(n_6816),
.Y(n_9426)
);

INVx2_ASAP7_75t_L g9427 ( 
.A(n_8964),
.Y(n_9427)
);

INVx1_ASAP7_75t_L g9428 ( 
.A(n_8040),
.Y(n_9428)
);

BUFx3_ASAP7_75t_L g9429 ( 
.A(n_8242),
.Y(n_9429)
);

CKINVDCx20_ASAP7_75t_R g9430 ( 
.A(n_7854),
.Y(n_9430)
);

AOI22xp33_ASAP7_75t_L g9431 ( 
.A1(n_7833),
.A2(n_7307),
.B1(n_7256),
.B2(n_7498),
.Y(n_9431)
);

AOI22xp33_ASAP7_75t_L g9432 ( 
.A1(n_7710),
.A2(n_7307),
.B1(n_7507),
.B2(n_7498),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_8040),
.Y(n_9433)
);

BUFx12f_ASAP7_75t_L g9434 ( 
.A(n_8242),
.Y(n_9434)
);

INVx2_ASAP7_75t_L g9435 ( 
.A(n_8964),
.Y(n_9435)
);

HB1xp67_ASAP7_75t_L g9436 ( 
.A(n_8034),
.Y(n_9436)
);

INVx2_ASAP7_75t_L g9437 ( 
.A(n_9019),
.Y(n_9437)
);

INVx3_ASAP7_75t_L g9438 ( 
.A(n_7977),
.Y(n_9438)
);

BUFx3_ASAP7_75t_L g9439 ( 
.A(n_8976),
.Y(n_9439)
);

INVx2_ASAP7_75t_L g9440 ( 
.A(n_9019),
.Y(n_9440)
);

INVx2_ASAP7_75t_L g9441 ( 
.A(n_9019),
.Y(n_9441)
);

CKINVDCx11_ASAP7_75t_R g9442 ( 
.A(n_7876),
.Y(n_9442)
);

INVx2_ASAP7_75t_L g9443 ( 
.A(n_9019),
.Y(n_9443)
);

BUFx12f_ASAP7_75t_L g9444 ( 
.A(n_8976),
.Y(n_9444)
);

AO21x2_ASAP7_75t_L g9445 ( 
.A1(n_8078),
.A2(n_6641),
.B(n_6638),
.Y(n_9445)
);

INVx1_ASAP7_75t_SL g9446 ( 
.A(n_7924),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_8052),
.Y(n_9447)
);

BUFx2_ASAP7_75t_R g9448 ( 
.A(n_8049),
.Y(n_9448)
);

OR2x6_ASAP7_75t_L g9449 ( 
.A(n_8459),
.B(n_6807),
.Y(n_9449)
);

AOI22xp33_ASAP7_75t_L g9450 ( 
.A1(n_7837),
.A2(n_7307),
.B1(n_7507),
.B2(n_7021),
.Y(n_9450)
);

HB1xp67_ASAP7_75t_L g9451 ( 
.A(n_8034),
.Y(n_9451)
);

HB1xp67_ASAP7_75t_L g9452 ( 
.A(n_8075),
.Y(n_9452)
);

OAI22xp5_ASAP7_75t_L g9453 ( 
.A1(n_8321),
.A2(n_7061),
.B1(n_7297),
.B2(n_7288),
.Y(n_9453)
);

CKINVDCx6p67_ASAP7_75t_R g9454 ( 
.A(n_7821),
.Y(n_9454)
);

INVx11_ASAP7_75t_L g9455 ( 
.A(n_8023),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_8052),
.Y(n_9456)
);

AOI22xp33_ASAP7_75t_L g9457 ( 
.A1(n_7728),
.A2(n_7021),
.B1(n_6727),
.B2(n_6732),
.Y(n_9457)
);

NAND2x1p5_ASAP7_75t_L g9458 ( 
.A(n_7759),
.B(n_7117),
.Y(n_9458)
);

AOI22xp5_ASAP7_75t_SL g9459 ( 
.A1(n_7871),
.A2(n_7675),
.B1(n_7525),
.B2(n_7627),
.Y(n_9459)
);

OAI22xp33_ASAP7_75t_SL g9460 ( 
.A1(n_8284),
.A2(n_7533),
.B1(n_7405),
.B2(n_6816),
.Y(n_9460)
);

AOI21x1_ASAP7_75t_L g9461 ( 
.A1(n_7986),
.A2(n_6641),
.B(n_6638),
.Y(n_9461)
);

NAND2xp5_ASAP7_75t_L g9462 ( 
.A(n_7838),
.B(n_7399),
.Y(n_9462)
);

BUFx8_ASAP7_75t_SL g9463 ( 
.A(n_7794),
.Y(n_9463)
);

AND2x2_ASAP7_75t_L g9464 ( 
.A(n_8864),
.B(n_6966),
.Y(n_9464)
);

OAI21x1_ASAP7_75t_L g9465 ( 
.A1(n_8346),
.A2(n_6872),
.B(n_6868),
.Y(n_9465)
);

CKINVDCx8_ASAP7_75t_R g9466 ( 
.A(n_7863),
.Y(n_9466)
);

CKINVDCx11_ASAP7_75t_R g9467 ( 
.A(n_7876),
.Y(n_9467)
);

INVx1_ASAP7_75t_L g9468 ( 
.A(n_8058),
.Y(n_9468)
);

INVx4_ASAP7_75t_L g9469 ( 
.A(n_8898),
.Y(n_9469)
);

INVx1_ASAP7_75t_L g9470 ( 
.A(n_8058),
.Y(n_9470)
);

BUFx8_ASAP7_75t_L g9471 ( 
.A(n_8043),
.Y(n_9471)
);

INVx3_ASAP7_75t_L g9472 ( 
.A(n_7977),
.Y(n_9472)
);

HB1xp67_ASAP7_75t_L g9473 ( 
.A(n_8075),
.Y(n_9473)
);

CKINVDCx5p33_ASAP7_75t_R g9474 ( 
.A(n_7901),
.Y(n_9474)
);

AND2x2_ASAP7_75t_L g9475 ( 
.A(n_8006),
.B(n_6966),
.Y(n_9475)
);

INVx3_ASAP7_75t_L g9476 ( 
.A(n_7977),
.Y(n_9476)
);

INVx1_ASAP7_75t_L g9477 ( 
.A(n_8060),
.Y(n_9477)
);

INVx1_ASAP7_75t_L g9478 ( 
.A(n_8060),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_8061),
.Y(n_9479)
);

AO21x1_ASAP7_75t_SL g9480 ( 
.A1(n_8221),
.A2(n_6779),
.B(n_6793),
.Y(n_9480)
);

AND2x4_ASAP7_75t_L g9481 ( 
.A(n_8859),
.B(n_8933),
.Y(n_9481)
);

INVx1_ASAP7_75t_L g9482 ( 
.A(n_8061),
.Y(n_9482)
);

OAI21xp5_ASAP7_75t_L g9483 ( 
.A1(n_7970),
.A2(n_7299),
.B(n_7621),
.Y(n_9483)
);

AO21x2_ASAP7_75t_L g9484 ( 
.A1(n_8739),
.A2(n_6666),
.B(n_6654),
.Y(n_9484)
);

AOI22xp33_ASAP7_75t_L g9485 ( 
.A1(n_7849),
.A2(n_6727),
.B1(n_6732),
.B2(n_6717),
.Y(n_9485)
);

BUFx2_ASAP7_75t_R g9486 ( 
.A(n_8065),
.Y(n_9486)
);

BUFx10_ASAP7_75t_L g9487 ( 
.A(n_8281),
.Y(n_9487)
);

CKINVDCx6p67_ASAP7_75t_R g9488 ( 
.A(n_7821),
.Y(n_9488)
);

AO21x1_ASAP7_75t_SL g9489 ( 
.A1(n_8221),
.A2(n_6793),
.B(n_7424),
.Y(n_9489)
);

BUFx4f_ASAP7_75t_L g9490 ( 
.A(n_8898),
.Y(n_9490)
);

AOI22xp33_ASAP7_75t_L g9491 ( 
.A1(n_8232),
.A2(n_6727),
.B1(n_6732),
.B2(n_6717),
.Y(n_9491)
);

INVx1_ASAP7_75t_L g9492 ( 
.A(n_8079),
.Y(n_9492)
);

INVx1_ASAP7_75t_SL g9493 ( 
.A(n_7980),
.Y(n_9493)
);

AND2x2_ASAP7_75t_L g9494 ( 
.A(n_8006),
.B(n_6966),
.Y(n_9494)
);

AND2x2_ASAP7_75t_L g9495 ( 
.A(n_8006),
.B(n_6971),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_8079),
.Y(n_9496)
);

AOI22xp33_ASAP7_75t_L g9497 ( 
.A1(n_8232),
.A2(n_6727),
.B1(n_6732),
.B2(n_6717),
.Y(n_9497)
);

BUFx3_ASAP7_75t_L g9498 ( 
.A(n_8024),
.Y(n_9498)
);

CKINVDCx5p33_ASAP7_75t_R g9499 ( 
.A(n_7901),
.Y(n_9499)
);

AOI22xp5_ASAP7_75t_L g9500 ( 
.A1(n_7746),
.A2(n_7340),
.B1(n_6689),
.B2(n_7530),
.Y(n_9500)
);

INVx4_ASAP7_75t_L g9501 ( 
.A(n_8912),
.Y(n_9501)
);

BUFx2_ASAP7_75t_R g9502 ( 
.A(n_8446),
.Y(n_9502)
);

BUFx8_ASAP7_75t_L g9503 ( 
.A(n_8043),
.Y(n_9503)
);

OAI21x1_ASAP7_75t_L g9504 ( 
.A1(n_8346),
.A2(n_6872),
.B(n_6868),
.Y(n_9504)
);

NAND2xp5_ASAP7_75t_L g9505 ( 
.A(n_7900),
.B(n_7399),
.Y(n_9505)
);

AOI21x1_ASAP7_75t_L g9506 ( 
.A1(n_7952),
.A2(n_6666),
.B(n_6654),
.Y(n_9506)
);

AOI22xp33_ASAP7_75t_L g9507 ( 
.A1(n_8866),
.A2(n_6727),
.B1(n_6732),
.B2(n_6717),
.Y(n_9507)
);

INVx1_ASAP7_75t_L g9508 ( 
.A(n_8080),
.Y(n_9508)
);

INVx1_ASAP7_75t_L g9509 ( 
.A(n_8080),
.Y(n_9509)
);

AOI22xp33_ASAP7_75t_L g9510 ( 
.A1(n_8866),
.A2(n_6727),
.B1(n_6732),
.B2(n_6717),
.Y(n_9510)
);

INVx2_ASAP7_75t_L g9511 ( 
.A(n_9026),
.Y(n_9511)
);

AOI22xp33_ASAP7_75t_L g9512 ( 
.A1(n_8543),
.A2(n_7767),
.B1(n_7764),
.B2(n_7795),
.Y(n_9512)
);

AOI22xp33_ASAP7_75t_L g9513 ( 
.A1(n_8543),
.A2(n_6737),
.B1(n_6776),
.B2(n_6717),
.Y(n_9513)
);

INVx5_ASAP7_75t_L g9514 ( 
.A(n_8044),
.Y(n_9514)
);

INVx2_ASAP7_75t_L g9515 ( 
.A(n_9019),
.Y(n_9515)
);

INVx2_ASAP7_75t_SL g9516 ( 
.A(n_8050),
.Y(n_9516)
);

OA21x2_ASAP7_75t_L g9517 ( 
.A1(n_8029),
.A2(n_6822),
.B(n_6816),
.Y(n_9517)
);

BUFx2_ASAP7_75t_SL g9518 ( 
.A(n_8254),
.Y(n_9518)
);

HB1xp67_ASAP7_75t_SL g9519 ( 
.A(n_8765),
.Y(n_9519)
);

INVx2_ASAP7_75t_L g9520 ( 
.A(n_9030),
.Y(n_9520)
);

HB1xp67_ASAP7_75t_L g9521 ( 
.A(n_8101),
.Y(n_9521)
);

NAND2x1p5_ASAP7_75t_L g9522 ( 
.A(n_7759),
.B(n_7133),
.Y(n_9522)
);

OAI22x1_ASAP7_75t_L g9523 ( 
.A1(n_8294),
.A2(n_7627),
.B1(n_7631),
.B2(n_7617),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_8081),
.Y(n_9524)
);

INVx2_ASAP7_75t_L g9525 ( 
.A(n_9030),
.Y(n_9525)
);

BUFx6f_ASAP7_75t_L g9526 ( 
.A(n_8044),
.Y(n_9526)
);

BUFx2_ASAP7_75t_L g9527 ( 
.A(n_8742),
.Y(n_9527)
);

OAI22xp5_ASAP7_75t_L g9528 ( 
.A1(n_7889),
.A2(n_7405),
.B1(n_7533),
.B2(n_7530),
.Y(n_9528)
);

INVx2_ASAP7_75t_L g9529 ( 
.A(n_9030),
.Y(n_9529)
);

OAI22xp33_ASAP7_75t_L g9530 ( 
.A1(n_7946),
.A2(n_8294),
.B1(n_8195),
.B2(n_8117),
.Y(n_9530)
);

HB1xp67_ASAP7_75t_L g9531 ( 
.A(n_8101),
.Y(n_9531)
);

AOI22xp33_ASAP7_75t_SL g9532 ( 
.A1(n_8744),
.A2(n_7571),
.B1(n_7601),
.B2(n_7500),
.Y(n_9532)
);

AOI22xp33_ASAP7_75t_SL g9533 ( 
.A1(n_8744),
.A2(n_7571),
.B1(n_7601),
.B2(n_7500),
.Y(n_9533)
);

NAND2x1p5_ASAP7_75t_L g9534 ( 
.A(n_7759),
.B(n_7133),
.Y(n_9534)
);

AOI22xp33_ASAP7_75t_SL g9535 ( 
.A1(n_7764),
.A2(n_7571),
.B1(n_7601),
.B2(n_7500),
.Y(n_9535)
);

OAI22xp5_ASAP7_75t_L g9536 ( 
.A1(n_7889),
.A2(n_7405),
.B1(n_7533),
.B2(n_6689),
.Y(n_9536)
);

CKINVDCx20_ASAP7_75t_R g9537 ( 
.A(n_7983),
.Y(n_9537)
);

OAI22xp5_ASAP7_75t_L g9538 ( 
.A1(n_7989),
.A2(n_7533),
.B1(n_7405),
.B2(n_7447),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_8081),
.Y(n_9539)
);

INVx2_ASAP7_75t_L g9540 ( 
.A(n_7720),
.Y(n_9540)
);

NAND2x1p5_ASAP7_75t_L g9541 ( 
.A(n_7759),
.B(n_7133),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_8088),
.Y(n_9542)
);

AOI21x1_ASAP7_75t_L g9543 ( 
.A1(n_7952),
.A2(n_6666),
.B(n_6654),
.Y(n_9543)
);

AOI22xp33_ASAP7_75t_SL g9544 ( 
.A1(n_8109),
.A2(n_7615),
.B1(n_7601),
.B2(n_7701),
.Y(n_9544)
);

INVx2_ASAP7_75t_L g9545 ( 
.A(n_7720),
.Y(n_9545)
);

BUFx2_ASAP7_75t_L g9546 ( 
.A(n_8742),
.Y(n_9546)
);

INVx5_ASAP7_75t_L g9547 ( 
.A(n_8044),
.Y(n_9547)
);

INVx1_ASAP7_75t_L g9548 ( 
.A(n_8088),
.Y(n_9548)
);

NAND2xp5_ASAP7_75t_L g9549 ( 
.A(n_7900),
.B(n_7407),
.Y(n_9549)
);

INVxp67_ASAP7_75t_SL g9550 ( 
.A(n_8313),
.Y(n_9550)
);

BUFx2_ASAP7_75t_R g9551 ( 
.A(n_8113),
.Y(n_9551)
);

BUFx2_ASAP7_75t_L g9552 ( 
.A(n_8742),
.Y(n_9552)
);

INVx1_ASAP7_75t_SL g9553 ( 
.A(n_7980),
.Y(n_9553)
);

AOI21x1_ASAP7_75t_L g9554 ( 
.A1(n_7952),
.A2(n_6696),
.B(n_6687),
.Y(n_9554)
);

INVx2_ASAP7_75t_SL g9555 ( 
.A(n_8050),
.Y(n_9555)
);

AOI22xp33_ASAP7_75t_L g9556 ( 
.A1(n_7767),
.A2(n_7795),
.B1(n_8136),
.B2(n_8164),
.Y(n_9556)
);

OAI22xp5_ASAP7_75t_L g9557 ( 
.A1(n_7989),
.A2(n_7946),
.B1(n_8768),
.B2(n_7950),
.Y(n_9557)
);

AO21x1_ASAP7_75t_L g9558 ( 
.A1(n_8972),
.A2(n_7143),
.B(n_7088),
.Y(n_9558)
);

NAND2xp5_ASAP7_75t_L g9559 ( 
.A(n_8532),
.B(n_7407),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_8089),
.Y(n_9560)
);

NAND2xp33_ASAP7_75t_SL g9561 ( 
.A(n_8888),
.B(n_7675),
.Y(n_9561)
);

NAND2xp5_ASAP7_75t_L g9562 ( 
.A(n_8532),
.B(n_7407),
.Y(n_9562)
);

AOI22xp33_ASAP7_75t_L g9563 ( 
.A1(n_7795),
.A2(n_6776),
.B1(n_6737),
.B2(n_7485),
.Y(n_9563)
);

NAND2x1p5_ASAP7_75t_L g9564 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9564)
);

OAI21x1_ASAP7_75t_SL g9565 ( 
.A1(n_8313),
.A2(n_7519),
.B(n_7502),
.Y(n_9565)
);

INVx1_ASAP7_75t_L g9566 ( 
.A(n_8089),
.Y(n_9566)
);

CKINVDCx6p67_ASAP7_75t_R g9567 ( 
.A(n_7821),
.Y(n_9567)
);

AOI22xp33_ASAP7_75t_L g9568 ( 
.A1(n_8136),
.A2(n_6776),
.B1(n_6737),
.B2(n_7485),
.Y(n_9568)
);

AOI22xp33_ASAP7_75t_SL g9569 ( 
.A1(n_8109),
.A2(n_7615),
.B1(n_7701),
.B2(n_7603),
.Y(n_9569)
);

HB1xp67_ASAP7_75t_L g9570 ( 
.A(n_8111),
.Y(n_9570)
);

BUFx3_ASAP7_75t_L g9571 ( 
.A(n_8024),
.Y(n_9571)
);

INVxp67_ASAP7_75t_SL g9572 ( 
.A(n_8313),
.Y(n_9572)
);

INVx1_ASAP7_75t_L g9573 ( 
.A(n_8102),
.Y(n_9573)
);

BUFx3_ASAP7_75t_L g9574 ( 
.A(n_8024),
.Y(n_9574)
);

INVx1_ASAP7_75t_L g9575 ( 
.A(n_8102),
.Y(n_9575)
);

INVx2_ASAP7_75t_L g9576 ( 
.A(n_7720),
.Y(n_9576)
);

INVx2_ASAP7_75t_L g9577 ( 
.A(n_7737),
.Y(n_9577)
);

AOI22xp33_ASAP7_75t_SL g9578 ( 
.A1(n_8164),
.A2(n_7615),
.B1(n_7603),
.B2(n_7261),
.Y(n_9578)
);

OAI22xp33_ASAP7_75t_L g9579 ( 
.A1(n_8195),
.A2(n_7556),
.B1(n_7554),
.B2(n_7519),
.Y(n_9579)
);

INVx1_ASAP7_75t_L g9580 ( 
.A(n_8108),
.Y(n_9580)
);

CKINVDCx5p33_ASAP7_75t_R g9581 ( 
.A(n_7983),
.Y(n_9581)
);

AOI21x1_ASAP7_75t_L g9582 ( 
.A1(n_8614),
.A2(n_6696),
.B(n_6687),
.Y(n_9582)
);

INVx1_ASAP7_75t_L g9583 ( 
.A(n_8108),
.Y(n_9583)
);

INVx6_ASAP7_75t_L g9584 ( 
.A(n_7850),
.Y(n_9584)
);

OAI21xp5_ASAP7_75t_L g9585 ( 
.A1(n_7970),
.A2(n_7699),
.B(n_7513),
.Y(n_9585)
);

BUFx8_ASAP7_75t_SL g9586 ( 
.A(n_8546),
.Y(n_9586)
);

BUFx3_ASAP7_75t_L g9587 ( 
.A(n_8024),
.Y(n_9587)
);

INVx1_ASAP7_75t_L g9588 ( 
.A(n_8112),
.Y(n_9588)
);

INVx2_ASAP7_75t_L g9589 ( 
.A(n_7737),
.Y(n_9589)
);

AND2x4_ASAP7_75t_L g9590 ( 
.A(n_8859),
.B(n_6971),
.Y(n_9590)
);

INVx5_ASAP7_75t_L g9591 ( 
.A(n_8044),
.Y(n_9591)
);

INVx2_ASAP7_75t_L g9592 ( 
.A(n_7737),
.Y(n_9592)
);

AOI21x1_ASAP7_75t_L g9593 ( 
.A1(n_8614),
.A2(n_6696),
.B(n_6687),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_7745),
.Y(n_9594)
);

INVx1_ASAP7_75t_L g9595 ( 
.A(n_8112),
.Y(n_9595)
);

HB1xp67_ASAP7_75t_L g9596 ( 
.A(n_8111),
.Y(n_9596)
);

NAND2xp5_ASAP7_75t_L g9597 ( 
.A(n_8815),
.B(n_7233),
.Y(n_9597)
);

INVx2_ASAP7_75t_L g9598 ( 
.A(n_7745),
.Y(n_9598)
);

AOI22xp33_ASAP7_75t_L g9599 ( 
.A1(n_8944),
.A2(n_6776),
.B1(n_6737),
.B2(n_7494),
.Y(n_9599)
);

INVx2_ASAP7_75t_L g9600 ( 
.A(n_7745),
.Y(n_9600)
);

BUFx8_ASAP7_75t_L g9601 ( 
.A(n_8239),
.Y(n_9601)
);

INVx4_ASAP7_75t_L g9602 ( 
.A(n_8912),
.Y(n_9602)
);

CKINVDCx5p33_ASAP7_75t_R g9603 ( 
.A(n_8003),
.Y(n_9603)
);

BUFx6f_ASAP7_75t_L g9604 ( 
.A(n_8044),
.Y(n_9604)
);

INVx2_ASAP7_75t_L g9605 ( 
.A(n_7777),
.Y(n_9605)
);

INVx2_ASAP7_75t_L g9606 ( 
.A(n_7777),
.Y(n_9606)
);

INVx1_ASAP7_75t_L g9607 ( 
.A(n_8124),
.Y(n_9607)
);

INVxp67_ASAP7_75t_SL g9608 ( 
.A(n_8551),
.Y(n_9608)
);

BUFx2_ASAP7_75t_L g9609 ( 
.A(n_8742),
.Y(n_9609)
);

INVx2_ASAP7_75t_L g9610 ( 
.A(n_7777),
.Y(n_9610)
);

INVx1_ASAP7_75t_L g9611 ( 
.A(n_8124),
.Y(n_9611)
);

INVx3_ASAP7_75t_L g9612 ( 
.A(n_8044),
.Y(n_9612)
);

AO21x1_ASAP7_75t_L g9613 ( 
.A1(n_8972),
.A2(n_7328),
.B(n_7284),
.Y(n_9613)
);

INVx2_ASAP7_75t_L g9614 ( 
.A(n_7789),
.Y(n_9614)
);

NAND2xp5_ASAP7_75t_L g9615 ( 
.A(n_8906),
.B(n_8917),
.Y(n_9615)
);

HB1xp67_ASAP7_75t_L g9616 ( 
.A(n_8170),
.Y(n_9616)
);

INVx1_ASAP7_75t_L g9617 ( 
.A(n_8129),
.Y(n_9617)
);

HB1xp67_ASAP7_75t_L g9618 ( 
.A(n_8170),
.Y(n_9618)
);

CKINVDCx16_ASAP7_75t_R g9619 ( 
.A(n_8771),
.Y(n_9619)
);

INVx2_ASAP7_75t_L g9620 ( 
.A(n_7789),
.Y(n_9620)
);

CKINVDCx20_ASAP7_75t_R g9621 ( 
.A(n_8003),
.Y(n_9621)
);

INVx2_ASAP7_75t_L g9622 ( 
.A(n_7789),
.Y(n_9622)
);

INVx2_ASAP7_75t_SL g9623 ( 
.A(n_8050),
.Y(n_9623)
);

AOI22xp33_ASAP7_75t_SL g9624 ( 
.A1(n_8100),
.A2(n_7615),
.B1(n_7603),
.B2(n_7261),
.Y(n_9624)
);

AND2x4_ASAP7_75t_L g9625 ( 
.A(n_8933),
.B(n_6971),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_8129),
.Y(n_9626)
);

AND2x2_ASAP7_75t_L g9627 ( 
.A(n_8104),
.B(n_8115),
.Y(n_9627)
);

BUFx3_ASAP7_75t_L g9628 ( 
.A(n_8024),
.Y(n_9628)
);

HB1xp67_ASAP7_75t_L g9629 ( 
.A(n_8226),
.Y(n_9629)
);

INVx3_ASAP7_75t_L g9630 ( 
.A(n_8044),
.Y(n_9630)
);

AOI22xp33_ASAP7_75t_SL g9631 ( 
.A1(n_8100),
.A2(n_7603),
.B1(n_7261),
.B2(n_7321),
.Y(n_9631)
);

INVx1_ASAP7_75t_L g9632 ( 
.A(n_8131),
.Y(n_9632)
);

INVx1_ASAP7_75t_SL g9633 ( 
.A(n_8096),
.Y(n_9633)
);

CKINVDCx20_ASAP7_75t_R g9634 ( 
.A(n_8067),
.Y(n_9634)
);

INVx2_ASAP7_75t_L g9635 ( 
.A(n_7800),
.Y(n_9635)
);

INVx2_ASAP7_75t_L g9636 ( 
.A(n_7800),
.Y(n_9636)
);

INVx4_ASAP7_75t_L g9637 ( 
.A(n_8912),
.Y(n_9637)
);

INVx1_ASAP7_75t_L g9638 ( 
.A(n_8131),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_8138),
.Y(n_9639)
);

INVx1_ASAP7_75t_L g9640 ( 
.A(n_8138),
.Y(n_9640)
);

OAI21x1_ASAP7_75t_L g9641 ( 
.A1(n_8346),
.A2(n_6924),
.B(n_6872),
.Y(n_9641)
);

AND2x2_ASAP7_75t_L g9642 ( 
.A(n_8104),
.B(n_6971),
.Y(n_9642)
);

OAI21xp5_ASAP7_75t_L g9643 ( 
.A1(n_8211),
.A2(n_7699),
.B(n_7513),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_8155),
.Y(n_9644)
);

AOI22xp33_ASAP7_75t_L g9645 ( 
.A1(n_8944),
.A2(n_6776),
.B1(n_6737),
.B2(n_7494),
.Y(n_9645)
);

AND2x2_ASAP7_75t_L g9646 ( 
.A(n_8104),
.B(n_7001),
.Y(n_9646)
);

OAI22xp5_ASAP7_75t_L g9647 ( 
.A1(n_8768),
.A2(n_7447),
.B1(n_7463),
.B2(n_7456),
.Y(n_9647)
);

INVx1_ASAP7_75t_L g9648 ( 
.A(n_8155),
.Y(n_9648)
);

AOI22xp33_ASAP7_75t_L g9649 ( 
.A1(n_8147),
.A2(n_6776),
.B1(n_6737),
.B2(n_7103),
.Y(n_9649)
);

BUFx3_ASAP7_75t_L g9650 ( 
.A(n_8024),
.Y(n_9650)
);

OAI21x1_ASAP7_75t_L g9651 ( 
.A1(n_8907),
.A2(n_7446),
.B(n_6924),
.Y(n_9651)
);

AOI22xp5_ASAP7_75t_L g9652 ( 
.A1(n_7932),
.A2(n_7540),
.B1(n_7281),
.B2(n_7151),
.Y(n_9652)
);

OAI21x1_ASAP7_75t_L g9653 ( 
.A1(n_8941),
.A2(n_7446),
.B(n_6924),
.Y(n_9653)
);

INVx1_ASAP7_75t_L g9654 ( 
.A(n_8157),
.Y(n_9654)
);

OA21x2_ASAP7_75t_L g9655 ( 
.A1(n_8029),
.A2(n_6822),
.B(n_7284),
.Y(n_9655)
);

INVx2_ASAP7_75t_SL g9656 ( 
.A(n_8362),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_8157),
.Y(n_9657)
);

AOI21x1_ASAP7_75t_L g9658 ( 
.A1(n_8682),
.A2(n_6711),
.B(n_6708),
.Y(n_9658)
);

INVx1_ASAP7_75t_L g9659 ( 
.A(n_8159),
.Y(n_9659)
);

INVx4_ASAP7_75t_L g9660 ( 
.A(n_8024),
.Y(n_9660)
);

AOI22xp5_ASAP7_75t_L g9661 ( 
.A1(n_7932),
.A2(n_7540),
.B1(n_7103),
.B2(n_7161),
.Y(n_9661)
);

HB1xp67_ASAP7_75t_L g9662 ( 
.A(n_8226),
.Y(n_9662)
);

OAI21x1_ASAP7_75t_L g9663 ( 
.A1(n_8632),
.A2(n_6924),
.B(n_6872),
.Y(n_9663)
);

INVx2_ASAP7_75t_L g9664 ( 
.A(n_7800),
.Y(n_9664)
);

INVx2_ASAP7_75t_L g9665 ( 
.A(n_7809),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8159),
.Y(n_9666)
);

HB1xp67_ASAP7_75t_L g9667 ( 
.A(n_8273),
.Y(n_9667)
);

OAI22xp5_ASAP7_75t_L g9668 ( 
.A1(n_7950),
.A2(n_7456),
.B1(n_7463),
.B2(n_7478),
.Y(n_9668)
);

BUFx3_ASAP7_75t_L g9669 ( 
.A(n_8386),
.Y(n_9669)
);

INVx1_ASAP7_75t_L g9670 ( 
.A(n_8174),
.Y(n_9670)
);

AND2x2_ASAP7_75t_L g9671 ( 
.A(n_8115),
.B(n_7001),
.Y(n_9671)
);

INVx6_ASAP7_75t_L g9672 ( 
.A(n_7850),
.Y(n_9672)
);

INVx1_ASAP7_75t_L g9673 ( 
.A(n_8174),
.Y(n_9673)
);

CKINVDCx11_ASAP7_75t_R g9674 ( 
.A(n_8067),
.Y(n_9674)
);

INVx6_ASAP7_75t_L g9675 ( 
.A(n_7850),
.Y(n_9675)
);

INVx1_ASAP7_75t_L g9676 ( 
.A(n_8203),
.Y(n_9676)
);

NAND2x1p5_ASAP7_75t_L g9677 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9677)
);

BUFx10_ASAP7_75t_L g9678 ( 
.A(n_8158),
.Y(n_9678)
);

INVx8_ASAP7_75t_L g9679 ( 
.A(n_8386),
.Y(n_9679)
);

BUFx3_ASAP7_75t_L g9680 ( 
.A(n_8386),
.Y(n_9680)
);

BUFx6f_ASAP7_75t_L g9681 ( 
.A(n_8044),
.Y(n_9681)
);

HB1xp67_ASAP7_75t_L g9682 ( 
.A(n_8273),
.Y(n_9682)
);

AOI22xp33_ASAP7_75t_SL g9683 ( 
.A1(n_8100),
.A2(n_7603),
.B1(n_7261),
.B2(n_7321),
.Y(n_9683)
);

NAND2xp5_ASAP7_75t_L g9684 ( 
.A(n_8906),
.B(n_7233),
.Y(n_9684)
);

OAI21xp5_ASAP7_75t_L g9685 ( 
.A1(n_8211),
.A2(n_7513),
.B(n_7694),
.Y(n_9685)
);

BUFx3_ASAP7_75t_L g9686 ( 
.A(n_8386),
.Y(n_9686)
);

INVx1_ASAP7_75t_L g9687 ( 
.A(n_8203),
.Y(n_9687)
);

AND2x2_ASAP7_75t_L g9688 ( 
.A(n_8115),
.B(n_7001),
.Y(n_9688)
);

AOI22xp33_ASAP7_75t_SL g9689 ( 
.A1(n_8100),
.A2(n_7603),
.B1(n_7261),
.B2(n_7321),
.Y(n_9689)
);

BUFx2_ASAP7_75t_R g9690 ( 
.A(n_8231),
.Y(n_9690)
);

OAI21x1_ASAP7_75t_L g9691 ( 
.A1(n_8632),
.A2(n_6924),
.B(n_6872),
.Y(n_9691)
);

INVx1_ASAP7_75t_L g9692 ( 
.A(n_8209),
.Y(n_9692)
);

AOI22xp33_ASAP7_75t_L g9693 ( 
.A1(n_8147),
.A2(n_7337),
.B1(n_7314),
.B2(n_7205),
.Y(n_9693)
);

INVx2_ASAP7_75t_L g9694 ( 
.A(n_7809),
.Y(n_9694)
);

NAND2xp5_ASAP7_75t_L g9695 ( 
.A(n_8917),
.B(n_6767),
.Y(n_9695)
);

INVx1_ASAP7_75t_L g9696 ( 
.A(n_8209),
.Y(n_9696)
);

INVx2_ASAP7_75t_L g9697 ( 
.A(n_7809),
.Y(n_9697)
);

INVx2_ASAP7_75t_L g9698 ( 
.A(n_7831),
.Y(n_9698)
);

INVx1_ASAP7_75t_SL g9699 ( 
.A(n_8096),
.Y(n_9699)
);

OAI22xp5_ASAP7_75t_L g9700 ( 
.A1(n_7999),
.A2(n_7478),
.B1(n_7694),
.B2(n_7537),
.Y(n_9700)
);

INVx1_ASAP7_75t_L g9701 ( 
.A(n_8210),
.Y(n_9701)
);

CKINVDCx6p67_ASAP7_75t_R g9702 ( 
.A(n_7821),
.Y(n_9702)
);

CKINVDCx20_ASAP7_75t_R g9703 ( 
.A(n_8308),
.Y(n_9703)
);

INVx2_ASAP7_75t_L g9704 ( 
.A(n_7831),
.Y(n_9704)
);

INVx1_ASAP7_75t_L g9705 ( 
.A(n_8210),
.Y(n_9705)
);

NOR2xp33_ASAP7_75t_L g9706 ( 
.A(n_8957),
.B(n_7396),
.Y(n_9706)
);

INVx2_ASAP7_75t_L g9707 ( 
.A(n_7831),
.Y(n_9707)
);

BUFx6f_ASAP7_75t_L g9708 ( 
.A(n_8082),
.Y(n_9708)
);

INVx1_ASAP7_75t_SL g9709 ( 
.A(n_8135),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_8216),
.Y(n_9710)
);

NOR2xp33_ASAP7_75t_L g9711 ( 
.A(n_8992),
.B(n_7396),
.Y(n_9711)
);

BUFx3_ASAP7_75t_L g9712 ( 
.A(n_8386),
.Y(n_9712)
);

BUFx2_ASAP7_75t_SL g9713 ( 
.A(n_8538),
.Y(n_9713)
);

CKINVDCx20_ASAP7_75t_R g9714 ( 
.A(n_8308),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_8216),
.Y(n_9715)
);

INVx1_ASAP7_75t_L g9716 ( 
.A(n_8255),
.Y(n_9716)
);

AND2x2_ASAP7_75t_L g9717 ( 
.A(n_7864),
.B(n_7001),
.Y(n_9717)
);

BUFx10_ASAP7_75t_L g9718 ( 
.A(n_8926),
.Y(n_9718)
);

HB1xp67_ASAP7_75t_L g9719 ( 
.A(n_8347),
.Y(n_9719)
);

OAI21xp5_ASAP7_75t_SL g9720 ( 
.A1(n_7788),
.A2(n_7339),
.B(n_7554),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_8255),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_8260),
.Y(n_9722)
);

BUFx4f_ASAP7_75t_SL g9723 ( 
.A(n_8573),
.Y(n_9723)
);

OAI21x1_ASAP7_75t_L g9724 ( 
.A1(n_8632),
.A2(n_6984),
.B(n_6924),
.Y(n_9724)
);

BUFx2_ASAP7_75t_L g9725 ( 
.A(n_8742),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_8260),
.Y(n_9726)
);

AND2x2_ASAP7_75t_L g9727 ( 
.A(n_7864),
.B(n_7880),
.Y(n_9727)
);

OAI21x1_ASAP7_75t_L g9728 ( 
.A1(n_8697),
.A2(n_6986),
.B(n_6984),
.Y(n_9728)
);

AND2x2_ASAP7_75t_L g9729 ( 
.A(n_7864),
.B(n_7020),
.Y(n_9729)
);

BUFx6f_ASAP7_75t_L g9730 ( 
.A(n_8082),
.Y(n_9730)
);

AOI22xp33_ASAP7_75t_L g9731 ( 
.A1(n_7943),
.A2(n_7337),
.B1(n_7314),
.B2(n_7205),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_8265),
.Y(n_9732)
);

AOI22xp33_ASAP7_75t_L g9733 ( 
.A1(n_7943),
.A2(n_7314),
.B1(n_7205),
.B2(n_7261),
.Y(n_9733)
);

INVx2_ASAP7_75t_L g9734 ( 
.A(n_7839),
.Y(n_9734)
);

AO21x1_ASAP7_75t_L g9735 ( 
.A1(n_8218),
.A2(n_7328),
.B(n_7609),
.Y(n_9735)
);

AOI22xp33_ASAP7_75t_L g9736 ( 
.A1(n_8426),
.A2(n_7314),
.B1(n_7205),
.B2(n_7167),
.Y(n_9736)
);

INVx1_ASAP7_75t_L g9737 ( 
.A(n_8265),
.Y(n_9737)
);

INVx1_ASAP7_75t_L g9738 ( 
.A(n_8267),
.Y(n_9738)
);

AOI22xp33_ASAP7_75t_L g9739 ( 
.A1(n_8426),
.A2(n_7314),
.B1(n_7205),
.B2(n_7167),
.Y(n_9739)
);

INVx1_ASAP7_75t_L g9740 ( 
.A(n_8267),
.Y(n_9740)
);

INVxp67_ASAP7_75t_SL g9741 ( 
.A(n_8551),
.Y(n_9741)
);

INVx2_ASAP7_75t_L g9742 ( 
.A(n_7839),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_7839),
.Y(n_9743)
);

OAI21xp5_ASAP7_75t_SL g9744 ( 
.A1(n_7788),
.A2(n_7556),
.B(n_7537),
.Y(n_9744)
);

INVx2_ASAP7_75t_SL g9745 ( 
.A(n_8362),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_8269),
.Y(n_9746)
);

INVx2_ASAP7_75t_L g9747 ( 
.A(n_7853),
.Y(n_9747)
);

AO21x2_ASAP7_75t_L g9748 ( 
.A1(n_8739),
.A2(n_8047),
.B(n_7988),
.Y(n_9748)
);

INVx2_ASAP7_75t_L g9749 ( 
.A(n_7853),
.Y(n_9749)
);

OAI22xp5_ASAP7_75t_L g9750 ( 
.A1(n_7999),
.A2(n_7542),
.B1(n_7599),
.B2(n_7574),
.Y(n_9750)
);

INVx2_ASAP7_75t_SL g9751 ( 
.A(n_8362),
.Y(n_9751)
);

BUFx6f_ASAP7_75t_L g9752 ( 
.A(n_8082),
.Y(n_9752)
);

OA21x2_ASAP7_75t_L g9753 ( 
.A1(n_8033),
.A2(n_7718),
.B(n_8685),
.Y(n_9753)
);

BUFx6f_ASAP7_75t_L g9754 ( 
.A(n_8082),
.Y(n_9754)
);

NOR2xp33_ASAP7_75t_L g9755 ( 
.A(n_8992),
.B(n_7396),
.Y(n_9755)
);

INVx2_ASAP7_75t_L g9756 ( 
.A(n_7853),
.Y(n_9756)
);

AO21x2_ASAP7_75t_L g9757 ( 
.A1(n_8739),
.A2(n_6711),
.B(n_6708),
.Y(n_9757)
);

INVx2_ASAP7_75t_L g9758 ( 
.A(n_7857),
.Y(n_9758)
);

AOI222xp33_ASAP7_75t_L g9759 ( 
.A1(n_8246),
.A2(n_7542),
.B1(n_7516),
.B2(n_7499),
.C1(n_7222),
.C2(n_6825),
.Y(n_9759)
);

INVx2_ASAP7_75t_L g9760 ( 
.A(n_7857),
.Y(n_9760)
);

AOI22xp33_ASAP7_75t_L g9761 ( 
.A1(n_7797),
.A2(n_7314),
.B1(n_7205),
.B2(n_7167),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_8269),
.Y(n_9762)
);

HB1xp67_ASAP7_75t_L g9763 ( 
.A(n_8347),
.Y(n_9763)
);

OR2x6_ASAP7_75t_L g9764 ( 
.A(n_8404),
.B(n_6807),
.Y(n_9764)
);

INVx2_ASAP7_75t_L g9765 ( 
.A(n_7857),
.Y(n_9765)
);

AOI22xp33_ASAP7_75t_SL g9766 ( 
.A1(n_8218),
.A2(n_7603),
.B1(n_7321),
.B2(n_7335),
.Y(n_9766)
);

BUFx8_ASAP7_75t_SL g9767 ( 
.A(n_8573),
.Y(n_9767)
);

BUFx6f_ASAP7_75t_L g9768 ( 
.A(n_8082),
.Y(n_9768)
);

AOI22xp33_ASAP7_75t_L g9769 ( 
.A1(n_7797),
.A2(n_7314),
.B1(n_7205),
.B2(n_7167),
.Y(n_9769)
);

AOI21xp5_ASAP7_75t_L g9770 ( 
.A1(n_8047),
.A2(n_7430),
.B(n_7609),
.Y(n_9770)
);

HB1xp67_ASAP7_75t_L g9771 ( 
.A(n_8367),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_8283),
.Y(n_9772)
);

INVx2_ASAP7_75t_L g9773 ( 
.A(n_7910),
.Y(n_9773)
);

CKINVDCx20_ASAP7_75t_R g9774 ( 
.A(n_8692),
.Y(n_9774)
);

INVx1_ASAP7_75t_L g9775 ( 
.A(n_8283),
.Y(n_9775)
);

HB1xp67_ASAP7_75t_L g9776 ( 
.A(n_8367),
.Y(n_9776)
);

INVx8_ASAP7_75t_L g9777 ( 
.A(n_8386),
.Y(n_9777)
);

INVx2_ASAP7_75t_L g9778 ( 
.A(n_7910),
.Y(n_9778)
);

BUFx3_ASAP7_75t_L g9779 ( 
.A(n_8386),
.Y(n_9779)
);

INVx2_ASAP7_75t_L g9780 ( 
.A(n_7910),
.Y(n_9780)
);

OAI21x1_ASAP7_75t_L g9781 ( 
.A1(n_8697),
.A2(n_6986),
.B(n_6984),
.Y(n_9781)
);

INVx2_ASAP7_75t_L g9782 ( 
.A(n_7919),
.Y(n_9782)
);

INVx1_ASAP7_75t_L g9783 ( 
.A(n_8291),
.Y(n_9783)
);

NAND2xp5_ASAP7_75t_L g9784 ( 
.A(n_9011),
.B(n_6767),
.Y(n_9784)
);

INVx1_ASAP7_75t_L g9785 ( 
.A(n_8291),
.Y(n_9785)
);

AOI22xp33_ASAP7_75t_L g9786 ( 
.A1(n_7927),
.A2(n_7314),
.B1(n_7205),
.B2(n_7167),
.Y(n_9786)
);

INVx1_ASAP7_75t_L g9787 ( 
.A(n_8297),
.Y(n_9787)
);

AOI22xp33_ASAP7_75t_L g9788 ( 
.A1(n_7927),
.A2(n_8246),
.B1(n_8130),
.B2(n_8149),
.Y(n_9788)
);

AOI22xp5_ASAP7_75t_L g9789 ( 
.A1(n_7928),
.A2(n_7161),
.B1(n_7365),
.B2(n_7556),
.Y(n_9789)
);

BUFx2_ASAP7_75t_R g9790 ( 
.A(n_8711),
.Y(n_9790)
);

INVx2_ASAP7_75t_L g9791 ( 
.A(n_7919),
.Y(n_9791)
);

INVx1_ASAP7_75t_L g9792 ( 
.A(n_8297),
.Y(n_9792)
);

OAI21x1_ASAP7_75t_L g9793 ( 
.A1(n_8697),
.A2(n_6986),
.B(n_6984),
.Y(n_9793)
);

AOI22xp5_ASAP7_75t_L g9794 ( 
.A1(n_7928),
.A2(n_7365),
.B1(n_7599),
.B2(n_7574),
.Y(n_9794)
);

OAI22xp5_ASAP7_75t_L g9795 ( 
.A1(n_8139),
.A2(n_7599),
.B1(n_7574),
.B2(n_7516),
.Y(n_9795)
);

CKINVDCx5p33_ASAP7_75t_R g9796 ( 
.A(n_8692),
.Y(n_9796)
);

BUFx3_ASAP7_75t_L g9797 ( 
.A(n_8429),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_8303),
.Y(n_9798)
);

INVx1_ASAP7_75t_L g9799 ( 
.A(n_8303),
.Y(n_9799)
);

INVx1_ASAP7_75t_L g9800 ( 
.A(n_8306),
.Y(n_9800)
);

INVx4_ASAP7_75t_L g9801 ( 
.A(n_8429),
.Y(n_9801)
);

INVx2_ASAP7_75t_L g9802 ( 
.A(n_7919),
.Y(n_9802)
);

OAI22xp33_ASAP7_75t_L g9803 ( 
.A1(n_8117),
.A2(n_7502),
.B1(n_7529),
.B2(n_7519),
.Y(n_9803)
);

INVx3_ASAP7_75t_L g9804 ( 
.A(n_8082),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_9011),
.B(n_6825),
.Y(n_9805)
);

INVx1_ASAP7_75t_L g9806 ( 
.A(n_8306),
.Y(n_9806)
);

OAI22xp5_ASAP7_75t_L g9807 ( 
.A1(n_8139),
.A2(n_7499),
.B1(n_7222),
.B2(n_7660),
.Y(n_9807)
);

OA21x2_ASAP7_75t_L g9808 ( 
.A1(n_8033),
.A2(n_6711),
.B(n_6708),
.Y(n_9808)
);

HB1xp67_ASAP7_75t_L g9809 ( 
.A(n_8376),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_8307),
.Y(n_9810)
);

OAI21x1_ASAP7_75t_L g9811 ( 
.A1(n_8697),
.A2(n_6986),
.B(n_6984),
.Y(n_9811)
);

BUFx2_ASAP7_75t_L g9812 ( 
.A(n_8742),
.Y(n_9812)
);

INVx4_ASAP7_75t_L g9813 ( 
.A(n_8429),
.Y(n_9813)
);

NAND2x1p5_ASAP7_75t_L g9814 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_8307),
.Y(n_9815)
);

BUFx3_ASAP7_75t_L g9816 ( 
.A(n_8429),
.Y(n_9816)
);

INVx1_ASAP7_75t_L g9817 ( 
.A(n_8309),
.Y(n_9817)
);

INVx2_ASAP7_75t_L g9818 ( 
.A(n_7936),
.Y(n_9818)
);

HB1xp67_ASAP7_75t_L g9819 ( 
.A(n_8376),
.Y(n_9819)
);

CKINVDCx11_ASAP7_75t_R g9820 ( 
.A(n_8788),
.Y(n_9820)
);

INVx2_ASAP7_75t_L g9821 ( 
.A(n_7936),
.Y(n_9821)
);

HB1xp67_ASAP7_75t_L g9822 ( 
.A(n_8392),
.Y(n_9822)
);

AOI22xp33_ASAP7_75t_SL g9823 ( 
.A1(n_8394),
.A2(n_7603),
.B1(n_7321),
.B2(n_7335),
.Y(n_9823)
);

INVx2_ASAP7_75t_L g9824 ( 
.A(n_7936),
.Y(n_9824)
);

INVx2_ASAP7_75t_L g9825 ( 
.A(n_7940),
.Y(n_9825)
);

INVx1_ASAP7_75t_L g9826 ( 
.A(n_8309),
.Y(n_9826)
);

NAND2x1_ASAP7_75t_L g9827 ( 
.A(n_7988),
.B(n_7278),
.Y(n_9827)
);

NAND2xp5_ASAP7_75t_L g9828 ( 
.A(n_9012),
.B(n_7236),
.Y(n_9828)
);

AOI22xp33_ASAP7_75t_L g9829 ( 
.A1(n_8130),
.A2(n_7321),
.B1(n_7335),
.B2(n_7167),
.Y(n_9829)
);

NAND2xp5_ASAP7_75t_L g9830 ( 
.A(n_9012),
.B(n_7236),
.Y(n_9830)
);

BUFx2_ASAP7_75t_L g9831 ( 
.A(n_7939),
.Y(n_9831)
);

INVx1_ASAP7_75t_L g9832 ( 
.A(n_8310),
.Y(n_9832)
);

INVx1_ASAP7_75t_L g9833 ( 
.A(n_8310),
.Y(n_9833)
);

AOI22xp33_ASAP7_75t_L g9834 ( 
.A1(n_8149),
.A2(n_7360),
.B1(n_7438),
.B2(n_7335),
.Y(n_9834)
);

AO21x2_ASAP7_75t_L g9835 ( 
.A1(n_8739),
.A2(n_6653),
.B(n_6652),
.Y(n_9835)
);

AO21x2_ASAP7_75t_L g9836 ( 
.A1(n_8739),
.A2(n_6653),
.B(n_6652),
.Y(n_9836)
);

OAI22xp33_ASAP7_75t_L g9837 ( 
.A1(n_8066),
.A2(n_7502),
.B1(n_7529),
.B2(n_7400),
.Y(n_9837)
);

INVx1_ASAP7_75t_L g9838 ( 
.A(n_8314),
.Y(n_9838)
);

INVx2_ASAP7_75t_L g9839 ( 
.A(n_7940),
.Y(n_9839)
);

BUFx2_ASAP7_75t_L g9840 ( 
.A(n_8160),
.Y(n_9840)
);

INVx2_ASAP7_75t_L g9841 ( 
.A(n_7940),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_8314),
.Y(n_9842)
);

INVx1_ASAP7_75t_L g9843 ( 
.A(n_8333),
.Y(n_9843)
);

AOI21xp5_ASAP7_75t_L g9844 ( 
.A1(n_7744),
.A2(n_7664),
.B(n_7497),
.Y(n_9844)
);

AND2x2_ASAP7_75t_L g9845 ( 
.A(n_7880),
.B(n_7020),
.Y(n_9845)
);

AND2x2_ASAP7_75t_L g9846 ( 
.A(n_7880),
.B(n_7020),
.Y(n_9846)
);

CKINVDCx11_ASAP7_75t_R g9847 ( 
.A(n_8788),
.Y(n_9847)
);

AOI22xp33_ASAP7_75t_L g9848 ( 
.A1(n_8691),
.A2(n_7360),
.B1(n_7438),
.B2(n_7335),
.Y(n_9848)
);

INVx2_ASAP7_75t_L g9849 ( 
.A(n_7949),
.Y(n_9849)
);

AND2x2_ASAP7_75t_L g9850 ( 
.A(n_8002),
.B(n_7020),
.Y(n_9850)
);

BUFx3_ASAP7_75t_L g9851 ( 
.A(n_8429),
.Y(n_9851)
);

INVx1_ASAP7_75t_L g9852 ( 
.A(n_8333),
.Y(n_9852)
);

AOI22xp33_ASAP7_75t_L g9853 ( 
.A1(n_8691),
.A2(n_7360),
.B1(n_7438),
.B2(n_7335),
.Y(n_9853)
);

INVx2_ASAP7_75t_L g9854 ( 
.A(n_7949),
.Y(n_9854)
);

INVx1_ASAP7_75t_L g9855 ( 
.A(n_8339),
.Y(n_9855)
);

INVxp67_ASAP7_75t_SL g9856 ( 
.A(n_8551),
.Y(n_9856)
);

INVx1_ASAP7_75t_L g9857 ( 
.A(n_8339),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_L g9858 ( 
.A(n_7907),
.B(n_7241),
.Y(n_9858)
);

HB1xp67_ASAP7_75t_L g9859 ( 
.A(n_8392),
.Y(n_9859)
);

CKINVDCx11_ASAP7_75t_R g9860 ( 
.A(n_8818),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_8341),
.Y(n_9861)
);

OA21x2_ASAP7_75t_L g9862 ( 
.A1(n_8033),
.A2(n_6667),
.B(n_6659),
.Y(n_9862)
);

AND2x4_ASAP7_75t_L g9863 ( 
.A(n_8933),
.B(n_7023),
.Y(n_9863)
);

AO21x2_ASAP7_75t_L g9864 ( 
.A1(n_7988),
.A2(n_6653),
.B(n_6652),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_8341),
.Y(n_9865)
);

OAI21x1_ASAP7_75t_L g9866 ( 
.A1(n_8814),
.A2(n_6986),
.B(n_6984),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_8343),
.Y(n_9867)
);

BUFx2_ASAP7_75t_L g9868 ( 
.A(n_8208),
.Y(n_9868)
);

AOI22xp33_ASAP7_75t_SL g9869 ( 
.A1(n_8394),
.A2(n_7603),
.B1(n_7360),
.B2(n_7460),
.Y(n_9869)
);

INVx1_ASAP7_75t_L g9870 ( 
.A(n_8343),
.Y(n_9870)
);

INVx1_ASAP7_75t_L g9871 ( 
.A(n_8345),
.Y(n_9871)
);

INVx1_ASAP7_75t_L g9872 ( 
.A(n_8345),
.Y(n_9872)
);

CKINVDCx20_ASAP7_75t_R g9873 ( 
.A(n_8818),
.Y(n_9873)
);

BUFx6f_ASAP7_75t_L g9874 ( 
.A(n_8082),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_8348),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_8348),
.Y(n_9876)
);

NAND2x1p5_ASAP7_75t_L g9877 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9877)
);

HB1xp67_ASAP7_75t_L g9878 ( 
.A(n_8464),
.Y(n_9878)
);

INVx1_ASAP7_75t_L g9879 ( 
.A(n_8360),
.Y(n_9879)
);

CKINVDCx5p33_ASAP7_75t_R g9880 ( 
.A(n_8723),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_8360),
.Y(n_9881)
);

INVx2_ASAP7_75t_L g9882 ( 
.A(n_7949),
.Y(n_9882)
);

INVx2_ASAP7_75t_L g9883 ( 
.A(n_7962),
.Y(n_9883)
);

INVx3_ASAP7_75t_L g9884 ( 
.A(n_8082),
.Y(n_9884)
);

INVx1_ASAP7_75t_L g9885 ( 
.A(n_8363),
.Y(n_9885)
);

AND2x2_ASAP7_75t_L g9886 ( 
.A(n_8002),
.B(n_7023),
.Y(n_9886)
);

INVx3_ASAP7_75t_L g9887 ( 
.A(n_8114),
.Y(n_9887)
);

AND2x2_ASAP7_75t_L g9888 ( 
.A(n_8002),
.B(n_8144),
.Y(n_9888)
);

HB1xp67_ASAP7_75t_L g9889 ( 
.A(n_8464),
.Y(n_9889)
);

BUFx2_ASAP7_75t_L g9890 ( 
.A(n_7939),
.Y(n_9890)
);

AOI21xp5_ASAP7_75t_L g9891 ( 
.A1(n_7744),
.A2(n_7664),
.B(n_7497),
.Y(n_9891)
);

INVx2_ASAP7_75t_L g9892 ( 
.A(n_7962),
.Y(n_9892)
);

AOI22xp33_ASAP7_75t_SL g9893 ( 
.A1(n_7930),
.A2(n_7984),
.B1(n_8070),
.B2(n_8414),
.Y(n_9893)
);

INVx2_ASAP7_75t_L g9894 ( 
.A(n_7962),
.Y(n_9894)
);

AND2x4_ASAP7_75t_L g9895 ( 
.A(n_8933),
.B(n_7023),
.Y(n_9895)
);

INVx2_ASAP7_75t_L g9896 ( 
.A(n_7969),
.Y(n_9896)
);

AND2x4_ASAP7_75t_L g9897 ( 
.A(n_8940),
.B(n_7023),
.Y(n_9897)
);

AOI22xp5_ASAP7_75t_L g9898 ( 
.A1(n_8172),
.A2(n_7635),
.B1(n_7613),
.B2(n_7400),
.Y(n_9898)
);

HB1xp67_ASAP7_75t_L g9899 ( 
.A(n_8540),
.Y(n_9899)
);

HB1xp67_ASAP7_75t_L g9900 ( 
.A(n_8540),
.Y(n_9900)
);

INVx1_ASAP7_75t_L g9901 ( 
.A(n_8363),
.Y(n_9901)
);

BUFx3_ASAP7_75t_L g9902 ( 
.A(n_8429),
.Y(n_9902)
);

INVx4_ASAP7_75t_L g9903 ( 
.A(n_8429),
.Y(n_9903)
);

HB1xp67_ASAP7_75t_L g9904 ( 
.A(n_8660),
.Y(n_9904)
);

OAI21x1_ASAP7_75t_L g9905 ( 
.A1(n_8941),
.A2(n_7446),
.B(n_7027),
.Y(n_9905)
);

AOI22xp33_ASAP7_75t_SL g9906 ( 
.A1(n_7930),
.A2(n_7603),
.B1(n_7360),
.B2(n_7460),
.Y(n_9906)
);

NAND2xp5_ASAP7_75t_L g9907 ( 
.A(n_7907),
.B(n_7241),
.Y(n_9907)
);

AOI22xp33_ASAP7_75t_L g9908 ( 
.A1(n_8241),
.A2(n_7438),
.B1(n_7460),
.B2(n_7360),
.Y(n_9908)
);

INVx2_ASAP7_75t_L g9909 ( 
.A(n_7969),
.Y(n_9909)
);

INVx1_ASAP7_75t_L g9910 ( 
.A(n_8374),
.Y(n_9910)
);

INVx2_ASAP7_75t_SL g9911 ( 
.A(n_8362),
.Y(n_9911)
);

INVx2_ASAP7_75t_L g9912 ( 
.A(n_7969),
.Y(n_9912)
);

AOI22xp33_ASAP7_75t_SL g9913 ( 
.A1(n_7984),
.A2(n_7603),
.B1(n_7438),
.B2(n_7460),
.Y(n_9913)
);

INVx2_ASAP7_75t_L g9914 ( 
.A(n_7991),
.Y(n_9914)
);

HB1xp67_ASAP7_75t_L g9915 ( 
.A(n_8660),
.Y(n_9915)
);

BUFx2_ASAP7_75t_L g9916 ( 
.A(n_8208),
.Y(n_9916)
);

BUFx2_ASAP7_75t_L g9917 ( 
.A(n_8208),
.Y(n_9917)
);

AOI22xp33_ASAP7_75t_L g9918 ( 
.A1(n_8241),
.A2(n_7460),
.B1(n_7438),
.B2(n_7613),
.Y(n_9918)
);

INVx3_ASAP7_75t_L g9919 ( 
.A(n_8114),
.Y(n_9919)
);

INVx1_ASAP7_75t_L g9920 ( 
.A(n_8374),
.Y(n_9920)
);

AND2x2_ASAP7_75t_L g9921 ( 
.A(n_8144),
.B(n_7460),
.Y(n_9921)
);

INVx1_ASAP7_75t_L g9922 ( 
.A(n_8380),
.Y(n_9922)
);

INVx1_ASAP7_75t_L g9923 ( 
.A(n_8380),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_8383),
.Y(n_9924)
);

BUFx3_ASAP7_75t_L g9925 ( 
.A(n_8711),
.Y(n_9925)
);

CKINVDCx11_ASAP7_75t_R g9926 ( 
.A(n_8711),
.Y(n_9926)
);

AND2x2_ASAP7_75t_L g9927 ( 
.A(n_8144),
.B(n_6827),
.Y(n_9927)
);

INVx6_ASAP7_75t_L g9928 ( 
.A(n_7850),
.Y(n_9928)
);

INVx1_ASAP7_75t_L g9929 ( 
.A(n_8383),
.Y(n_9929)
);

INVx2_ASAP7_75t_L g9930 ( 
.A(n_7991),
.Y(n_9930)
);

INVx8_ASAP7_75t_L g9931 ( 
.A(n_8965),
.Y(n_9931)
);

INVx2_ASAP7_75t_L g9932 ( 
.A(n_7991),
.Y(n_9932)
);

AND2x4_ASAP7_75t_L g9933 ( 
.A(n_8940),
.B(n_7384),
.Y(n_9933)
);

BUFx2_ASAP7_75t_L g9934 ( 
.A(n_7939),
.Y(n_9934)
);

INVxp33_ASAP7_75t_L g9935 ( 
.A(n_8612),
.Y(n_9935)
);

AOI22xp33_ASAP7_75t_L g9936 ( 
.A1(n_8512),
.A2(n_7635),
.B1(n_5809),
.B2(n_5808),
.Y(n_9936)
);

OAI22xp33_ASAP7_75t_L g9937 ( 
.A1(n_8066),
.A2(n_7529),
.B1(n_7400),
.B2(n_7614),
.Y(n_9937)
);

AOI22xp33_ASAP7_75t_L g9938 ( 
.A1(n_8512),
.A2(n_5809),
.B1(n_5808),
.B2(n_7278),
.Y(n_9938)
);

INVx2_ASAP7_75t_L g9939 ( 
.A(n_8007),
.Y(n_9939)
);

INVx2_ASAP7_75t_L g9940 ( 
.A(n_8007),
.Y(n_9940)
);

AO21x1_ASAP7_75t_L g9941 ( 
.A1(n_8062),
.A2(n_6934),
.B(n_7062),
.Y(n_9941)
);

INVx2_ASAP7_75t_L g9942 ( 
.A(n_8007),
.Y(n_9942)
);

OAI21x1_ASAP7_75t_L g9943 ( 
.A1(n_8681),
.A2(n_7027),
.B(n_6986),
.Y(n_9943)
);

INVx2_ASAP7_75t_L g9944 ( 
.A(n_8013),
.Y(n_9944)
);

AOI22xp33_ASAP7_75t_SL g9945 ( 
.A1(n_7984),
.A2(n_8070),
.B1(n_8452),
.B2(n_8414),
.Y(n_9945)
);

AOI22xp33_ASAP7_75t_L g9946 ( 
.A1(n_8698),
.A2(n_5809),
.B1(n_5808),
.B2(n_5719),
.Y(n_9946)
);

OA21x2_ASAP7_75t_L g9947 ( 
.A1(n_7718),
.A2(n_6667),
.B(n_6659),
.Y(n_9947)
);

AOI22xp33_ASAP7_75t_SL g9948 ( 
.A1(n_7984),
.A2(n_7603),
.B1(n_7590),
.B2(n_7583),
.Y(n_9948)
);

AO21x1_ASAP7_75t_L g9949 ( 
.A1(n_8062),
.A2(n_8452),
.B(n_7963),
.Y(n_9949)
);

INVx4_ASAP7_75t_L g9950 ( 
.A(n_8711),
.Y(n_9950)
);

NAND2x1p5_ASAP7_75t_L g9951 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9951)
);

INVx2_ASAP7_75t_SL g9952 ( 
.A(n_8362),
.Y(n_9952)
);

INVx2_ASAP7_75t_L g9953 ( 
.A(n_8013),
.Y(n_9953)
);

OAI22xp5_ASAP7_75t_L g9954 ( 
.A1(n_7956),
.A2(n_7660),
.B1(n_7392),
.B2(n_7370),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_8387),
.Y(n_9955)
);

BUFx2_ASAP7_75t_L g9956 ( 
.A(n_7939),
.Y(n_9956)
);

INVx2_ASAP7_75t_SL g9957 ( 
.A(n_8362),
.Y(n_9957)
);

INVx1_ASAP7_75t_L g9958 ( 
.A(n_8387),
.Y(n_9958)
);

INVx4_ASAP7_75t_L g9959 ( 
.A(n_8919),
.Y(n_9959)
);

INVx3_ASAP7_75t_L g9960 ( 
.A(n_8114),
.Y(n_9960)
);

INVx1_ASAP7_75t_L g9961 ( 
.A(n_8410),
.Y(n_9961)
);

NAND2x1p5_ASAP7_75t_L g9962 ( 
.A(n_8738),
.B(n_7133),
.Y(n_9962)
);

BUFx6f_ASAP7_75t_L g9963 ( 
.A(n_8114),
.Y(n_9963)
);

INVx2_ASAP7_75t_L g9964 ( 
.A(n_8013),
.Y(n_9964)
);

AND2x4_ASAP7_75t_L g9965 ( 
.A(n_8940),
.B(n_7389),
.Y(n_9965)
);

INVxp67_ASAP7_75t_L g9966 ( 
.A(n_7937),
.Y(n_9966)
);

INVx1_ASAP7_75t_L g9967 ( 
.A(n_8410),
.Y(n_9967)
);

NAND2xp5_ASAP7_75t_L g9968 ( 
.A(n_8361),
.B(n_7283),
.Y(n_9968)
);

INVx2_ASAP7_75t_SL g9969 ( 
.A(n_8820),
.Y(n_9969)
);

INVx1_ASAP7_75t_L g9970 ( 
.A(n_8417),
.Y(n_9970)
);

AOI22xp33_ASAP7_75t_L g9971 ( 
.A1(n_8698),
.A2(n_5809),
.B1(n_5808),
.B2(n_5719),
.Y(n_9971)
);

INVx1_ASAP7_75t_L g9972 ( 
.A(n_8417),
.Y(n_9972)
);

BUFx3_ASAP7_75t_L g9973 ( 
.A(n_8919),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_8432),
.Y(n_9974)
);

INVx2_ASAP7_75t_L g9975 ( 
.A(n_8017),
.Y(n_9975)
);

CKINVDCx5p33_ASAP7_75t_R g9976 ( 
.A(n_8842),
.Y(n_9976)
);

BUFx2_ASAP7_75t_R g9977 ( 
.A(n_8919),
.Y(n_9977)
);

NAND2xp5_ASAP7_75t_L g9978 ( 
.A(n_8361),
.B(n_7283),
.Y(n_9978)
);

AO21x2_ASAP7_75t_L g9979 ( 
.A1(n_7834),
.A2(n_7559),
.B(n_7534),
.Y(n_9979)
);

INVx4_ASAP7_75t_L g9980 ( 
.A(n_8919),
.Y(n_9980)
);

INVx1_ASAP7_75t_L g9981 ( 
.A(n_8432),
.Y(n_9981)
);

INVx2_ASAP7_75t_L g9982 ( 
.A(n_8017),
.Y(n_9982)
);

BUFx6f_ASAP7_75t_L g9983 ( 
.A(n_8114),
.Y(n_9983)
);

OR2x6_ASAP7_75t_L g9984 ( 
.A(n_8404),
.B(n_6807),
.Y(n_9984)
);

AO21x2_ASAP7_75t_L g9985 ( 
.A1(n_7834),
.A2(n_7835),
.B(n_8685),
.Y(n_9985)
);

BUFx3_ASAP7_75t_L g9986 ( 
.A(n_8126),
.Y(n_9986)
);

OAI22xp5_ASAP7_75t_L g9987 ( 
.A1(n_7956),
.A2(n_7392),
.B1(n_7370),
.B2(n_7369),
.Y(n_9987)
);

INVx2_ASAP7_75t_L g9988 ( 
.A(n_8017),
.Y(n_9988)
);

AOI22xp33_ASAP7_75t_L g9989 ( 
.A1(n_8355),
.A2(n_5719),
.B1(n_5742),
.B2(n_5739),
.Y(n_9989)
);

BUFx6f_ASAP7_75t_L g9990 ( 
.A(n_8114),
.Y(n_9990)
);

INVx2_ASAP7_75t_L g9991 ( 
.A(n_8039),
.Y(n_9991)
);

HB1xp67_ASAP7_75t_L g9992 ( 
.A(n_8721),
.Y(n_9992)
);

HB1xp67_ASAP7_75t_L g9993 ( 
.A(n_8721),
.Y(n_9993)
);

OA21x2_ASAP7_75t_L g9994 ( 
.A1(n_7718),
.A2(n_8746),
.B(n_7813),
.Y(n_9994)
);

HB1xp67_ASAP7_75t_L g9995 ( 
.A(n_8116),
.Y(n_9995)
);

BUFx12f_ASAP7_75t_L g9996 ( 
.A(n_8069),
.Y(n_9996)
);

OAI22xp5_ASAP7_75t_L g9997 ( 
.A1(n_8086),
.A2(n_7369),
.B1(n_7243),
.B2(n_7614),
.Y(n_9997)
);

INVx1_ASAP7_75t_L g9998 ( 
.A(n_8445),
.Y(n_9998)
);

AOI22xp5_ASAP7_75t_L g9999 ( 
.A1(n_8172),
.A2(n_7592),
.B1(n_7663),
.B2(n_7661),
.Y(n_9999)
);

NAND2xp5_ASAP7_75t_L g10000 ( 
.A(n_8409),
.B(n_7305),
.Y(n_10000)
);

HB1xp67_ASAP7_75t_L g10001 ( 
.A(n_8116),
.Y(n_10001)
);

INVx2_ASAP7_75t_L g10002 ( 
.A(n_8039),
.Y(n_10002)
);

BUFx8_ASAP7_75t_L g10003 ( 
.A(n_8239),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_8445),
.Y(n_10004)
);

BUFx4f_ASAP7_75t_SL g10005 ( 
.A(n_8069),
.Y(n_10005)
);

BUFx3_ASAP7_75t_L g10006 ( 
.A(n_8126),
.Y(n_10006)
);

AOI21x1_ASAP7_75t_L g10007 ( 
.A1(n_8682),
.A2(n_6947),
.B(n_6945),
.Y(n_10007)
);

OAI22xp33_ASAP7_75t_L g10008 ( 
.A1(n_8839),
.A2(n_7658),
.B1(n_7691),
.B2(n_7614),
.Y(n_10008)
);

CKINVDCx9p33_ASAP7_75t_R g10009 ( 
.A(n_8765),
.Y(n_10009)
);

INVx1_ASAP7_75t_L g10010 ( 
.A(n_8449),
.Y(n_10010)
);

BUFx6f_ASAP7_75t_L g10011 ( 
.A(n_8114),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_8449),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_8450),
.Y(n_10013)
);

OAI21x1_ASAP7_75t_L g10014 ( 
.A1(n_8248),
.A2(n_7036),
.B(n_7027),
.Y(n_10014)
);

INVx1_ASAP7_75t_L g10015 ( 
.A(n_8450),
.Y(n_10015)
);

INVx1_ASAP7_75t_L g10016 ( 
.A(n_8460),
.Y(n_10016)
);

INVx2_ASAP7_75t_L g10017 ( 
.A(n_8039),
.Y(n_10017)
);

INVx1_ASAP7_75t_L g10018 ( 
.A(n_8460),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_8465),
.Y(n_10019)
);

INVx1_ASAP7_75t_L g10020 ( 
.A(n_8465),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_8470),
.Y(n_10021)
);

INVx2_ASAP7_75t_L g10022 ( 
.A(n_8051),
.Y(n_10022)
);

INVx1_ASAP7_75t_L g10023 ( 
.A(n_8470),
.Y(n_10023)
);

AOI22xp5_ASAP7_75t_L g10024 ( 
.A1(n_7865),
.A2(n_7592),
.B1(n_7663),
.B2(n_7661),
.Y(n_10024)
);

INVx2_ASAP7_75t_L g10025 ( 
.A(n_8051),
.Y(n_10025)
);

HB1xp67_ASAP7_75t_L g10026 ( 
.A(n_8223),
.Y(n_10026)
);

INVx2_ASAP7_75t_L g10027 ( 
.A(n_8051),
.Y(n_10027)
);

OAI21x1_ASAP7_75t_L g10028 ( 
.A1(n_8323),
.A2(n_7036),
.B(n_7027),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_8487),
.Y(n_10029)
);

BUFx3_ASAP7_75t_L g10030 ( 
.A(n_8126),
.Y(n_10030)
);

BUFx3_ASAP7_75t_L g10031 ( 
.A(n_8126),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_8487),
.Y(n_10032)
);

OAI22xp5_ASAP7_75t_L g10033 ( 
.A1(n_8086),
.A2(n_7243),
.B1(n_7691),
.B2(n_7658),
.Y(n_10033)
);

INVxp67_ASAP7_75t_SL g10034 ( 
.A(n_8152),
.Y(n_10034)
);

INVx1_ASAP7_75t_L g10035 ( 
.A(n_8510),
.Y(n_10035)
);

OAI21x1_ASAP7_75t_L g10036 ( 
.A1(n_7753),
.A2(n_7446),
.B(n_7036),
.Y(n_10036)
);

BUFx6f_ASAP7_75t_L g10037 ( 
.A(n_8114),
.Y(n_10037)
);

OAI22xp5_ASAP7_75t_L g10038 ( 
.A1(n_8020),
.A2(n_7658),
.B1(n_7691),
.B2(n_7135),
.Y(n_10038)
);

AOI21x1_ASAP7_75t_L g10039 ( 
.A1(n_8193),
.A2(n_6947),
.B(n_6945),
.Y(n_10039)
);

AOI22xp33_ASAP7_75t_SL g10040 ( 
.A1(n_8070),
.A2(n_7603),
.B1(n_7590),
.B2(n_7583),
.Y(n_10040)
);

INVx2_ASAP7_75t_L g10041 ( 
.A(n_8064),
.Y(n_10041)
);

INVx1_ASAP7_75t_L g10042 ( 
.A(n_8510),
.Y(n_10042)
);

BUFx6f_ASAP7_75t_SL g10043 ( 
.A(n_8069),
.Y(n_10043)
);

AND2x4_ASAP7_75t_L g10044 ( 
.A(n_8940),
.B(n_7389),
.Y(n_10044)
);

OAI21x1_ASAP7_75t_SL g10045 ( 
.A1(n_8152),
.A2(n_6939),
.B(n_6912),
.Y(n_10045)
);

NAND2xp5_ASAP7_75t_L g10046 ( 
.A(n_8409),
.B(n_7305),
.Y(n_10046)
);

INVx1_ASAP7_75t_L g10047 ( 
.A(n_8514),
.Y(n_10047)
);

INVx5_ASAP7_75t_L g10048 ( 
.A(n_8191),
.Y(n_10048)
);

INVx2_ASAP7_75t_L g10049 ( 
.A(n_8064),
.Y(n_10049)
);

OAI22xp33_ASAP7_75t_L g10050 ( 
.A1(n_8839),
.A2(n_7590),
.B1(n_7612),
.B2(n_7583),
.Y(n_10050)
);

INVx3_ASAP7_75t_L g10051 ( 
.A(n_8191),
.Y(n_10051)
);

INVx2_ASAP7_75t_SL g10052 ( 
.A(n_8820),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_8514),
.Y(n_10053)
);

AOI22xp5_ASAP7_75t_L g10054 ( 
.A1(n_7865),
.A2(n_7592),
.B1(n_7700),
.B2(n_7553),
.Y(n_10054)
);

OA21x2_ASAP7_75t_L g10055 ( 
.A1(n_8746),
.A2(n_6667),
.B(n_6659),
.Y(n_10055)
);

OAI21x1_ASAP7_75t_L g10056 ( 
.A1(n_8248),
.A2(n_7036),
.B(n_7027),
.Y(n_10056)
);

INVx3_ASAP7_75t_L g10057 ( 
.A(n_8191),
.Y(n_10057)
);

AND2x2_ASAP7_75t_L g10058 ( 
.A(n_8169),
.B(n_6827),
.Y(n_10058)
);

INVx1_ASAP7_75t_L g10059 ( 
.A(n_8525),
.Y(n_10059)
);

INVx2_ASAP7_75t_L g10060 ( 
.A(n_8064),
.Y(n_10060)
);

AND2x2_ASAP7_75t_L g10061 ( 
.A(n_8169),
.B(n_6827),
.Y(n_10061)
);

INVx3_ASAP7_75t_L g10062 ( 
.A(n_8191),
.Y(n_10062)
);

INVx2_ASAP7_75t_SL g10063 ( 
.A(n_8820),
.Y(n_10063)
);

BUFx3_ASAP7_75t_L g10064 ( 
.A(n_8126),
.Y(n_10064)
);

CKINVDCx20_ASAP7_75t_R g10065 ( 
.A(n_8846),
.Y(n_10065)
);

AND2x2_ASAP7_75t_L g10066 ( 
.A(n_8169),
.B(n_6827),
.Y(n_10066)
);

OAI22xp5_ASAP7_75t_L g10067 ( 
.A1(n_8020),
.A2(n_7135),
.B1(n_7641),
.B2(n_7631),
.Y(n_10067)
);

INVx1_ASAP7_75t_L g10068 ( 
.A(n_8525),
.Y(n_10068)
);

BUFx2_ASAP7_75t_R g10069 ( 
.A(n_8863),
.Y(n_10069)
);

AOI22xp33_ASAP7_75t_L g10070 ( 
.A1(n_8355),
.A2(n_5719),
.B1(n_5742),
.B2(n_5739),
.Y(n_10070)
);

INVx1_ASAP7_75t_SL g10071 ( 
.A(n_8135),
.Y(n_10071)
);

INVx3_ASAP7_75t_L g10072 ( 
.A(n_8191),
.Y(n_10072)
);

INVx2_ASAP7_75t_L g10073 ( 
.A(n_8091),
.Y(n_10073)
);

INVx2_ASAP7_75t_L g10074 ( 
.A(n_8091),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_8091),
.Y(n_10075)
);

NAND2xp5_ASAP7_75t_L g10076 ( 
.A(n_9015),
.B(n_7324),
.Y(n_10076)
);

INVx2_ASAP7_75t_L g10077 ( 
.A(n_8132),
.Y(n_10077)
);

BUFx3_ASAP7_75t_L g10078 ( 
.A(n_8834),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_8529),
.Y(n_10079)
);

INVx1_ASAP7_75t_L g10080 ( 
.A(n_8529),
.Y(n_10080)
);

INVx2_ASAP7_75t_SL g10081 ( 
.A(n_8820),
.Y(n_10081)
);

AOI21x1_ASAP7_75t_L g10082 ( 
.A1(n_8193),
.A2(n_6947),
.B(n_6945),
.Y(n_10082)
);

INVx1_ASAP7_75t_L g10083 ( 
.A(n_8539),
.Y(n_10083)
);

INVx2_ASAP7_75t_L g10084 ( 
.A(n_8132),
.Y(n_10084)
);

NAND2xp5_ASAP7_75t_L g10085 ( 
.A(n_9015),
.B(n_7324),
.Y(n_10085)
);

OAI22xp5_ASAP7_75t_L g10086 ( 
.A1(n_8200),
.A2(n_7645),
.B1(n_7662),
.B2(n_7641),
.Y(n_10086)
);

INVx3_ASAP7_75t_L g10087 ( 
.A(n_8191),
.Y(n_10087)
);

HB1xp67_ASAP7_75t_SL g10088 ( 
.A(n_8822),
.Y(n_10088)
);

OAI21xp5_ASAP7_75t_L g10089 ( 
.A1(n_8219),
.A2(n_7415),
.B(n_6934),
.Y(n_10089)
);

INVx3_ASAP7_75t_L g10090 ( 
.A(n_8191),
.Y(n_10090)
);

OAI22xp5_ASAP7_75t_L g10091 ( 
.A1(n_8200),
.A2(n_7995),
.B1(n_8184),
.B2(n_8438),
.Y(n_10091)
);

OAI21x1_ASAP7_75t_L g10092 ( 
.A1(n_8248),
.A2(n_7036),
.B(n_7027),
.Y(n_10092)
);

OAI21xp5_ASAP7_75t_SL g10093 ( 
.A1(n_8929),
.A2(n_7643),
.B(n_7402),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_8539),
.Y(n_10094)
);

INVx2_ASAP7_75t_SL g10095 ( 
.A(n_8820),
.Y(n_10095)
);

HB1xp67_ASAP7_75t_L g10096 ( 
.A(n_8223),
.Y(n_10096)
);

INVx2_ASAP7_75t_SL g10097 ( 
.A(n_8820),
.Y(n_10097)
);

AO21x2_ASAP7_75t_L g10098 ( 
.A1(n_7834),
.A2(n_7559),
.B(n_7534),
.Y(n_10098)
);

INVx1_ASAP7_75t_SL g10099 ( 
.A(n_8418),
.Y(n_10099)
);

AND2x2_ASAP7_75t_L g10100 ( 
.A(n_8272),
.B(n_6827),
.Y(n_10100)
);

CKINVDCx8_ASAP7_75t_R g10101 ( 
.A(n_8891),
.Y(n_10101)
);

BUFx8_ASAP7_75t_L g10102 ( 
.A(n_8444),
.Y(n_10102)
);

AND2x2_ASAP7_75t_L g10103 ( 
.A(n_8272),
.B(n_6827),
.Y(n_10103)
);

OA21x2_ASAP7_75t_L g10104 ( 
.A1(n_7813),
.A2(n_6667),
.B(n_6659),
.Y(n_10104)
);

HB1xp67_ASAP7_75t_L g10105 ( 
.A(n_8280),
.Y(n_10105)
);

OAI22xp5_ASAP7_75t_L g10106 ( 
.A1(n_7995),
.A2(n_7662),
.B1(n_7679),
.B2(n_7645),
.Y(n_10106)
);

INVx2_ASAP7_75t_L g10107 ( 
.A(n_8132),
.Y(n_10107)
);

BUFx12f_ASAP7_75t_L g10108 ( 
.A(n_8069),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_8542),
.Y(n_10109)
);

INVx3_ASAP7_75t_L g10110 ( 
.A(n_8191),
.Y(n_10110)
);

INVx1_ASAP7_75t_L g10111 ( 
.A(n_8542),
.Y(n_10111)
);

INVx11_ASAP7_75t_L g10112 ( 
.A(n_8444),
.Y(n_10112)
);

INVx1_ASAP7_75t_L g10113 ( 
.A(n_8563),
.Y(n_10113)
);

INVxp67_ASAP7_75t_L g10114 ( 
.A(n_7937),
.Y(n_10114)
);

INVx2_ASAP7_75t_L g10115 ( 
.A(n_8141),
.Y(n_10115)
);

INVx1_ASAP7_75t_L g10116 ( 
.A(n_8563),
.Y(n_10116)
);

OR2x6_ASAP7_75t_L g10117 ( 
.A(n_8586),
.B(n_6807),
.Y(n_10117)
);

INVx2_ASAP7_75t_L g10118 ( 
.A(n_9014),
.Y(n_10118)
);

INVx2_ASAP7_75t_L g10119 ( 
.A(n_9014),
.Y(n_10119)
);

INVx2_ASAP7_75t_L g10120 ( 
.A(n_9014),
.Y(n_10120)
);

AOI22xp33_ASAP7_75t_L g10121 ( 
.A1(n_7890),
.A2(n_5739),
.B1(n_5746),
.B2(n_5742),
.Y(n_10121)
);

HB1xp67_ASAP7_75t_L g10122 ( 
.A(n_8280),
.Y(n_10122)
);

INVx2_ASAP7_75t_L g10123 ( 
.A(n_8141),
.Y(n_10123)
);

INVx1_ASAP7_75t_L g10124 ( 
.A(n_8564),
.Y(n_10124)
);

OAI21x1_ASAP7_75t_SL g10125 ( 
.A1(n_8152),
.A2(n_6939),
.B(n_6912),
.Y(n_10125)
);

BUFx3_ASAP7_75t_L g10126 ( 
.A(n_8069),
.Y(n_10126)
);

INVx2_ASAP7_75t_L g10127 ( 
.A(n_8141),
.Y(n_10127)
);

INVx1_ASAP7_75t_L g10128 ( 
.A(n_8564),
.Y(n_10128)
);

AND2x2_ASAP7_75t_L g10129 ( 
.A(n_8272),
.B(n_8312),
.Y(n_10129)
);

INVx2_ASAP7_75t_L g10130 ( 
.A(n_8145),
.Y(n_10130)
);

OAI22xp5_ASAP7_75t_L g10131 ( 
.A1(n_7995),
.A2(n_7693),
.B1(n_7679),
.B2(n_7700),
.Y(n_10131)
);

INVx2_ASAP7_75t_L g10132 ( 
.A(n_8145),
.Y(n_10132)
);

AOI22xp33_ASAP7_75t_L g10133 ( 
.A1(n_7890),
.A2(n_5739),
.B1(n_5746),
.B2(n_5742),
.Y(n_10133)
);

INVx1_ASAP7_75t_L g10134 ( 
.A(n_8567),
.Y(n_10134)
);

INVx1_ASAP7_75t_L g10135 ( 
.A(n_8567),
.Y(n_10135)
);

AOI22xp33_ASAP7_75t_SL g10136 ( 
.A1(n_8070),
.A2(n_7603),
.B1(n_7590),
.B2(n_7583),
.Y(n_10136)
);

BUFx3_ASAP7_75t_L g10137 ( 
.A(n_8148),
.Y(n_10137)
);

INVx1_ASAP7_75t_L g10138 ( 
.A(n_8570),
.Y(n_10138)
);

BUFx2_ASAP7_75t_R g10139 ( 
.A(n_8897),
.Y(n_10139)
);

BUFx2_ASAP7_75t_L g10140 ( 
.A(n_7939),
.Y(n_10140)
);

BUFx4_ASAP7_75t_SL g10141 ( 
.A(n_8822),
.Y(n_10141)
);

INVx2_ASAP7_75t_L g10142 ( 
.A(n_8145),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_8570),
.Y(n_10143)
);

INVx1_ASAP7_75t_L g10144 ( 
.A(n_8572),
.Y(n_10144)
);

INVx2_ASAP7_75t_L g10145 ( 
.A(n_8165),
.Y(n_10145)
);

CKINVDCx5p33_ASAP7_75t_R g10146 ( 
.A(n_8358),
.Y(n_10146)
);

INVx1_ASAP7_75t_L g10147 ( 
.A(n_8572),
.Y(n_10147)
);

BUFx8_ASAP7_75t_L g10148 ( 
.A(n_8612),
.Y(n_10148)
);

OAI21xp5_ASAP7_75t_L g10149 ( 
.A1(n_8219),
.A2(n_7415),
.B(n_7410),
.Y(n_10149)
);

OA21x2_ASAP7_75t_L g10150 ( 
.A1(n_7813),
.A2(n_6702),
.B(n_6681),
.Y(n_10150)
);

OAI21x1_ASAP7_75t_L g10151 ( 
.A1(n_8814),
.A2(n_7048),
.B(n_7036),
.Y(n_10151)
);

INVx1_ASAP7_75t_L g10152 ( 
.A(n_8579),
.Y(n_10152)
);

HB1xp67_ASAP7_75t_L g10153 ( 
.A(n_8298),
.Y(n_10153)
);

INVx3_ASAP7_75t_L g10154 ( 
.A(n_8278),
.Y(n_10154)
);

INVx1_ASAP7_75t_L g10155 ( 
.A(n_8579),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_8165),
.Y(n_10156)
);

BUFx8_ASAP7_75t_L g10157 ( 
.A(n_8684),
.Y(n_10157)
);

AOI22xp33_ASAP7_75t_L g10158 ( 
.A1(n_8467),
.A2(n_5746),
.B1(n_5761),
.B2(n_6014),
.Y(n_10158)
);

NAND2xp5_ASAP7_75t_L g10159 ( 
.A(n_8014),
.B(n_7332),
.Y(n_10159)
);

AOI22xp33_ASAP7_75t_L g10160 ( 
.A1(n_8467),
.A2(n_5746),
.B1(n_5761),
.B2(n_6014),
.Y(n_10160)
);

INVx1_ASAP7_75t_L g10161 ( 
.A(n_8584),
.Y(n_10161)
);

CKINVDCx11_ASAP7_75t_R g10162 ( 
.A(n_8148),
.Y(n_10162)
);

AOI21x1_ASAP7_75t_L g10163 ( 
.A1(n_8193),
.A2(n_6961),
.B(n_6947),
.Y(n_10163)
);

INVx1_ASAP7_75t_L g10164 ( 
.A(n_8584),
.Y(n_10164)
);

BUFx2_ASAP7_75t_R g10165 ( 
.A(n_8586),
.Y(n_10165)
);

INVx2_ASAP7_75t_SL g10166 ( 
.A(n_8988),
.Y(n_10166)
);

BUFx3_ASAP7_75t_L g10167 ( 
.A(n_8148),
.Y(n_10167)
);

AND2x4_ASAP7_75t_L g10168 ( 
.A(n_9024),
.B(n_7389),
.Y(n_10168)
);

AND2x4_ASAP7_75t_L g10169 ( 
.A(n_9024),
.B(n_7389),
.Y(n_10169)
);

INVx2_ASAP7_75t_SL g10170 ( 
.A(n_8988),
.Y(n_10170)
);

INVx2_ASAP7_75t_L g10171 ( 
.A(n_8165),
.Y(n_10171)
);

INVx1_ASAP7_75t_L g10172 ( 
.A(n_8596),
.Y(n_10172)
);

INVx2_ASAP7_75t_L g10173 ( 
.A(n_8180),
.Y(n_10173)
);

INVx6_ASAP7_75t_L g10174 ( 
.A(n_8148),
.Y(n_10174)
);

BUFx2_ASAP7_75t_L g10175 ( 
.A(n_7939),
.Y(n_10175)
);

AOI22xp33_ASAP7_75t_SL g10176 ( 
.A1(n_8315),
.A2(n_7603),
.B1(n_7644),
.B2(n_7612),
.Y(n_10176)
);

BUFx2_ASAP7_75t_R g10177 ( 
.A(n_8716),
.Y(n_10177)
);

CKINVDCx5p33_ASAP7_75t_R g10178 ( 
.A(n_8358),
.Y(n_10178)
);

INVx1_ASAP7_75t_L g10179 ( 
.A(n_8596),
.Y(n_10179)
);

AO21x1_ASAP7_75t_L g10180 ( 
.A1(n_7963),
.A2(n_7067),
.B(n_7062),
.Y(n_10180)
);

AOI21xp33_ASAP7_75t_L g10181 ( 
.A1(n_8027),
.A2(n_7415),
.B(n_7468),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_8599),
.Y(n_10182)
);

HB1xp67_ASAP7_75t_L g10183 ( 
.A(n_8298),
.Y(n_10183)
);

BUFx12f_ASAP7_75t_L g10184 ( 
.A(n_8148),
.Y(n_10184)
);

INVx1_ASAP7_75t_L g10185 ( 
.A(n_8599),
.Y(n_10185)
);

INVx2_ASAP7_75t_L g10186 ( 
.A(n_8180),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_8180),
.Y(n_10187)
);

OAI21x1_ASAP7_75t_L g10188 ( 
.A1(n_8323),
.A2(n_7055),
.B(n_7048),
.Y(n_10188)
);

AOI21x1_ASAP7_75t_L g10189 ( 
.A1(n_7829),
.A2(n_6963),
.B(n_6961),
.Y(n_10189)
);

OR2x6_ASAP7_75t_L g10190 ( 
.A(n_8716),
.B(n_6807),
.Y(n_10190)
);

INVx2_ASAP7_75t_L g10191 ( 
.A(n_8236),
.Y(n_10191)
);

INVx2_ASAP7_75t_SL g10192 ( 
.A(n_8988),
.Y(n_10192)
);

INVx1_ASAP7_75t_L g10193 ( 
.A(n_8600),
.Y(n_10193)
);

CKINVDCx11_ASAP7_75t_R g10194 ( 
.A(n_8215),
.Y(n_10194)
);

INVx1_ASAP7_75t_L g10195 ( 
.A(n_8600),
.Y(n_10195)
);

INVx4_ASAP7_75t_L g10196 ( 
.A(n_8215),
.Y(n_10196)
);

INVx2_ASAP7_75t_L g10197 ( 
.A(n_8236),
.Y(n_10197)
);

AND2x4_ASAP7_75t_L g10198 ( 
.A(n_9024),
.B(n_7426),
.Y(n_10198)
);

INVx1_ASAP7_75t_L g10199 ( 
.A(n_8608),
.Y(n_10199)
);

BUFx3_ASAP7_75t_L g10200 ( 
.A(n_8215),
.Y(n_10200)
);

INVx1_ASAP7_75t_SL g10201 ( 
.A(n_8418),
.Y(n_10201)
);

AND2x2_ASAP7_75t_L g10202 ( 
.A(n_8312),
.B(n_6829),
.Y(n_10202)
);

INVx1_ASAP7_75t_L g10203 ( 
.A(n_8608),
.Y(n_10203)
);

AOI22xp33_ASAP7_75t_L g10204 ( 
.A1(n_8277),
.A2(n_5746),
.B1(n_5761),
.B2(n_6014),
.Y(n_10204)
);

INVx2_ASAP7_75t_L g10205 ( 
.A(n_8236),
.Y(n_10205)
);

OAI22xp33_ASAP7_75t_L g10206 ( 
.A1(n_8544),
.A2(n_7644),
.B1(n_7647),
.B2(n_7612),
.Y(n_10206)
);

AOI22xp33_ASAP7_75t_L g10207 ( 
.A1(n_8277),
.A2(n_5761),
.B1(n_6021),
.B2(n_6014),
.Y(n_10207)
);

INVx1_ASAP7_75t_L g10208 ( 
.A(n_8611),
.Y(n_10208)
);

AOI22xp33_ASAP7_75t_SL g10209 ( 
.A1(n_8315),
.A2(n_7644),
.B1(n_7647),
.B2(n_7612),
.Y(n_10209)
);

INVx5_ASAP7_75t_L g10210 ( 
.A(n_8278),
.Y(n_10210)
);

INVx2_ASAP7_75t_SL g10211 ( 
.A(n_8988),
.Y(n_10211)
);

INVx2_ASAP7_75t_L g10212 ( 
.A(n_8253),
.Y(n_10212)
);

AND2x2_ASAP7_75t_L g10213 ( 
.A(n_8312),
.B(n_6829),
.Y(n_10213)
);

AOI22xp33_ASAP7_75t_L g10214 ( 
.A1(n_8857),
.A2(n_5761),
.B1(n_6021),
.B2(n_6014),
.Y(n_10214)
);

INVxp67_ASAP7_75t_SL g10215 ( 
.A(n_8401),
.Y(n_10215)
);

INVx3_ASAP7_75t_L g10216 ( 
.A(n_8278),
.Y(n_10216)
);

INVx1_ASAP7_75t_L g10217 ( 
.A(n_8611),
.Y(n_10217)
);

INVx2_ASAP7_75t_L g10218 ( 
.A(n_8253),
.Y(n_10218)
);

BUFx2_ASAP7_75t_R g10219 ( 
.A(n_9010),
.Y(n_10219)
);

INVx6_ASAP7_75t_L g10220 ( 
.A(n_8215),
.Y(n_10220)
);

NAND2xp5_ASAP7_75t_L g10221 ( 
.A(n_8014),
.B(n_7332),
.Y(n_10221)
);

INVx2_ASAP7_75t_SL g10222 ( 
.A(n_8988),
.Y(n_10222)
);

AO21x1_ASAP7_75t_SL g10223 ( 
.A1(n_8338),
.A2(n_7473),
.B(n_7468),
.Y(n_10223)
);

BUFx2_ASAP7_75t_L g10224 ( 
.A(n_7939),
.Y(n_10224)
);

AOI22xp33_ASAP7_75t_L g10225 ( 
.A1(n_8857),
.A2(n_6021),
.B1(n_6051),
.B2(n_6025),
.Y(n_10225)
);

INVx2_ASAP7_75t_L g10226 ( 
.A(n_8253),
.Y(n_10226)
);

AO21x2_ASAP7_75t_L g10227 ( 
.A1(n_7835),
.A2(n_7653),
.B(n_7623),
.Y(n_10227)
);

AO21x2_ASAP7_75t_L g10228 ( 
.A1(n_7835),
.A2(n_7653),
.B(n_7623),
.Y(n_10228)
);

OAI22xp33_ASAP7_75t_R g10229 ( 
.A1(n_7754),
.A2(n_7402),
.B1(n_7553),
.B2(n_7552),
.Y(n_10229)
);

INVx2_ASAP7_75t_L g10230 ( 
.A(n_8268),
.Y(n_10230)
);

INVx1_ASAP7_75t_L g10231 ( 
.A(n_8618),
.Y(n_10231)
);

AO22x1_ASAP7_75t_L g10232 ( 
.A1(n_7871),
.A2(n_7693),
.B1(n_7385),
.B2(n_7397),
.Y(n_10232)
);

NAND2x1p5_ASAP7_75t_L g10233 ( 
.A(n_8738),
.B(n_7133),
.Y(n_10233)
);

BUFx6f_ASAP7_75t_L g10234 ( 
.A(n_8278),
.Y(n_10234)
);

AOI22xp33_ASAP7_75t_L g10235 ( 
.A1(n_8634),
.A2(n_6021),
.B1(n_6051),
.B2(n_6025),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_8618),
.Y(n_10236)
);

AOI22xp33_ASAP7_75t_L g10237 ( 
.A1(n_8634),
.A2(n_6021),
.B1(n_6051),
.B2(n_6025),
.Y(n_10237)
);

INVx1_ASAP7_75t_SL g10238 ( 
.A(n_8435),
.Y(n_10238)
);

BUFx12f_ASAP7_75t_L g10239 ( 
.A(n_8215),
.Y(n_10239)
);

OAI21xp33_ASAP7_75t_SL g10240 ( 
.A1(n_8319),
.A2(n_7643),
.B(n_7075),
.Y(n_10240)
);

AOI22xp33_ASAP7_75t_L g10241 ( 
.A1(n_8616),
.A2(n_6021),
.B1(n_6051),
.B2(n_6025),
.Y(n_10241)
);

INVx2_ASAP7_75t_L g10242 ( 
.A(n_8268),
.Y(n_10242)
);

AND2x2_ASAP7_75t_L g10243 ( 
.A(n_8342),
.B(n_6829),
.Y(n_10243)
);

INVx2_ASAP7_75t_L g10244 ( 
.A(n_8268),
.Y(n_10244)
);

INVx4_ASAP7_75t_L g10245 ( 
.A(n_8481),
.Y(n_10245)
);

AOI22xp33_ASAP7_75t_L g10246 ( 
.A1(n_8616),
.A2(n_8090),
.B1(n_8026),
.B2(n_7973),
.Y(n_10246)
);

INVx2_ASAP7_75t_L g10247 ( 
.A(n_8295),
.Y(n_10247)
);

OAI21x1_ASAP7_75t_L g10248 ( 
.A1(n_7753),
.A2(n_7055),
.B(n_7048),
.Y(n_10248)
);

INVx2_ASAP7_75t_L g10249 ( 
.A(n_8295),
.Y(n_10249)
);

AOI22xp33_ASAP7_75t_L g10250 ( 
.A1(n_8090),
.A2(n_6021),
.B1(n_6051),
.B2(n_6025),
.Y(n_10250)
);

AND2x2_ASAP7_75t_L g10251 ( 
.A(n_8342),
.B(n_6829),
.Y(n_10251)
);

OAI22xp5_ASAP7_75t_L g10252 ( 
.A1(n_8184),
.A2(n_7647),
.B1(n_7644),
.B2(n_7385),
.Y(n_10252)
);

BUFx2_ASAP7_75t_L g10253 ( 
.A(n_8160),
.Y(n_10253)
);

HB1xp67_ASAP7_75t_L g10254 ( 
.A(n_8504),
.Y(n_10254)
);

INVx3_ASAP7_75t_L g10255 ( 
.A(n_8278),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_8619),
.Y(n_10256)
);

INVx1_ASAP7_75t_L g10257 ( 
.A(n_8619),
.Y(n_10257)
);

INVx2_ASAP7_75t_L g10258 ( 
.A(n_8295),
.Y(n_10258)
);

INVx1_ASAP7_75t_L g10259 ( 
.A(n_8620),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_8620),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_8621),
.Y(n_10261)
);

INVx2_ASAP7_75t_L g10262 ( 
.A(n_8305),
.Y(n_10262)
);

BUFx4f_ASAP7_75t_SL g10263 ( 
.A(n_8481),
.Y(n_10263)
);

INVx2_ASAP7_75t_L g10264 ( 
.A(n_8305),
.Y(n_10264)
);

OAI22xp5_ASAP7_75t_L g10265 ( 
.A1(n_8438),
.A2(n_7647),
.B1(n_7397),
.B2(n_7404),
.Y(n_10265)
);

INVx2_ASAP7_75t_L g10266 ( 
.A(n_8305),
.Y(n_10266)
);

INVx2_ASAP7_75t_L g10267 ( 
.A(n_8388),
.Y(n_10267)
);

INVx5_ASAP7_75t_L g10268 ( 
.A(n_8278),
.Y(n_10268)
);

AND2x2_ASAP7_75t_L g10269 ( 
.A(n_8342),
.B(n_6829),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_8621),
.Y(n_10270)
);

AND2x4_ASAP7_75t_L g10271 ( 
.A(n_9024),
.B(n_8959),
.Y(n_10271)
);

AOI22xp33_ASAP7_75t_SL g10272 ( 
.A1(n_8894),
.A2(n_6025),
.B1(n_6051),
.B2(n_6021),
.Y(n_10272)
);

AOI22xp33_ASAP7_75t_L g10273 ( 
.A1(n_8026),
.A2(n_6025),
.B1(n_6065),
.B2(n_6051),
.Y(n_10273)
);

INVx1_ASAP7_75t_L g10274 ( 
.A(n_8627),
.Y(n_10274)
);

INVx1_ASAP7_75t_L g10275 ( 
.A(n_8627),
.Y(n_10275)
);

INVx1_ASAP7_75t_L g10276 ( 
.A(n_8640),
.Y(n_10276)
);

BUFx6f_ASAP7_75t_L g10277 ( 
.A(n_8278),
.Y(n_10277)
);

AO21x1_ASAP7_75t_L g10278 ( 
.A1(n_8401),
.A2(n_8929),
.B(n_8214),
.Y(n_10278)
);

AO21x1_ASAP7_75t_SL g10279 ( 
.A1(n_8338),
.A2(n_7473),
.B(n_7468),
.Y(n_10279)
);

AOI21x1_ASAP7_75t_L g10280 ( 
.A1(n_7829),
.A2(n_6963),
.B(n_6961),
.Y(n_10280)
);

INVx1_ASAP7_75t_L g10281 ( 
.A(n_8640),
.Y(n_10281)
);

HB1xp67_ASAP7_75t_L g10282 ( 
.A(n_8504),
.Y(n_10282)
);

INVx2_ASAP7_75t_L g10283 ( 
.A(n_8388),
.Y(n_10283)
);

AOI22xp33_ASAP7_75t_L g10284 ( 
.A1(n_8026),
.A2(n_7973),
.B1(n_7782),
.B2(n_8993),
.Y(n_10284)
);

INVx1_ASAP7_75t_L g10285 ( 
.A(n_8644),
.Y(n_10285)
);

AND2x2_ASAP7_75t_L g10286 ( 
.A(n_8375),
.B(n_8377),
.Y(n_10286)
);

INVx2_ASAP7_75t_L g10287 ( 
.A(n_8388),
.Y(n_10287)
);

AOI22xp33_ASAP7_75t_SL g10288 ( 
.A1(n_8894),
.A2(n_6051),
.B1(n_6065),
.B2(n_6025),
.Y(n_10288)
);

OAI22xp5_ASAP7_75t_L g10289 ( 
.A1(n_8194),
.A2(n_7404),
.B1(n_7406),
.B2(n_7374),
.Y(n_10289)
);

AOI22xp33_ASAP7_75t_SL g10290 ( 
.A1(n_8894),
.A2(n_6071),
.B1(n_6065),
.B2(n_6965),
.Y(n_10290)
);

INVx2_ASAP7_75t_L g10291 ( 
.A(n_8412),
.Y(n_10291)
);

HB1xp67_ASAP7_75t_L g10292 ( 
.A(n_8751),
.Y(n_10292)
);

INVx1_ASAP7_75t_L g10293 ( 
.A(n_8644),
.Y(n_10293)
);

HB1xp67_ASAP7_75t_L g10294 ( 
.A(n_8751),
.Y(n_10294)
);

CKINVDCx5p33_ASAP7_75t_R g10295 ( 
.A(n_7807),
.Y(n_10295)
);

INVx1_ASAP7_75t_L g10296 ( 
.A(n_8649),
.Y(n_10296)
);

OAI21x1_ASAP7_75t_L g10297 ( 
.A1(n_8935),
.A2(n_7055),
.B(n_7048),
.Y(n_10297)
);

INVx2_ASAP7_75t_L g10298 ( 
.A(n_8412),
.Y(n_10298)
);

AO21x1_ASAP7_75t_SL g10299 ( 
.A1(n_9002),
.A2(n_7491),
.B(n_7473),
.Y(n_10299)
);

INVx1_ASAP7_75t_L g10300 ( 
.A(n_8649),
.Y(n_10300)
);

AOI22xp33_ASAP7_75t_SL g10301 ( 
.A1(n_8004),
.A2(n_6071),
.B1(n_6065),
.B2(n_6965),
.Y(n_10301)
);

INVx1_ASAP7_75t_L g10302 ( 
.A(n_8662),
.Y(n_10302)
);

INVx3_ASAP7_75t_L g10303 ( 
.A(n_8278),
.Y(n_10303)
);

AOI22xp33_ASAP7_75t_L g10304 ( 
.A1(n_7973),
.A2(n_6065),
.B1(n_6071),
.B2(n_7552),
.Y(n_10304)
);

INVx2_ASAP7_75t_L g10305 ( 
.A(n_8412),
.Y(n_10305)
);

HB1xp67_ASAP7_75t_L g10306 ( 
.A(n_8751),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_8662),
.Y(n_10307)
);

AND2x2_ASAP7_75t_L g10308 ( 
.A(n_8375),
.B(n_6829),
.Y(n_10308)
);

INVx1_ASAP7_75t_L g10309 ( 
.A(n_8680),
.Y(n_10309)
);

INVx1_ASAP7_75t_L g10310 ( 
.A(n_8680),
.Y(n_10310)
);

INVx2_ASAP7_75t_L g10311 ( 
.A(n_8443),
.Y(n_10311)
);

BUFx2_ASAP7_75t_L g10312 ( 
.A(n_8160),
.Y(n_10312)
);

INVx3_ASAP7_75t_L g10313 ( 
.A(n_8282),
.Y(n_10313)
);

AOI21x1_ASAP7_75t_L g10314 ( 
.A1(n_7829),
.A2(n_6963),
.B(n_6961),
.Y(n_10314)
);

AOI22xp33_ASAP7_75t_L g10315 ( 
.A1(n_7782),
.A2(n_6065),
.B1(n_6071),
.B2(n_6449),
.Y(n_10315)
);

CKINVDCx20_ASAP7_75t_R g10316 ( 
.A(n_7807),
.Y(n_10316)
);

CKINVDCx5p33_ASAP7_75t_R g10317 ( 
.A(n_8481),
.Y(n_10317)
);

INVx2_ASAP7_75t_L g10318 ( 
.A(n_8443),
.Y(n_10318)
);

INVx2_ASAP7_75t_L g10319 ( 
.A(n_8443),
.Y(n_10319)
);

INVx2_ASAP7_75t_L g10320 ( 
.A(n_8448),
.Y(n_10320)
);

OAI21x1_ASAP7_75t_L g10321 ( 
.A1(n_7753),
.A2(n_7055),
.B(n_7048),
.Y(n_10321)
);

INVx2_ASAP7_75t_L g10322 ( 
.A(n_8448),
.Y(n_10322)
);

INVx2_ASAP7_75t_L g10323 ( 
.A(n_8448),
.Y(n_10323)
);

INVx1_ASAP7_75t_L g10324 ( 
.A(n_8687),
.Y(n_10324)
);

INVxp33_ASAP7_75t_L g10325 ( 
.A(n_8684),
.Y(n_10325)
);

INVx1_ASAP7_75t_L g10326 ( 
.A(n_8687),
.Y(n_10326)
);

INVx2_ASAP7_75t_L g10327 ( 
.A(n_8455),
.Y(n_10327)
);

NAND2x1p5_ASAP7_75t_L g10328 ( 
.A(n_8738),
.B(n_7199),
.Y(n_10328)
);

CKINVDCx8_ASAP7_75t_R g10329 ( 
.A(n_9010),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_8693),
.Y(n_10330)
);

INVx1_ASAP7_75t_L g10331 ( 
.A(n_8693),
.Y(n_10331)
);

INVx2_ASAP7_75t_L g10332 ( 
.A(n_8455),
.Y(n_10332)
);

INVx3_ASAP7_75t_L g10333 ( 
.A(n_8282),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_8694),
.Y(n_10334)
);

INVx1_ASAP7_75t_L g10335 ( 
.A(n_8694),
.Y(n_10335)
);

INVx1_ASAP7_75t_L g10336 ( 
.A(n_8702),
.Y(n_10336)
);

OAI21x1_ASAP7_75t_L g10337 ( 
.A1(n_8569),
.A2(n_7055),
.B(n_7048),
.Y(n_10337)
);

INVx1_ASAP7_75t_L g10338 ( 
.A(n_8702),
.Y(n_10338)
);

INVxp33_ASAP7_75t_L g10339 ( 
.A(n_8771),
.Y(n_10339)
);

HB1xp67_ASAP7_75t_L g10340 ( 
.A(n_8751),
.Y(n_10340)
);

INVx1_ASAP7_75t_SL g10341 ( 
.A(n_8435),
.Y(n_10341)
);

INVx1_ASAP7_75t_L g10342 ( 
.A(n_8705),
.Y(n_10342)
);

INVx1_ASAP7_75t_L g10343 ( 
.A(n_8705),
.Y(n_10343)
);

OAI22xp33_ASAP7_75t_L g10344 ( 
.A1(n_8544),
.A2(n_8772),
.B1(n_8777),
.B2(n_8767),
.Y(n_10344)
);

NAND2xp5_ASAP7_75t_L g10345 ( 
.A(n_8143),
.B(n_8171),
.Y(n_10345)
);

INVx1_ASAP7_75t_L g10346 ( 
.A(n_8709),
.Y(n_10346)
);

OAI22xp33_ASAP7_75t_L g10347 ( 
.A1(n_8767),
.A2(n_7140),
.B1(n_6982),
.B2(n_6065),
.Y(n_10347)
);

OAI21x1_ASAP7_75t_L g10348 ( 
.A1(n_8248),
.A2(n_7057),
.B(n_7055),
.Y(n_10348)
);

INVx2_ASAP7_75t_L g10349 ( 
.A(n_8455),
.Y(n_10349)
);

NAND2xp5_ASAP7_75t_L g10350 ( 
.A(n_8143),
.B(n_7344),
.Y(n_10350)
);

INVx2_ASAP7_75t_L g10351 ( 
.A(n_8472),
.Y(n_10351)
);

OAI22xp5_ASAP7_75t_L g10352 ( 
.A1(n_8194),
.A2(n_7406),
.B1(n_7416),
.B2(n_7374),
.Y(n_10352)
);

NAND2x1p5_ASAP7_75t_L g10353 ( 
.A(n_8805),
.B(n_7199),
.Y(n_10353)
);

BUFx2_ASAP7_75t_SL g10354 ( 
.A(n_8538),
.Y(n_10354)
);

OAI21xp5_ASAP7_75t_L g10355 ( 
.A1(n_8224),
.A2(n_7417),
.B(n_7410),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_8709),
.Y(n_10356)
);

INVx2_ASAP7_75t_L g10357 ( 
.A(n_8472),
.Y(n_10357)
);

INVx2_ASAP7_75t_L g10358 ( 
.A(n_8472),
.Y(n_10358)
);

INVx1_ASAP7_75t_L g10359 ( 
.A(n_8712),
.Y(n_10359)
);

AOI22xp33_ASAP7_75t_SL g10360 ( 
.A1(n_8004),
.A2(n_6071),
.B1(n_6065),
.B2(n_6965),
.Y(n_10360)
);

BUFx2_ASAP7_75t_SL g10361 ( 
.A(n_8666),
.Y(n_10361)
);

INVx1_ASAP7_75t_L g10362 ( 
.A(n_8712),
.Y(n_10362)
);

INVx1_ASAP7_75t_SL g10363 ( 
.A(n_8439),
.Y(n_10363)
);

AOI22xp33_ASAP7_75t_SL g10364 ( 
.A1(n_8004),
.A2(n_6071),
.B1(n_7139),
.B2(n_6965),
.Y(n_10364)
);

HB1xp67_ASAP7_75t_L g10365 ( 
.A(n_8751),
.Y(n_10365)
);

INVx1_ASAP7_75t_L g10366 ( 
.A(n_8713),
.Y(n_10366)
);

INVx2_ASAP7_75t_L g10367 ( 
.A(n_8480),
.Y(n_10367)
);

AOI22xp33_ASAP7_75t_L g10368 ( 
.A1(n_8993),
.A2(n_8330),
.B1(n_8562),
.B2(n_8545),
.Y(n_10368)
);

BUFx12f_ASAP7_75t_L g10369 ( 
.A(n_8481),
.Y(n_10369)
);

AND2x4_ASAP7_75t_L g10370 ( 
.A(n_8959),
.B(n_7426),
.Y(n_10370)
);

INVx2_ASAP7_75t_L g10371 ( 
.A(n_8480),
.Y(n_10371)
);

CKINVDCx6p67_ASAP7_75t_R g10372 ( 
.A(n_8481),
.Y(n_10372)
);

BUFx10_ASAP7_75t_L g10373 ( 
.A(n_8988),
.Y(n_10373)
);

INVx1_ASAP7_75t_L g10374 ( 
.A(n_8713),
.Y(n_10374)
);

AOI22xp33_ASAP7_75t_SL g10375 ( 
.A1(n_8332),
.A2(n_6071),
.B1(n_7139),
.B2(n_6965),
.Y(n_10375)
);

OAI22xp5_ASAP7_75t_L g10376 ( 
.A1(n_7840),
.A2(n_7416),
.B1(n_6894),
.B2(n_7067),
.Y(n_10376)
);

HB1xp67_ASAP7_75t_L g10377 ( 
.A(n_8812),
.Y(n_10377)
);

BUFx6f_ASAP7_75t_L g10378 ( 
.A(n_8282),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_8719),
.Y(n_10379)
);

INVx1_ASAP7_75t_L g10380 ( 
.A(n_8719),
.Y(n_10380)
);

INVx1_ASAP7_75t_L g10381 ( 
.A(n_8735),
.Y(n_10381)
);

INVx1_ASAP7_75t_L g10382 ( 
.A(n_9033),
.Y(n_10382)
);

OAI21x1_ASAP7_75t_L g10383 ( 
.A1(n_9053),
.A2(n_8238),
.B(n_8327),
.Y(n_10383)
);

INVx1_ASAP7_75t_L g10384 ( 
.A(n_9033),
.Y(n_10384)
);

INVx2_ASAP7_75t_L g10385 ( 
.A(n_9582),
.Y(n_10385)
);

AND2x2_ASAP7_75t_L g10386 ( 
.A(n_9727),
.B(n_7774),
.Y(n_10386)
);

NOR2xp33_ASAP7_75t_L g10387 ( 
.A(n_9144),
.B(n_9249),
.Y(n_10387)
);

INVx1_ASAP7_75t_L g10388 ( 
.A(n_9041),
.Y(n_10388)
);

NAND2xp5_ASAP7_75t_L g10389 ( 
.A(n_9119),
.B(n_7814),
.Y(n_10389)
);

BUFx3_ASAP7_75t_L g10390 ( 
.A(n_9338),
.Y(n_10390)
);

HB1xp67_ASAP7_75t_L g10391 ( 
.A(n_9995),
.Y(n_10391)
);

OR2x2_ASAP7_75t_L g10392 ( 
.A(n_9615),
.B(n_8076),
.Y(n_10392)
);

OAI21x1_ASAP7_75t_L g10393 ( 
.A1(n_9053),
.A2(n_8238),
.B(n_8327),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_9041),
.Y(n_10394)
);

AND2x2_ASAP7_75t_L g10395 ( 
.A(n_9727),
.B(n_7774),
.Y(n_10395)
);

INVx2_ASAP7_75t_L g10396 ( 
.A(n_9582),
.Y(n_10396)
);

HB1xp67_ASAP7_75t_L g10397 ( 
.A(n_10001),
.Y(n_10397)
);

INVx5_ASAP7_75t_L g10398 ( 
.A(n_9098),
.Y(n_10398)
);

INVx1_ASAP7_75t_L g10399 ( 
.A(n_9052),
.Y(n_10399)
);

INVx1_ASAP7_75t_L g10400 ( 
.A(n_9052),
.Y(n_10400)
);

INVx2_ASAP7_75t_L g10401 ( 
.A(n_9593),
.Y(n_10401)
);

INVx3_ASAP7_75t_L g10402 ( 
.A(n_10329),
.Y(n_10402)
);

AND2x2_ASAP7_75t_L g10403 ( 
.A(n_10215),
.B(n_8110),
.Y(n_10403)
);

CKINVDCx5p33_ASAP7_75t_R g10404 ( 
.A(n_10141),
.Y(n_10404)
);

OAI21x1_ASAP7_75t_L g10405 ( 
.A1(n_9053),
.A2(n_8238),
.B(n_8327),
.Y(n_10405)
);

INVx2_ASAP7_75t_L g10406 ( 
.A(n_9593),
.Y(n_10406)
);

INVx2_ASAP7_75t_L g10407 ( 
.A(n_9658),
.Y(n_10407)
);

INVx2_ASAP7_75t_SL g10408 ( 
.A(n_9931),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_9058),
.Y(n_10409)
);

INVx3_ASAP7_75t_L g10410 ( 
.A(n_10329),
.Y(n_10410)
);

AND2x2_ASAP7_75t_L g10411 ( 
.A(n_9888),
.B(n_8110),
.Y(n_10411)
);

INVx2_ASAP7_75t_L g10412 ( 
.A(n_9658),
.Y(n_10412)
);

INVx1_ASAP7_75t_L g10413 ( 
.A(n_9058),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_9059),
.Y(n_10414)
);

NAND2xp5_ASAP7_75t_L g10415 ( 
.A(n_9391),
.B(n_9155),
.Y(n_10415)
);

INVx2_ASAP7_75t_SL g10416 ( 
.A(n_9931),
.Y(n_10416)
);

INVx2_ASAP7_75t_SL g10417 ( 
.A(n_9931),
.Y(n_10417)
);

AOI221xp5_ASAP7_75t_L g10418 ( 
.A1(n_9530),
.A2(n_8234),
.B1(n_9002),
.B2(n_8631),
.C(n_8986),
.Y(n_10418)
);

INVx1_ASAP7_75t_L g10419 ( 
.A(n_9059),
.Y(n_10419)
);

INVx3_ASAP7_75t_L g10420 ( 
.A(n_9295),
.Y(n_10420)
);

BUFx2_ASAP7_75t_L g10421 ( 
.A(n_9254),
.Y(n_10421)
);

CKINVDCx11_ASAP7_75t_R g10422 ( 
.A(n_9057),
.Y(n_10422)
);

OAI22xp5_ASAP7_75t_L g10423 ( 
.A1(n_9512),
.A2(n_8562),
.B1(n_8628),
.B2(n_8545),
.Y(n_10423)
);

INVx3_ASAP7_75t_L g10424 ( 
.A(n_9295),
.Y(n_10424)
);

BUFx12f_ASAP7_75t_L g10425 ( 
.A(n_9338),
.Y(n_10425)
);

INVx2_ASAP7_75t_L g10426 ( 
.A(n_10007),
.Y(n_10426)
);

INVx1_ASAP7_75t_L g10427 ( 
.A(n_9060),
.Y(n_10427)
);

INVx1_ASAP7_75t_L g10428 ( 
.A(n_9060),
.Y(n_10428)
);

OR2x2_ASAP7_75t_L g10429 ( 
.A(n_9315),
.B(n_8171),
.Y(n_10429)
);

INVx1_ASAP7_75t_L g10430 ( 
.A(n_9061),
.Y(n_10430)
);

INVx1_ASAP7_75t_L g10431 ( 
.A(n_9061),
.Y(n_10431)
);

HB1xp67_ASAP7_75t_L g10432 ( 
.A(n_10026),
.Y(n_10432)
);

AOI21xp5_ASAP7_75t_L g10433 ( 
.A1(n_9418),
.A2(n_10091),
.B(n_9309),
.Y(n_10433)
);

AND2x2_ASAP7_75t_L g10434 ( 
.A(n_9888),
.B(n_8167),
.Y(n_10434)
);

INVx2_ASAP7_75t_SL g10435 ( 
.A(n_9931),
.Y(n_10435)
);

AOI22xp5_ASAP7_75t_SL g10436 ( 
.A1(n_10091),
.A2(n_8012),
.B1(n_8761),
.B2(n_8531),
.Y(n_10436)
);

INVx2_ASAP7_75t_L g10437 ( 
.A(n_10007),
.Y(n_10437)
);

AND2x2_ASAP7_75t_L g10438 ( 
.A(n_9034),
.B(n_8167),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_9064),
.Y(n_10439)
);

INVx1_ASAP7_75t_L g10440 ( 
.A(n_9064),
.Y(n_10440)
);

AND2x2_ASAP7_75t_L g10441 ( 
.A(n_9034),
.B(n_8285),
.Y(n_10441)
);

AND2x2_ASAP7_75t_L g10442 ( 
.A(n_9043),
.B(n_8285),
.Y(n_10442)
);

INVx1_ASAP7_75t_L g10443 ( 
.A(n_9065),
.Y(n_10443)
);

INVx1_ASAP7_75t_L g10444 ( 
.A(n_9065),
.Y(n_10444)
);

INVx2_ASAP7_75t_L g10445 ( 
.A(n_9040),
.Y(n_10445)
);

INVx2_ASAP7_75t_SL g10446 ( 
.A(n_9931),
.Y(n_10446)
);

INVx1_ASAP7_75t_L g10447 ( 
.A(n_9069),
.Y(n_10447)
);

INVx1_ASAP7_75t_L g10448 ( 
.A(n_9069),
.Y(n_10448)
);

INVx2_ASAP7_75t_SL g10449 ( 
.A(n_9295),
.Y(n_10449)
);

OAI21x1_ASAP7_75t_L g10450 ( 
.A1(n_9094),
.A2(n_8304),
.B(n_8469),
.Y(n_10450)
);

AOI21x1_ASAP7_75t_L g10451 ( 
.A1(n_10232),
.A2(n_8945),
.B(n_8801),
.Y(n_10451)
);

OA21x2_ASAP7_75t_L g10452 ( 
.A1(n_10034),
.A2(n_8792),
.B(n_8750),
.Y(n_10452)
);

INVx2_ASAP7_75t_L g10453 ( 
.A(n_9040),
.Y(n_10453)
);

CKINVDCx6p67_ASAP7_75t_R g10454 ( 
.A(n_9057),
.Y(n_10454)
);

HB1xp67_ASAP7_75t_L g10455 ( 
.A(n_10096),
.Y(n_10455)
);

HB1xp67_ASAP7_75t_L g10456 ( 
.A(n_10105),
.Y(n_10456)
);

INVx2_ASAP7_75t_L g10457 ( 
.A(n_9040),
.Y(n_10457)
);

INVx2_ASAP7_75t_L g10458 ( 
.A(n_9050),
.Y(n_10458)
);

BUFx2_ASAP7_75t_SL g10459 ( 
.A(n_10065),
.Y(n_10459)
);

INVx2_ASAP7_75t_L g10460 ( 
.A(n_9050),
.Y(n_10460)
);

BUFx3_ASAP7_75t_L g10461 ( 
.A(n_9338),
.Y(n_10461)
);

INVx2_ASAP7_75t_L g10462 ( 
.A(n_9050),
.Y(n_10462)
);

INVx1_ASAP7_75t_L g10463 ( 
.A(n_9071),
.Y(n_10463)
);

AOI21x1_ASAP7_75t_L g10464 ( 
.A1(n_10232),
.A2(n_8945),
.B(n_8801),
.Y(n_10464)
);

INVx2_ASAP7_75t_L g10465 ( 
.A(n_9054),
.Y(n_10465)
);

INVx1_ASAP7_75t_L g10466 ( 
.A(n_9071),
.Y(n_10466)
);

A2O1A1Ixp33_ASAP7_75t_L g10467 ( 
.A1(n_9418),
.A2(n_8234),
.B(n_8639),
.C(n_8214),
.Y(n_10467)
);

AND2x2_ASAP7_75t_L g10468 ( 
.A(n_9043),
.B(n_8490),
.Y(n_10468)
);

INVx2_ASAP7_75t_L g10469 ( 
.A(n_9054),
.Y(n_10469)
);

AND2x2_ASAP7_75t_L g10470 ( 
.A(n_9049),
.B(n_9717),
.Y(n_10470)
);

INVx2_ASAP7_75t_L g10471 ( 
.A(n_9054),
.Y(n_10471)
);

INVx2_ASAP7_75t_L g10472 ( 
.A(n_9063),
.Y(n_10472)
);

INVx4_ASAP7_75t_L g10473 ( 
.A(n_9098),
.Y(n_10473)
);

BUFx3_ASAP7_75t_L g10474 ( 
.A(n_9338),
.Y(n_10474)
);

INVx1_ASAP7_75t_L g10475 ( 
.A(n_9072),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_9072),
.Y(n_10476)
);

OAI21x1_ASAP7_75t_L g10477 ( 
.A1(n_9094),
.A2(n_8304),
.B(n_8469),
.Y(n_10477)
);

AO21x2_ASAP7_75t_L g10478 ( 
.A1(n_9550),
.A2(n_9572),
.B(n_9608),
.Y(n_10478)
);

INVx1_ASAP7_75t_L g10479 ( 
.A(n_9074),
.Y(n_10479)
);

AOI21xp5_ASAP7_75t_L g10480 ( 
.A1(n_9309),
.A2(n_8027),
.B(n_7776),
.Y(n_10480)
);

BUFx2_ASAP7_75t_L g10481 ( 
.A(n_9254),
.Y(n_10481)
);

BUFx2_ASAP7_75t_L g10482 ( 
.A(n_9254),
.Y(n_10482)
);

INVx1_ASAP7_75t_L g10483 ( 
.A(n_9074),
.Y(n_10483)
);

OAI21x1_ASAP7_75t_L g10484 ( 
.A1(n_9207),
.A2(n_8304),
.B(n_8469),
.Y(n_10484)
);

INVx2_ASAP7_75t_L g10485 ( 
.A(n_9063),
.Y(n_10485)
);

INVx3_ASAP7_75t_L g10486 ( 
.A(n_9295),
.Y(n_10486)
);

INVx2_ASAP7_75t_L g10487 ( 
.A(n_9063),
.Y(n_10487)
);

INVx2_ASAP7_75t_L g10488 ( 
.A(n_9078),
.Y(n_10488)
);

INVx1_ASAP7_75t_L g10489 ( 
.A(n_9075),
.Y(n_10489)
);

BUFx2_ASAP7_75t_L g10490 ( 
.A(n_9434),
.Y(n_10490)
);

INVx2_ASAP7_75t_L g10491 ( 
.A(n_9078),
.Y(n_10491)
);

INVx2_ASAP7_75t_SL g10492 ( 
.A(n_9295),
.Y(n_10492)
);

INVx2_ASAP7_75t_L g10493 ( 
.A(n_9078),
.Y(n_10493)
);

AO31x2_ASAP7_75t_L g10494 ( 
.A1(n_9949),
.A2(n_8416),
.A3(n_8300),
.B(n_7955),
.Y(n_10494)
);

INVx3_ASAP7_75t_L g10495 ( 
.A(n_9295),
.Y(n_10495)
);

AND2x2_ASAP7_75t_L g10496 ( 
.A(n_9049),
.B(n_8490),
.Y(n_10496)
);

BUFx3_ASAP7_75t_L g10497 ( 
.A(n_9471),
.Y(n_10497)
);

INVx2_ASAP7_75t_L g10498 ( 
.A(n_9079),
.Y(n_10498)
);

AND2x2_ASAP7_75t_L g10499 ( 
.A(n_9717),
.B(n_8490),
.Y(n_10499)
);

INVx1_ASAP7_75t_L g10500 ( 
.A(n_9075),
.Y(n_10500)
);

INVx1_ASAP7_75t_L g10501 ( 
.A(n_9076),
.Y(n_10501)
);

INVx1_ASAP7_75t_L g10502 ( 
.A(n_9076),
.Y(n_10502)
);

INVx1_ASAP7_75t_L g10503 ( 
.A(n_9082),
.Y(n_10503)
);

INVx2_ASAP7_75t_L g10504 ( 
.A(n_9079),
.Y(n_10504)
);

INVx2_ASAP7_75t_L g10505 ( 
.A(n_9079),
.Y(n_10505)
);

INVx1_ASAP7_75t_L g10506 ( 
.A(n_9082),
.Y(n_10506)
);

INVx2_ASAP7_75t_L g10507 ( 
.A(n_9520),
.Y(n_10507)
);

OA21x2_ASAP7_75t_L g10508 ( 
.A1(n_9741),
.A2(n_8792),
.B(n_8750),
.Y(n_10508)
);

AOI21x1_ASAP7_75t_L g10509 ( 
.A1(n_9374),
.A2(n_8666),
.B(n_8190),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9085),
.Y(n_10510)
);

INVx2_ASAP7_75t_SL g10511 ( 
.A(n_9591),
.Y(n_10511)
);

AND2x2_ASAP7_75t_L g10512 ( 
.A(n_9729),
.B(n_8490),
.Y(n_10512)
);

INVx2_ASAP7_75t_L g10513 ( 
.A(n_9520),
.Y(n_10513)
);

INVx1_ASAP7_75t_L g10514 ( 
.A(n_9085),
.Y(n_10514)
);

AND2x2_ASAP7_75t_L g10515 ( 
.A(n_9729),
.B(n_8490),
.Y(n_10515)
);

OAI21x1_ASAP7_75t_L g10516 ( 
.A1(n_9207),
.A2(n_8077),
.B(n_8826),
.Y(n_10516)
);

OA21x2_ASAP7_75t_L g10517 ( 
.A1(n_9856),
.A2(n_8792),
.B(n_8750),
.Y(n_10517)
);

AND2x2_ASAP7_75t_L g10518 ( 
.A(n_9845),
.B(n_8520),
.Y(n_10518)
);

INVx1_ASAP7_75t_L g10519 ( 
.A(n_9087),
.Y(n_10519)
);

NOR2xp33_ASAP7_75t_L g10520 ( 
.A(n_9144),
.B(n_8012),
.Y(n_10520)
);

HB1xp67_ASAP7_75t_L g10521 ( 
.A(n_10122),
.Y(n_10521)
);

INVx2_ASAP7_75t_L g10522 ( 
.A(n_9520),
.Y(n_10522)
);

AOI22xp33_ASAP7_75t_L g10523 ( 
.A1(n_9405),
.A2(n_7810),
.B1(n_8330),
.B2(n_8224),
.Y(n_10523)
);

NAND2xp5_ASAP7_75t_L g10524 ( 
.A(n_9155),
.B(n_8084),
.Y(n_10524)
);

INVx1_ASAP7_75t_L g10525 ( 
.A(n_9087),
.Y(n_10525)
);

INVx2_ASAP7_75t_L g10526 ( 
.A(n_9525),
.Y(n_10526)
);

INVx1_ASAP7_75t_L g10527 ( 
.A(n_9093),
.Y(n_10527)
);

AOI22xp5_ASAP7_75t_L g10528 ( 
.A1(n_10229),
.A2(n_9557),
.B1(n_9536),
.B2(n_9556),
.Y(n_10528)
);

INVx2_ASAP7_75t_SL g10529 ( 
.A(n_9295),
.Y(n_10529)
);

INVx1_ASAP7_75t_SL g10530 ( 
.A(n_9135),
.Y(n_10530)
);

INVx2_ASAP7_75t_L g10531 ( 
.A(n_9525),
.Y(n_10531)
);

BUFx2_ASAP7_75t_L g10532 ( 
.A(n_9434),
.Y(n_10532)
);

INVx1_ASAP7_75t_L g10533 ( 
.A(n_9093),
.Y(n_10533)
);

INVx3_ASAP7_75t_L g10534 ( 
.A(n_9514),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_9101),
.Y(n_10535)
);

INVx3_ASAP7_75t_L g10536 ( 
.A(n_9514),
.Y(n_10536)
);

INVx1_ASAP7_75t_L g10537 ( 
.A(n_9101),
.Y(n_10537)
);

OAI21xp5_ASAP7_75t_L g10538 ( 
.A1(n_9250),
.A2(n_8654),
.B(n_8986),
.Y(n_10538)
);

INVx2_ASAP7_75t_L g10539 ( 
.A(n_9525),
.Y(n_10539)
);

INVx2_ASAP7_75t_L g10540 ( 
.A(n_9529),
.Y(n_10540)
);

INVx2_ASAP7_75t_L g10541 ( 
.A(n_9529),
.Y(n_10541)
);

AND2x2_ASAP7_75t_L g10542 ( 
.A(n_9845),
.B(n_8520),
.Y(n_10542)
);

OAI21x1_ASAP7_75t_L g10543 ( 
.A1(n_9207),
.A2(n_8077),
.B(n_8826),
.Y(n_10543)
);

AND2x2_ASAP7_75t_L g10544 ( 
.A(n_9846),
.B(n_8520),
.Y(n_10544)
);

INVx2_ASAP7_75t_L g10545 ( 
.A(n_9529),
.Y(n_10545)
);

HB1xp67_ASAP7_75t_L g10546 ( 
.A(n_10153),
.Y(n_10546)
);

AND2x4_ASAP7_75t_L g10547 ( 
.A(n_9950),
.B(n_7719),
.Y(n_10547)
);

CKINVDCx5p33_ASAP7_75t_R g10548 ( 
.A(n_9471),
.Y(n_10548)
);

NAND2xp5_ASAP7_75t_L g10549 ( 
.A(n_9158),
.B(n_9170),
.Y(n_10549)
);

INVx2_ASAP7_75t_L g10550 ( 
.A(n_9540),
.Y(n_10550)
);

INVx1_ASAP7_75t_L g10551 ( 
.A(n_9107),
.Y(n_10551)
);

OR2x2_ASAP7_75t_L g10552 ( 
.A(n_9315),
.B(n_8185),
.Y(n_10552)
);

INVx1_ASAP7_75t_L g10553 ( 
.A(n_9107),
.Y(n_10553)
);

AND2x2_ASAP7_75t_L g10554 ( 
.A(n_9846),
.B(n_8520),
.Y(n_10554)
);

NOR2xp33_ASAP7_75t_L g10555 ( 
.A(n_9249),
.B(n_8084),
.Y(n_10555)
);

INVx2_ASAP7_75t_L g10556 ( 
.A(n_9540),
.Y(n_10556)
);

AND2x2_ASAP7_75t_L g10557 ( 
.A(n_9850),
.B(n_8520),
.Y(n_10557)
);

NAND2x1p5_ASAP7_75t_L g10558 ( 
.A(n_9514),
.B(n_8805),
.Y(n_10558)
);

INVx2_ASAP7_75t_L g10559 ( 
.A(n_9540),
.Y(n_10559)
);

BUFx3_ASAP7_75t_L g10560 ( 
.A(n_9471),
.Y(n_10560)
);

INVx1_ASAP7_75t_L g10561 ( 
.A(n_9109),
.Y(n_10561)
);

INVx1_ASAP7_75t_SL g10562 ( 
.A(n_9135),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_9545),
.Y(n_10563)
);

INVx2_ASAP7_75t_L g10564 ( 
.A(n_9545),
.Y(n_10564)
);

AND2x4_ASAP7_75t_SL g10565 ( 
.A(n_9454),
.B(n_8531),
.Y(n_10565)
);

BUFx2_ASAP7_75t_L g10566 ( 
.A(n_9434),
.Y(n_10566)
);

INVxp67_ASAP7_75t_L g10567 ( 
.A(n_9386),
.Y(n_10567)
);

INVx1_ASAP7_75t_L g10568 ( 
.A(n_9109),
.Y(n_10568)
);

INVx2_ASAP7_75t_L g10569 ( 
.A(n_9545),
.Y(n_10569)
);

NAND2x1p5_ASAP7_75t_L g10570 ( 
.A(n_9514),
.B(n_8805),
.Y(n_10570)
);

INVx1_ASAP7_75t_L g10571 ( 
.A(n_9111),
.Y(n_10571)
);

INVx1_ASAP7_75t_L g10572 ( 
.A(n_9111),
.Y(n_10572)
);

INVx1_ASAP7_75t_L g10573 ( 
.A(n_9113),
.Y(n_10573)
);

INVx2_ASAP7_75t_L g10574 ( 
.A(n_9576),
.Y(n_10574)
);

OAI22xp5_ASAP7_75t_L g10575 ( 
.A1(n_9788),
.A2(n_8671),
.B1(n_8628),
.B2(n_8122),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_9113),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_9116),
.Y(n_10577)
);

INVx1_ASAP7_75t_L g10578 ( 
.A(n_9116),
.Y(n_10578)
);

INVx1_ASAP7_75t_L g10579 ( 
.A(n_9124),
.Y(n_10579)
);

INVx2_ASAP7_75t_SL g10580 ( 
.A(n_9514),
.Y(n_10580)
);

NAND2xp5_ASAP7_75t_L g10581 ( 
.A(n_9158),
.B(n_8402),
.Y(n_10581)
);

INVx1_ASAP7_75t_L g10582 ( 
.A(n_9124),
.Y(n_10582)
);

OAI21x1_ASAP7_75t_L g10583 ( 
.A1(n_9070),
.A2(n_8077),
.B(n_8826),
.Y(n_10583)
);

INVx1_ASAP7_75t_L g10584 ( 
.A(n_9129),
.Y(n_10584)
);

OAI21x1_ASAP7_75t_L g10585 ( 
.A1(n_9070),
.A2(n_7845),
.B(n_8072),
.Y(n_10585)
);

A2O1A1Ixp33_ASAP7_75t_L g10586 ( 
.A1(n_9039),
.A2(n_8639),
.B(n_8319),
.C(n_8071),
.Y(n_10586)
);

OAI21x1_ASAP7_75t_L g10587 ( 
.A1(n_9154),
.A2(n_7845),
.B(n_8072),
.Y(n_10587)
);

INVx1_ASAP7_75t_L g10588 ( 
.A(n_9129),
.Y(n_10588)
);

OA21x2_ASAP7_75t_L g10589 ( 
.A1(n_10089),
.A2(n_8990),
.B(n_8985),
.Y(n_10589)
);

INVx1_ASAP7_75t_L g10590 ( 
.A(n_9138),
.Y(n_10590)
);

INVx1_ASAP7_75t_L g10591 ( 
.A(n_9138),
.Y(n_10591)
);

INVx4_ASAP7_75t_L g10592 ( 
.A(n_9098),
.Y(n_10592)
);

INVx2_ASAP7_75t_L g10593 ( 
.A(n_9576),
.Y(n_10593)
);

OAI21x1_ASAP7_75t_L g10594 ( 
.A1(n_9154),
.A2(n_7845),
.B(n_8072),
.Y(n_10594)
);

OAI21x1_ASAP7_75t_L g10595 ( 
.A1(n_9194),
.A2(n_8816),
.B(n_8991),
.Y(n_10595)
);

AND2x2_ASAP7_75t_L g10596 ( 
.A(n_9850),
.B(n_8468),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_9139),
.Y(n_10597)
);

OAI22xp5_ASAP7_75t_L g10598 ( 
.A1(n_9358),
.A2(n_8671),
.B1(n_8122),
.B2(n_8793),
.Y(n_10598)
);

INVx6_ASAP7_75t_L g10599 ( 
.A(n_9471),
.Y(n_10599)
);

BUFx3_ASAP7_75t_L g10600 ( 
.A(n_9503),
.Y(n_10600)
);

INVx2_ASAP7_75t_L g10601 ( 
.A(n_9576),
.Y(n_10601)
);

NOR2xp33_ASAP7_75t_L g10602 ( 
.A(n_9067),
.B(n_8531),
.Y(n_10602)
);

INVx1_ASAP7_75t_L g10603 ( 
.A(n_9139),
.Y(n_10603)
);

BUFx2_ASAP7_75t_L g10604 ( 
.A(n_9444),
.Y(n_10604)
);

INVx1_ASAP7_75t_L g10605 ( 
.A(n_9150),
.Y(n_10605)
);

INVx2_ASAP7_75t_L g10606 ( 
.A(n_9577),
.Y(n_10606)
);

INVx1_ASAP7_75t_L g10607 ( 
.A(n_9150),
.Y(n_10607)
);

HB1xp67_ASAP7_75t_L g10608 ( 
.A(n_10183),
.Y(n_10608)
);

INVx1_ASAP7_75t_L g10609 ( 
.A(n_9151),
.Y(n_10609)
);

INVx2_ASAP7_75t_L g10610 ( 
.A(n_9577),
.Y(n_10610)
);

INVx2_ASAP7_75t_L g10611 ( 
.A(n_9577),
.Y(n_10611)
);

CKINVDCx5p33_ASAP7_75t_R g10612 ( 
.A(n_9503),
.Y(n_10612)
);

BUFx6f_ASAP7_75t_L g10613 ( 
.A(n_9098),
.Y(n_10613)
);

BUFx2_ASAP7_75t_L g10614 ( 
.A(n_9444),
.Y(n_10614)
);

BUFx2_ASAP7_75t_L g10615 ( 
.A(n_9444),
.Y(n_10615)
);

HB1xp67_ASAP7_75t_L g10616 ( 
.A(n_10254),
.Y(n_10616)
);

AOI221xp5_ASAP7_75t_L g10617 ( 
.A1(n_9557),
.A2(n_8825),
.B1(n_8654),
.B2(n_8688),
.C(n_7882),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_9151),
.Y(n_10618)
);

INVx1_ASAP7_75t_L g10619 ( 
.A(n_9153),
.Y(n_10619)
);

AND2x4_ASAP7_75t_L g10620 ( 
.A(n_9950),
.B(n_7719),
.Y(n_10620)
);

AND2x2_ASAP7_75t_L g10621 ( 
.A(n_9886),
.B(n_8468),
.Y(n_10621)
);

INVxp67_ASAP7_75t_L g10622 ( 
.A(n_9386),
.Y(n_10622)
);

BUFx6f_ASAP7_75t_L g10623 ( 
.A(n_9098),
.Y(n_10623)
);

OAI21xp5_ASAP7_75t_L g10624 ( 
.A1(n_9535),
.A2(n_8633),
.B(n_7909),
.Y(n_10624)
);

INVx2_ASAP7_75t_L g10625 ( 
.A(n_9589),
.Y(n_10625)
);

INVx1_ASAP7_75t_L g10626 ( 
.A(n_9153),
.Y(n_10626)
);

INVx1_ASAP7_75t_L g10627 ( 
.A(n_9168),
.Y(n_10627)
);

BUFx2_ASAP7_75t_L g10628 ( 
.A(n_10148),
.Y(n_10628)
);

INVx1_ASAP7_75t_L g10629 ( 
.A(n_9168),
.Y(n_10629)
);

INVx2_ASAP7_75t_L g10630 ( 
.A(n_9589),
.Y(n_10630)
);

INVx2_ASAP7_75t_L g10631 ( 
.A(n_9589),
.Y(n_10631)
);

INVx8_ASAP7_75t_L g10632 ( 
.A(n_9136),
.Y(n_10632)
);

OR2x2_ASAP7_75t_L g10633 ( 
.A(n_9615),
.B(n_8076),
.Y(n_10633)
);

BUFx3_ASAP7_75t_L g10634 ( 
.A(n_9503),
.Y(n_10634)
);

BUFx3_ASAP7_75t_L g10635 ( 
.A(n_9503),
.Y(n_10635)
);

INVx1_ASAP7_75t_L g10636 ( 
.A(n_9169),
.Y(n_10636)
);

INVx1_ASAP7_75t_L g10637 ( 
.A(n_9169),
.Y(n_10637)
);

INVx2_ASAP7_75t_L g10638 ( 
.A(n_9592),
.Y(n_10638)
);

INVx1_ASAP7_75t_L g10639 ( 
.A(n_9176),
.Y(n_10639)
);

NAND2xp5_ASAP7_75t_L g10640 ( 
.A(n_9170),
.B(n_8402),
.Y(n_10640)
);

AOI22xp33_ASAP7_75t_L g10641 ( 
.A1(n_9348),
.A2(n_7810),
.B1(n_8899),
.B2(n_8836),
.Y(n_10641)
);

OAI31xp33_ASAP7_75t_SL g10642 ( 
.A1(n_9536),
.A2(n_8670),
.A3(n_8754),
.B(n_8708),
.Y(n_10642)
);

INVx2_ASAP7_75t_L g10643 ( 
.A(n_9592),
.Y(n_10643)
);

AOI22xp33_ASAP7_75t_SL g10644 ( 
.A1(n_10265),
.A2(n_7810),
.B1(n_7796),
.B2(n_8332),
.Y(n_10644)
);

INVx2_ASAP7_75t_L g10645 ( 
.A(n_9592),
.Y(n_10645)
);

INVx1_ASAP7_75t_L g10646 ( 
.A(n_9176),
.Y(n_10646)
);

INVx2_ASAP7_75t_L g10647 ( 
.A(n_9594),
.Y(n_10647)
);

INVx4_ASAP7_75t_SL g10648 ( 
.A(n_9098),
.Y(n_10648)
);

OAI22xp5_ASAP7_75t_L g10649 ( 
.A1(n_10246),
.A2(n_8793),
.B1(n_8653),
.B2(n_8385),
.Y(n_10649)
);

INVx1_ASAP7_75t_L g10650 ( 
.A(n_9177),
.Y(n_10650)
);

AND2x2_ASAP7_75t_L g10651 ( 
.A(n_9886),
.B(n_8468),
.Y(n_10651)
);

BUFx3_ASAP7_75t_L g10652 ( 
.A(n_9601),
.Y(n_10652)
);

INVx1_ASAP7_75t_L g10653 ( 
.A(n_9177),
.Y(n_10653)
);

INVx2_ASAP7_75t_L g10654 ( 
.A(n_9594),
.Y(n_10654)
);

BUFx3_ASAP7_75t_L g10655 ( 
.A(n_9601),
.Y(n_10655)
);

OR2x2_ASAP7_75t_L g10656 ( 
.A(n_9108),
.B(n_9112),
.Y(n_10656)
);

AND2x4_ASAP7_75t_L g10657 ( 
.A(n_9950),
.B(n_7719),
.Y(n_10657)
);

HB1xp67_ASAP7_75t_L g10658 ( 
.A(n_10282),
.Y(n_10658)
);

INVx1_ASAP7_75t_L g10659 ( 
.A(n_9178),
.Y(n_10659)
);

AND2x4_ASAP7_75t_L g10660 ( 
.A(n_9950),
.B(n_7719),
.Y(n_10660)
);

BUFx3_ASAP7_75t_L g10661 ( 
.A(n_9601),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_9178),
.Y(n_10662)
);

INVx3_ASAP7_75t_L g10663 ( 
.A(n_9514),
.Y(n_10663)
);

INVx1_ASAP7_75t_L g10664 ( 
.A(n_9183),
.Y(n_10664)
);

INVx1_ASAP7_75t_L g10665 ( 
.A(n_9183),
.Y(n_10665)
);

INVx1_ASAP7_75t_L g10666 ( 
.A(n_9184),
.Y(n_10666)
);

OAI211xp5_ASAP7_75t_L g10667 ( 
.A1(n_10284),
.A2(n_7824),
.B(n_7796),
.C(n_9025),
.Y(n_10667)
);

INVx1_ASAP7_75t_L g10668 ( 
.A(n_9184),
.Y(n_10668)
);

INVx1_ASAP7_75t_L g10669 ( 
.A(n_9185),
.Y(n_10669)
);

AOI22xp33_ASAP7_75t_SL g10670 ( 
.A1(n_10265),
.A2(n_7810),
.B1(n_7796),
.B2(n_7882),
.Y(n_10670)
);

AND2x4_ASAP7_75t_L g10671 ( 
.A(n_9959),
.B(n_7881),
.Y(n_10671)
);

AND2x4_ASAP7_75t_L g10672 ( 
.A(n_9959),
.B(n_7881),
.Y(n_10672)
);

INVx2_ASAP7_75t_L g10673 ( 
.A(n_9594),
.Y(n_10673)
);

HB1xp67_ASAP7_75t_L g10674 ( 
.A(n_9088),
.Y(n_10674)
);

AOI22xp33_ASAP7_75t_L g10675 ( 
.A1(n_9349),
.A2(n_7810),
.B1(n_8899),
.B2(n_8836),
.Y(n_10675)
);

BUFx2_ASAP7_75t_L g10676 ( 
.A(n_10148),
.Y(n_10676)
);

OR2x2_ASAP7_75t_L g10677 ( 
.A(n_9108),
.B(n_8076),
.Y(n_10677)
);

INVx1_ASAP7_75t_L g10678 ( 
.A(n_9185),
.Y(n_10678)
);

AND2x2_ASAP7_75t_L g10679 ( 
.A(n_9081),
.B(n_8524),
.Y(n_10679)
);

BUFx2_ASAP7_75t_L g10680 ( 
.A(n_10148),
.Y(n_10680)
);

INVx2_ASAP7_75t_L g10681 ( 
.A(n_9598),
.Y(n_10681)
);

INVx1_ASAP7_75t_L g10682 ( 
.A(n_9187),
.Y(n_10682)
);

INVx3_ASAP7_75t_L g10683 ( 
.A(n_9514),
.Y(n_10683)
);

INVx1_ASAP7_75t_L g10684 ( 
.A(n_9187),
.Y(n_10684)
);

INVx3_ASAP7_75t_L g10685 ( 
.A(n_9547),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_9191),
.Y(n_10686)
);

INVx3_ASAP7_75t_L g10687 ( 
.A(n_9547),
.Y(n_10687)
);

INVx2_ASAP7_75t_L g10688 ( 
.A(n_9598),
.Y(n_10688)
);

OAI21x1_ASAP7_75t_L g10689 ( 
.A1(n_9194),
.A2(n_8816),
.B(n_8991),
.Y(n_10689)
);

INVx2_ASAP7_75t_L g10690 ( 
.A(n_9598),
.Y(n_10690)
);

OR2x6_ASAP7_75t_L g10691 ( 
.A(n_9380),
.B(n_9959),
.Y(n_10691)
);

INVx3_ASAP7_75t_L g10692 ( 
.A(n_9547),
.Y(n_10692)
);

INVx1_ASAP7_75t_L g10693 ( 
.A(n_9191),
.Y(n_10693)
);

INVx4_ASAP7_75t_L g10694 ( 
.A(n_9100),
.Y(n_10694)
);

INVx1_ASAP7_75t_L g10695 ( 
.A(n_9197),
.Y(n_10695)
);

OR2x2_ASAP7_75t_L g10696 ( 
.A(n_9112),
.B(n_8430),
.Y(n_10696)
);

NAND2xp5_ASAP7_75t_L g10697 ( 
.A(n_9172),
.B(n_8541),
.Y(n_10697)
);

INVx1_ASAP7_75t_L g10698 ( 
.A(n_9197),
.Y(n_10698)
);

INVx2_ASAP7_75t_L g10699 ( 
.A(n_9600),
.Y(n_10699)
);

AND2x2_ASAP7_75t_L g10700 ( 
.A(n_9081),
.B(n_8524),
.Y(n_10700)
);

INVx3_ASAP7_75t_L g10701 ( 
.A(n_9547),
.Y(n_10701)
);

CKINVDCx20_ASAP7_75t_R g10702 ( 
.A(n_9442),
.Y(n_10702)
);

BUFx6f_ASAP7_75t_L g10703 ( 
.A(n_9100),
.Y(n_10703)
);

INVx2_ASAP7_75t_L g10704 ( 
.A(n_9600),
.Y(n_10704)
);

INVx2_ASAP7_75t_L g10705 ( 
.A(n_9600),
.Y(n_10705)
);

INVx1_ASAP7_75t_L g10706 ( 
.A(n_9202),
.Y(n_10706)
);

INVx1_ASAP7_75t_L g10707 ( 
.A(n_9202),
.Y(n_10707)
);

AOI21xp5_ASAP7_75t_L g10708 ( 
.A1(n_9483),
.A2(n_7776),
.B(n_7791),
.Y(n_10708)
);

INVx2_ASAP7_75t_L g10709 ( 
.A(n_9605),
.Y(n_10709)
);

INVx2_ASAP7_75t_L g10710 ( 
.A(n_9605),
.Y(n_10710)
);

OAI21x1_ASAP7_75t_L g10711 ( 
.A1(n_9325),
.A2(n_9017),
.B(n_8991),
.Y(n_10711)
);

INVx1_ASAP7_75t_L g10712 ( 
.A(n_9208),
.Y(n_10712)
);

INVx2_ASAP7_75t_L g10713 ( 
.A(n_9605),
.Y(n_10713)
);

INVx1_ASAP7_75t_L g10714 ( 
.A(n_9208),
.Y(n_10714)
);

NAND2x1p5_ASAP7_75t_L g10715 ( 
.A(n_9547),
.B(n_8805),
.Y(n_10715)
);

BUFx3_ASAP7_75t_L g10716 ( 
.A(n_9601),
.Y(n_10716)
);

NAND2xp5_ASAP7_75t_L g10717 ( 
.A(n_9172),
.B(n_8541),
.Y(n_10717)
);

INVx2_ASAP7_75t_L g10718 ( 
.A(n_9606),
.Y(n_10718)
);

AO21x2_ASAP7_75t_L g10719 ( 
.A1(n_9565),
.A2(n_7906),
.B(n_8416),
.Y(n_10719)
);

INVx2_ASAP7_75t_L g10720 ( 
.A(n_9606),
.Y(n_10720)
);

INVx1_ASAP7_75t_L g10721 ( 
.A(n_9213),
.Y(n_10721)
);

AND2x2_ASAP7_75t_L g10722 ( 
.A(n_9081),
.B(n_8524),
.Y(n_10722)
);

INVx2_ASAP7_75t_L g10723 ( 
.A(n_9606),
.Y(n_10723)
);

INVx1_ASAP7_75t_L g10724 ( 
.A(n_9213),
.Y(n_10724)
);

HB1xp67_ASAP7_75t_L g10725 ( 
.A(n_9090),
.Y(n_10725)
);

INVx1_ASAP7_75t_L g10726 ( 
.A(n_9217),
.Y(n_10726)
);

INVxp67_ASAP7_75t_L g10727 ( 
.A(n_9519),
.Y(n_10727)
);

AND2x2_ASAP7_75t_L g10728 ( 
.A(n_9081),
.B(n_8549),
.Y(n_10728)
);

INVx1_ASAP7_75t_L g10729 ( 
.A(n_9217),
.Y(n_10729)
);

INVx2_ASAP7_75t_L g10730 ( 
.A(n_9610),
.Y(n_10730)
);

INVx3_ASAP7_75t_L g10731 ( 
.A(n_9547),
.Y(n_10731)
);

INVx2_ASAP7_75t_L g10732 ( 
.A(n_9610),
.Y(n_10732)
);

AOI22xp33_ASAP7_75t_L g10733 ( 
.A1(n_9349),
.A2(n_8791),
.B1(n_7808),
.B2(n_7785),
.Y(n_10733)
);

CKINVDCx16_ASAP7_75t_R g10734 ( 
.A(n_10088),
.Y(n_10734)
);

OAI21x1_ASAP7_75t_L g10735 ( 
.A1(n_9325),
.A2(n_9017),
.B(n_8534),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_9218),
.Y(n_10736)
);

INVx1_ASAP7_75t_L g10737 ( 
.A(n_9218),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_9220),
.Y(n_10738)
);

INVx1_ASAP7_75t_L g10739 ( 
.A(n_9220),
.Y(n_10739)
);

AO31x2_ASAP7_75t_L g10740 ( 
.A1(n_9949),
.A2(n_8416),
.A3(n_8300),
.B(n_7955),
.Y(n_10740)
);

AND2x2_ASAP7_75t_L g10741 ( 
.A(n_9095),
.B(n_8549),
.Y(n_10741)
);

AND2x4_ASAP7_75t_L g10742 ( 
.A(n_9959),
.B(n_7881),
.Y(n_10742)
);

INVx1_ASAP7_75t_L g10743 ( 
.A(n_9225),
.Y(n_10743)
);

INVx3_ASAP7_75t_L g10744 ( 
.A(n_9547),
.Y(n_10744)
);

BUFx3_ASAP7_75t_L g10745 ( 
.A(n_10003),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_9225),
.Y(n_10746)
);

INVx2_ASAP7_75t_L g10747 ( 
.A(n_9610),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_9233),
.Y(n_10748)
);

AND2x2_ASAP7_75t_L g10749 ( 
.A(n_9095),
.B(n_8549),
.Y(n_10749)
);

OR2x2_ASAP7_75t_L g10750 ( 
.A(n_9120),
.B(n_8430),
.Y(n_10750)
);

HB1xp67_ASAP7_75t_L g10751 ( 
.A(n_9102),
.Y(n_10751)
);

INVx1_ASAP7_75t_L g10752 ( 
.A(n_9233),
.Y(n_10752)
);

INVx1_ASAP7_75t_L g10753 ( 
.A(n_9239),
.Y(n_10753)
);

INVx1_ASAP7_75t_L g10754 ( 
.A(n_9239),
.Y(n_10754)
);

INVx2_ASAP7_75t_L g10755 ( 
.A(n_9614),
.Y(n_10755)
);

INVx2_ASAP7_75t_L g10756 ( 
.A(n_9614),
.Y(n_10756)
);

NOR2x1_ASAP7_75t_SL g10757 ( 
.A(n_9518),
.B(n_8766),
.Y(n_10757)
);

INVx1_ASAP7_75t_L g10758 ( 
.A(n_9243),
.Y(n_10758)
);

INVx1_ASAP7_75t_L g10759 ( 
.A(n_9243),
.Y(n_10759)
);

INVx2_ASAP7_75t_SL g10760 ( 
.A(n_9591),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_9614),
.Y(n_10761)
);

INVx2_ASAP7_75t_L g10762 ( 
.A(n_9620),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_9244),
.Y(n_10763)
);

OR2x2_ASAP7_75t_L g10764 ( 
.A(n_9120),
.B(n_8430),
.Y(n_10764)
);

OR2x6_ASAP7_75t_L g10765 ( 
.A(n_9380),
.B(n_8531),
.Y(n_10765)
);

INVx2_ASAP7_75t_L g10766 ( 
.A(n_9620),
.Y(n_10766)
);

AO21x2_ASAP7_75t_L g10767 ( 
.A1(n_9565),
.A2(n_7906),
.B(n_7824),
.Y(n_10767)
);

INVx2_ASAP7_75t_SL g10768 ( 
.A(n_10210),
.Y(n_10768)
);

INVx3_ASAP7_75t_L g10769 ( 
.A(n_9591),
.Y(n_10769)
);

OAI21x1_ASAP7_75t_L g10770 ( 
.A1(n_9325),
.A2(n_9017),
.B(n_8534),
.Y(n_10770)
);

OR2x2_ASAP7_75t_L g10771 ( 
.A(n_9143),
.B(n_8484),
.Y(n_10771)
);

INVx2_ASAP7_75t_L g10772 ( 
.A(n_9620),
.Y(n_10772)
);

INVx1_ASAP7_75t_L g10773 ( 
.A(n_9244),
.Y(n_10773)
);

INVx1_ASAP7_75t_L g10774 ( 
.A(n_9247),
.Y(n_10774)
);

AND2x2_ASAP7_75t_L g10775 ( 
.A(n_9095),
.B(n_9141),
.Y(n_10775)
);

INVx1_ASAP7_75t_L g10776 ( 
.A(n_9247),
.Y(n_10776)
);

INVx2_ASAP7_75t_L g10777 ( 
.A(n_9622),
.Y(n_10777)
);

INVx1_ASAP7_75t_L g10778 ( 
.A(n_9248),
.Y(n_10778)
);

INVx2_ASAP7_75t_L g10779 ( 
.A(n_9622),
.Y(n_10779)
);

OR2x2_ASAP7_75t_L g10780 ( 
.A(n_9143),
.B(n_8484),
.Y(n_10780)
);

OAI22xp5_ASAP7_75t_L g10781 ( 
.A1(n_10024),
.A2(n_8653),
.B1(n_8385),
.B2(n_8406),
.Y(n_10781)
);

INVx1_ASAP7_75t_L g10782 ( 
.A(n_9248),
.Y(n_10782)
);

INVx1_ASAP7_75t_L g10783 ( 
.A(n_9251),
.Y(n_10783)
);

OR2x2_ASAP7_75t_L g10784 ( 
.A(n_9324),
.B(n_8185),
.Y(n_10784)
);

AOI21x1_ASAP7_75t_L g10785 ( 
.A1(n_9374),
.A2(n_8213),
.B(n_8190),
.Y(n_10785)
);

HB1xp67_ASAP7_75t_L g10786 ( 
.A(n_9133),
.Y(n_10786)
);

AND2x2_ASAP7_75t_L g10787 ( 
.A(n_9095),
.B(n_8588),
.Y(n_10787)
);

INVx1_ASAP7_75t_L g10788 ( 
.A(n_9251),
.Y(n_10788)
);

INVx1_ASAP7_75t_L g10789 ( 
.A(n_9253),
.Y(n_10789)
);

HB1xp67_ASAP7_75t_L g10790 ( 
.A(n_9164),
.Y(n_10790)
);

AND2x6_ASAP7_75t_L g10791 ( 
.A(n_9288),
.B(n_8282),
.Y(n_10791)
);

HB1xp67_ASAP7_75t_L g10792 ( 
.A(n_9181),
.Y(n_10792)
);

OR2x2_ASAP7_75t_L g10793 ( 
.A(n_9324),
.B(n_8213),
.Y(n_10793)
);

AND2x2_ASAP7_75t_L g10794 ( 
.A(n_9141),
.B(n_8588),
.Y(n_10794)
);

INVx2_ASAP7_75t_SL g10795 ( 
.A(n_10268),
.Y(n_10795)
);

INVx2_ASAP7_75t_L g10796 ( 
.A(n_9622),
.Y(n_10796)
);

HB1xp67_ASAP7_75t_L g10797 ( 
.A(n_9200),
.Y(n_10797)
);

HB1xp67_ASAP7_75t_L g10798 ( 
.A(n_9214),
.Y(n_10798)
);

INVx2_ASAP7_75t_L g10799 ( 
.A(n_9635),
.Y(n_10799)
);

INVx1_ASAP7_75t_L g10800 ( 
.A(n_9253),
.Y(n_10800)
);

INVx1_ASAP7_75t_L g10801 ( 
.A(n_9259),
.Y(n_10801)
);

OR2x2_ASAP7_75t_L g10802 ( 
.A(n_9142),
.B(n_8489),
.Y(n_10802)
);

INVx1_ASAP7_75t_SL g10803 ( 
.A(n_9551),
.Y(n_10803)
);

INVx1_ASAP7_75t_L g10804 ( 
.A(n_9259),
.Y(n_10804)
);

OR2x6_ASAP7_75t_L g10805 ( 
.A(n_9980),
.B(n_8531),
.Y(n_10805)
);

INVx4_ASAP7_75t_SL g10806 ( 
.A(n_9100),
.Y(n_10806)
);

INVx1_ASAP7_75t_L g10807 ( 
.A(n_9271),
.Y(n_10807)
);

BUFx2_ASAP7_75t_L g10808 ( 
.A(n_10148),
.Y(n_10808)
);

BUFx3_ASAP7_75t_L g10809 ( 
.A(n_10003),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_9271),
.Y(n_10810)
);

NAND2x1p5_ASAP7_75t_L g10811 ( 
.A(n_9591),
.B(n_8805),
.Y(n_10811)
);

INVx1_ASAP7_75t_L g10812 ( 
.A(n_9272),
.Y(n_10812)
);

OAI21xp5_ASAP7_75t_L g10813 ( 
.A1(n_9483),
.A2(n_8633),
.B(n_7909),
.Y(n_10813)
);

INVx1_ASAP7_75t_L g10814 ( 
.A(n_9272),
.Y(n_10814)
);

HB1xp67_ASAP7_75t_L g10815 ( 
.A(n_9224),
.Y(n_10815)
);

AND2x2_ASAP7_75t_L g10816 ( 
.A(n_9141),
.B(n_8588),
.Y(n_10816)
);

INVx2_ASAP7_75t_L g10817 ( 
.A(n_9635),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_9293),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_9293),
.Y(n_10819)
);

INVx1_ASAP7_75t_L g10820 ( 
.A(n_9294),
.Y(n_10820)
);

INVx1_ASAP7_75t_L g10821 ( 
.A(n_9294),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_9299),
.Y(n_10822)
);

INVx3_ASAP7_75t_L g10823 ( 
.A(n_9591),
.Y(n_10823)
);

HB1xp67_ASAP7_75t_L g10824 ( 
.A(n_9246),
.Y(n_10824)
);

AOI22xp33_ASAP7_75t_L g10825 ( 
.A1(n_9354),
.A2(n_8791),
.B1(n_7808),
.B2(n_7785),
.Y(n_10825)
);

AOI21x1_ASAP7_75t_L g10826 ( 
.A1(n_9205),
.A2(n_7955),
.B(n_7882),
.Y(n_10826)
);

OAI21x1_ASAP7_75t_L g10827 ( 
.A1(n_9458),
.A2(n_8534),
.B(n_8372),
.Y(n_10827)
);

INVx2_ASAP7_75t_L g10828 ( 
.A(n_9635),
.Y(n_10828)
);

HB1xp67_ASAP7_75t_L g10829 ( 
.A(n_9260),
.Y(n_10829)
);

BUFx6f_ASAP7_75t_L g10830 ( 
.A(n_9100),
.Y(n_10830)
);

INVx2_ASAP7_75t_L g10831 ( 
.A(n_9636),
.Y(n_10831)
);

AND2x2_ASAP7_75t_L g10832 ( 
.A(n_9141),
.B(n_8615),
.Y(n_10832)
);

AOI22xp5_ASAP7_75t_L g10833 ( 
.A1(n_10229),
.A2(n_7773),
.B1(n_8754),
.B2(n_8708),
.Y(n_10833)
);

AND2x2_ASAP7_75t_L g10834 ( 
.A(n_9147),
.B(n_8615),
.Y(n_10834)
);

AND2x4_ASAP7_75t_L g10835 ( 
.A(n_9980),
.B(n_9925),
.Y(n_10835)
);

INVx2_ASAP7_75t_L g10836 ( 
.A(n_9636),
.Y(n_10836)
);

INVx2_ASAP7_75t_L g10837 ( 
.A(n_9636),
.Y(n_10837)
);

AND2x2_ASAP7_75t_L g10838 ( 
.A(n_9147),
.B(n_9125),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_9966),
.B(n_10114),
.Y(n_10839)
);

INVx4_ASAP7_75t_L g10840 ( 
.A(n_9100),
.Y(n_10840)
);

INVx2_ASAP7_75t_L g10841 ( 
.A(n_9664),
.Y(n_10841)
);

INVx1_ASAP7_75t_L g10842 ( 
.A(n_9299),
.Y(n_10842)
);

INVx2_ASAP7_75t_L g10843 ( 
.A(n_9664),
.Y(n_10843)
);

INVx3_ASAP7_75t_L g10844 ( 
.A(n_9591),
.Y(n_10844)
);

HB1xp67_ASAP7_75t_L g10845 ( 
.A(n_9333),
.Y(n_10845)
);

HB1xp67_ASAP7_75t_L g10846 ( 
.A(n_9336),
.Y(n_10846)
);

HB1xp67_ASAP7_75t_L g10847 ( 
.A(n_9384),
.Y(n_10847)
);

INVx2_ASAP7_75t_L g10848 ( 
.A(n_9664),
.Y(n_10848)
);

HB1xp67_ASAP7_75t_L g10849 ( 
.A(n_9413),
.Y(n_10849)
);

INVx1_ASAP7_75t_L g10850 ( 
.A(n_9301),
.Y(n_10850)
);

BUFx2_ASAP7_75t_L g10851 ( 
.A(n_10157),
.Y(n_10851)
);

INVx2_ASAP7_75t_L g10852 ( 
.A(n_9665),
.Y(n_10852)
);

BUFx2_ASAP7_75t_L g10853 ( 
.A(n_10157),
.Y(n_10853)
);

INVx2_ASAP7_75t_L g10854 ( 
.A(n_9665),
.Y(n_10854)
);

OA21x2_ASAP7_75t_L g10855 ( 
.A1(n_10089),
.A2(n_9720),
.B(n_10149),
.Y(n_10855)
);

NAND2xp5_ASAP7_75t_SL g10856 ( 
.A(n_10278),
.B(n_8071),
.Y(n_10856)
);

INVx2_ASAP7_75t_SL g10857 ( 
.A(n_9591),
.Y(n_10857)
);

INVx2_ASAP7_75t_SL g10858 ( 
.A(n_10210),
.Y(n_10858)
);

AO21x2_ASAP7_75t_L g10859 ( 
.A1(n_9613),
.A2(n_7906),
.B(n_7824),
.Y(n_10859)
);

INVx2_ASAP7_75t_L g10860 ( 
.A(n_9665),
.Y(n_10860)
);

BUFx6f_ASAP7_75t_L g10861 ( 
.A(n_9100),
.Y(n_10861)
);

INVx2_ASAP7_75t_SL g10862 ( 
.A(n_10048),
.Y(n_10862)
);

INVx2_ASAP7_75t_L g10863 ( 
.A(n_9694),
.Y(n_10863)
);

BUFx6f_ASAP7_75t_L g10864 ( 
.A(n_9130),
.Y(n_10864)
);

INVx2_ASAP7_75t_L g10865 ( 
.A(n_9694),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_9301),
.Y(n_10866)
);

INVx1_ASAP7_75t_L g10867 ( 
.A(n_9306),
.Y(n_10867)
);

INVx1_ASAP7_75t_L g10868 ( 
.A(n_9306),
.Y(n_10868)
);

NAND2xp5_ASAP7_75t_L g10869 ( 
.A(n_9354),
.B(n_8554),
.Y(n_10869)
);

AOI21xp5_ASAP7_75t_L g10870 ( 
.A1(n_9528),
.A2(n_7791),
.B(n_8629),
.Y(n_10870)
);

INVx1_ASAP7_75t_L g10871 ( 
.A(n_9311),
.Y(n_10871)
);

OR2x6_ASAP7_75t_L g10872 ( 
.A(n_9980),
.B(n_8761),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_9311),
.Y(n_10873)
);

INVx2_ASAP7_75t_L g10874 ( 
.A(n_9694),
.Y(n_10874)
);

INVx1_ASAP7_75t_L g10875 ( 
.A(n_9316),
.Y(n_10875)
);

AND2x2_ASAP7_75t_L g10876 ( 
.A(n_9147),
.B(n_8615),
.Y(n_10876)
);

AND2x2_ASAP7_75t_L g10877 ( 
.A(n_9147),
.B(n_8635),
.Y(n_10877)
);

INVx2_ASAP7_75t_L g10878 ( 
.A(n_9697),
.Y(n_10878)
);

AND2x4_ASAP7_75t_L g10879 ( 
.A(n_9980),
.B(n_7881),
.Y(n_10879)
);

HB1xp67_ASAP7_75t_L g10880 ( 
.A(n_9422),
.Y(n_10880)
);

HB1xp67_ASAP7_75t_L g10881 ( 
.A(n_9436),
.Y(n_10881)
);

INVx2_ASAP7_75t_L g10882 ( 
.A(n_9697),
.Y(n_10882)
);

BUFx6f_ASAP7_75t_L g10883 ( 
.A(n_9130),
.Y(n_10883)
);

INVx1_ASAP7_75t_L g10884 ( 
.A(n_9316),
.Y(n_10884)
);

BUFx3_ASAP7_75t_L g10885 ( 
.A(n_10003),
.Y(n_10885)
);

BUFx4f_ASAP7_75t_SL g10886 ( 
.A(n_9211),
.Y(n_10886)
);

OR2x2_ASAP7_75t_L g10887 ( 
.A(n_9142),
.B(n_8489),
.Y(n_10887)
);

AO21x2_ASAP7_75t_L g10888 ( 
.A1(n_9613),
.A2(n_8757),
.B(n_8749),
.Y(n_10888)
);

OAI21x1_ASAP7_75t_L g10889 ( 
.A1(n_9458),
.A2(n_8372),
.B(n_8118),
.Y(n_10889)
);

INVx1_ASAP7_75t_L g10890 ( 
.A(n_9320),
.Y(n_10890)
);

AND2x2_ASAP7_75t_L g10891 ( 
.A(n_9125),
.B(n_8635),
.Y(n_10891)
);

HB1xp67_ASAP7_75t_L g10892 ( 
.A(n_9451),
.Y(n_10892)
);

HB1xp67_ASAP7_75t_L g10893 ( 
.A(n_9452),
.Y(n_10893)
);

INVx1_ASAP7_75t_L g10894 ( 
.A(n_9320),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_9322),
.Y(n_10895)
);

INVx2_ASAP7_75t_L g10896 ( 
.A(n_9697),
.Y(n_10896)
);

INVx1_ASAP7_75t_L g10897 ( 
.A(n_9322),
.Y(n_10897)
);

BUFx2_ASAP7_75t_L g10898 ( 
.A(n_10157),
.Y(n_10898)
);

INVx2_ASAP7_75t_L g10899 ( 
.A(n_9698),
.Y(n_10899)
);

BUFx4f_ASAP7_75t_SL g10900 ( 
.A(n_9211),
.Y(n_10900)
);

INVx3_ASAP7_75t_L g10901 ( 
.A(n_10048),
.Y(n_10901)
);

AND2x4_ASAP7_75t_L g10902 ( 
.A(n_9925),
.B(n_7905),
.Y(n_10902)
);

INVx2_ASAP7_75t_L g10903 ( 
.A(n_9698),
.Y(n_10903)
);

BUFx2_ASAP7_75t_L g10904 ( 
.A(n_10157),
.Y(n_10904)
);

OAI21xp5_ASAP7_75t_L g10905 ( 
.A1(n_10093),
.A2(n_7909),
.B(n_7902),
.Y(n_10905)
);

INVx2_ASAP7_75t_SL g10906 ( 
.A(n_10048),
.Y(n_10906)
);

INVx1_ASAP7_75t_L g10907 ( 
.A(n_9323),
.Y(n_10907)
);

INVx1_ASAP7_75t_L g10908 ( 
.A(n_9323),
.Y(n_10908)
);

OAI21x1_ASAP7_75t_L g10909 ( 
.A1(n_9458),
.A2(n_8372),
.B(n_8118),
.Y(n_10909)
);

INVx2_ASAP7_75t_L g10910 ( 
.A(n_9698),
.Y(n_10910)
);

INVx1_ASAP7_75t_L g10911 ( 
.A(n_9327),
.Y(n_10911)
);

INVx1_ASAP7_75t_L g10912 ( 
.A(n_9327),
.Y(n_10912)
);

OR2x2_ASAP7_75t_L g10913 ( 
.A(n_9559),
.B(n_8495),
.Y(n_10913)
);

INVxp67_ASAP7_75t_L g10914 ( 
.A(n_10223),
.Y(n_10914)
);

BUFx2_ASAP7_75t_L g10915 ( 
.A(n_9429),
.Y(n_10915)
);

INVx1_ASAP7_75t_L g10916 ( 
.A(n_9331),
.Y(n_10916)
);

BUFx3_ASAP7_75t_L g10917 ( 
.A(n_10003),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_9331),
.Y(n_10918)
);

AND2x2_ASAP7_75t_L g10919 ( 
.A(n_9166),
.B(n_8635),
.Y(n_10919)
);

AO21x2_ASAP7_75t_L g10920 ( 
.A1(n_10278),
.A2(n_8757),
.B(n_8749),
.Y(n_10920)
);

NAND2xp5_ASAP7_75t_L g10921 ( 
.A(n_9858),
.B(n_8554),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_9339),
.Y(n_10922)
);

INVx1_ASAP7_75t_L g10923 ( 
.A(n_9339),
.Y(n_10923)
);

OAI21x1_ASAP7_75t_L g10924 ( 
.A1(n_9522),
.A2(n_9541),
.B(n_9534),
.Y(n_10924)
);

OAI21x1_ASAP7_75t_L g10925 ( 
.A1(n_9522),
.A2(n_8118),
.B(n_8106),
.Y(n_10925)
);

OAI221xp5_ASAP7_75t_L g10926 ( 
.A1(n_9532),
.A2(n_8453),
.B1(n_8406),
.B2(n_8382),
.C(n_8688),
.Y(n_10926)
);

INVx2_ASAP7_75t_L g10927 ( 
.A(n_9704),
.Y(n_10927)
);

INVx1_ASAP7_75t_L g10928 ( 
.A(n_9346),
.Y(n_10928)
);

INVx1_ASAP7_75t_L g10929 ( 
.A(n_9346),
.Y(n_10929)
);

OAI211xp5_ASAP7_75t_L g10930 ( 
.A1(n_9744),
.A2(n_7796),
.B(n_9025),
.C(n_8125),
.Y(n_10930)
);

INVx2_ASAP7_75t_L g10931 ( 
.A(n_9704),
.Y(n_10931)
);

INVx2_ASAP7_75t_L g10932 ( 
.A(n_9704),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_9366),
.Y(n_10933)
);

BUFx2_ASAP7_75t_L g10934 ( 
.A(n_9429),
.Y(n_10934)
);

INVx2_ASAP7_75t_L g10935 ( 
.A(n_9707),
.Y(n_10935)
);

INVx1_ASAP7_75t_L g10936 ( 
.A(n_9366),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_9367),
.Y(n_10937)
);

OR2x2_ASAP7_75t_L g10938 ( 
.A(n_9559),
.B(n_8495),
.Y(n_10938)
);

INVx2_ASAP7_75t_L g10939 ( 
.A(n_9707),
.Y(n_10939)
);

NOR2xp33_ASAP7_75t_L g10940 ( 
.A(n_9310),
.B(n_8761),
.Y(n_10940)
);

INVx2_ASAP7_75t_L g10941 ( 
.A(n_9707),
.Y(n_10941)
);

HB1xp67_ASAP7_75t_L g10942 ( 
.A(n_9473),
.Y(n_10942)
);

AND2x2_ASAP7_75t_L g10943 ( 
.A(n_9166),
.B(n_8638),
.Y(n_10943)
);

INVx2_ASAP7_75t_L g10944 ( 
.A(n_9734),
.Y(n_10944)
);

INVx3_ASAP7_75t_L g10945 ( 
.A(n_10048),
.Y(n_10945)
);

INVx2_ASAP7_75t_L g10946 ( 
.A(n_9734),
.Y(n_10946)
);

HB1xp67_ASAP7_75t_L g10947 ( 
.A(n_9521),
.Y(n_10947)
);

AOI22xp33_ASAP7_75t_L g10948 ( 
.A1(n_9375),
.A2(n_7808),
.B1(n_7785),
.B2(n_7843),
.Y(n_10948)
);

INVx1_ASAP7_75t_L g10949 ( 
.A(n_9367),
.Y(n_10949)
);

INVx2_ASAP7_75t_L g10950 ( 
.A(n_9734),
.Y(n_10950)
);

INVx2_ASAP7_75t_L g10951 ( 
.A(n_9742),
.Y(n_10951)
);

INVx2_ASAP7_75t_L g10952 ( 
.A(n_9742),
.Y(n_10952)
);

HB1xp67_ASAP7_75t_L g10953 ( 
.A(n_9531),
.Y(n_10953)
);

HB1xp67_ASAP7_75t_L g10954 ( 
.A(n_9570),
.Y(n_10954)
);

BUFx3_ASAP7_75t_L g10955 ( 
.A(n_10102),
.Y(n_10955)
);

AOI21x1_ASAP7_75t_L g10956 ( 
.A1(n_9205),
.A2(n_8154),
.B(n_7967),
.Y(n_10956)
);

INVx1_ASAP7_75t_L g10957 ( 
.A(n_9368),
.Y(n_10957)
);

INVxp67_ASAP7_75t_L g10958 ( 
.A(n_10223),
.Y(n_10958)
);

INVx1_ASAP7_75t_L g10959 ( 
.A(n_9368),
.Y(n_10959)
);

BUFx3_ASAP7_75t_L g10960 ( 
.A(n_10102),
.Y(n_10960)
);

INVx2_ASAP7_75t_L g10961 ( 
.A(n_9742),
.Y(n_10961)
);

INVx1_ASAP7_75t_L g10962 ( 
.A(n_9372),
.Y(n_10962)
);

INVx2_ASAP7_75t_L g10963 ( 
.A(n_9743),
.Y(n_10963)
);

AND2x4_ASAP7_75t_L g10964 ( 
.A(n_9925),
.B(n_7905),
.Y(n_10964)
);

INVx2_ASAP7_75t_L g10965 ( 
.A(n_9743),
.Y(n_10965)
);

AND2x2_ASAP7_75t_L g10966 ( 
.A(n_9221),
.B(n_8638),
.Y(n_10966)
);

INVx1_ASAP7_75t_L g10967 ( 
.A(n_9372),
.Y(n_10967)
);

INVx1_ASAP7_75t_L g10968 ( 
.A(n_9376),
.Y(n_10968)
);

INVx1_ASAP7_75t_L g10969 ( 
.A(n_9376),
.Y(n_10969)
);

INVx1_ASAP7_75t_L g10970 ( 
.A(n_9379),
.Y(n_10970)
);

AND2x2_ASAP7_75t_L g10971 ( 
.A(n_9221),
.B(n_8638),
.Y(n_10971)
);

NOR2xp33_ASAP7_75t_L g10972 ( 
.A(n_9310),
.B(n_8761),
.Y(n_10972)
);

INVx1_ASAP7_75t_L g10973 ( 
.A(n_9379),
.Y(n_10973)
);

BUFx2_ASAP7_75t_L g10974 ( 
.A(n_9429),
.Y(n_10974)
);

OAI21x1_ASAP7_75t_L g10975 ( 
.A1(n_9522),
.A2(n_8120),
.B(n_8106),
.Y(n_10975)
);

INVx1_ASAP7_75t_L g10976 ( 
.A(n_9382),
.Y(n_10976)
);

BUFx2_ASAP7_75t_SL g10977 ( 
.A(n_10101),
.Y(n_10977)
);

AOI22xp33_ASAP7_75t_L g10978 ( 
.A1(n_9375),
.A2(n_7808),
.B1(n_7785),
.B2(n_7843),
.Y(n_10978)
);

INVx2_ASAP7_75t_L g10979 ( 
.A(n_9743),
.Y(n_10979)
);

AOI21xp33_ASAP7_75t_L g10980 ( 
.A1(n_9528),
.A2(n_7796),
.B(n_8212),
.Y(n_10980)
);

BUFx3_ASAP7_75t_L g10981 ( 
.A(n_10102),
.Y(n_10981)
);

INVx1_ASAP7_75t_L g10982 ( 
.A(n_9382),
.Y(n_10982)
);

NAND2xp5_ASAP7_75t_SL g10983 ( 
.A(n_9941),
.B(n_8670),
.Y(n_10983)
);

O2A1O1Ixp33_ASAP7_75t_L g10984 ( 
.A1(n_9720),
.A2(n_8420),
.B(n_8825),
.C(n_8629),
.Y(n_10984)
);

BUFx3_ASAP7_75t_L g10985 ( 
.A(n_10102),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_9385),
.Y(n_10986)
);

INVx2_ASAP7_75t_L g10987 ( 
.A(n_9747),
.Y(n_10987)
);

INVx2_ASAP7_75t_L g10988 ( 
.A(n_9747),
.Y(n_10988)
);

INVx2_ASAP7_75t_L g10989 ( 
.A(n_9747),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_9385),
.Y(n_10990)
);

AND2x2_ASAP7_75t_L g10991 ( 
.A(n_9238),
.B(n_8732),
.Y(n_10991)
);

INVx2_ASAP7_75t_L g10992 ( 
.A(n_9749),
.Y(n_10992)
);

HB1xp67_ASAP7_75t_L g10993 ( 
.A(n_9596),
.Y(n_10993)
);

INVx1_ASAP7_75t_L g10994 ( 
.A(n_9397),
.Y(n_10994)
);

INVx3_ASAP7_75t_L g10995 ( 
.A(n_10048),
.Y(n_10995)
);

NAND2xp5_ASAP7_75t_L g10996 ( 
.A(n_9858),
.B(n_8667),
.Y(n_10996)
);

INVx1_ASAP7_75t_L g10997 ( 
.A(n_9397),
.Y(n_10997)
);

INVx1_ASAP7_75t_L g10998 ( 
.A(n_9404),
.Y(n_10998)
);

INVxp33_ASAP7_75t_L g10999 ( 
.A(n_9459),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_9404),
.Y(n_11000)
);

NAND2x1p5_ASAP7_75t_L g11001 ( 
.A(n_10048),
.B(n_8805),
.Y(n_11001)
);

INVx2_ASAP7_75t_L g11002 ( 
.A(n_9749),
.Y(n_11002)
);

AND2x2_ASAP7_75t_L g11003 ( 
.A(n_9238),
.B(n_8732),
.Y(n_11003)
);

AND2x2_ASAP7_75t_L g11004 ( 
.A(n_9266),
.B(n_8732),
.Y(n_11004)
);

INVx2_ASAP7_75t_L g11005 ( 
.A(n_9749),
.Y(n_11005)
);

INVx3_ASAP7_75t_L g11006 ( 
.A(n_10048),
.Y(n_11006)
);

INVx1_ASAP7_75t_L g11007 ( 
.A(n_9407),
.Y(n_11007)
);

AND2x2_ASAP7_75t_L g11008 ( 
.A(n_9266),
.B(n_8758),
.Y(n_11008)
);

INVx1_ASAP7_75t_L g11009 ( 
.A(n_9407),
.Y(n_11009)
);

AO21x2_ASAP7_75t_L g11010 ( 
.A1(n_9558),
.A2(n_8749),
.B(n_8641),
.Y(n_11010)
);

CKINVDCx5p33_ASAP7_75t_R g11011 ( 
.A(n_9463),
.Y(n_11011)
);

INVx1_ASAP7_75t_L g11012 ( 
.A(n_9408),
.Y(n_11012)
);

INVx2_ASAP7_75t_L g11013 ( 
.A(n_9756),
.Y(n_11013)
);

INVx2_ASAP7_75t_L g11014 ( 
.A(n_9756),
.Y(n_11014)
);

NAND2xp5_ASAP7_75t_L g11015 ( 
.A(n_9907),
.B(n_8667),
.Y(n_11015)
);

OR2x2_ASAP7_75t_L g11016 ( 
.A(n_9562),
.B(n_8513),
.Y(n_11016)
);

AOI22xp33_ASAP7_75t_L g11017 ( 
.A1(n_9685),
.A2(n_7808),
.B1(n_7785),
.B2(n_7843),
.Y(n_11017)
);

INVx1_ASAP7_75t_L g11018 ( 
.A(n_9408),
.Y(n_11018)
);

INVx1_ASAP7_75t_L g11019 ( 
.A(n_9414),
.Y(n_11019)
);

AO21x1_ASAP7_75t_SL g11020 ( 
.A1(n_9789),
.A2(n_8453),
.B(n_8382),
.Y(n_11020)
);

OAI21x1_ASAP7_75t_L g11021 ( 
.A1(n_9534),
.A2(n_8120),
.B(n_8106),
.Y(n_11021)
);

OR2x2_ASAP7_75t_L g11022 ( 
.A(n_9562),
.B(n_8513),
.Y(n_11022)
);

AND2x4_ASAP7_75t_L g11023 ( 
.A(n_9973),
.B(n_7905),
.Y(n_11023)
);

BUFx6f_ASAP7_75t_L g11024 ( 
.A(n_9130),
.Y(n_11024)
);

OAI21x1_ASAP7_75t_L g11025 ( 
.A1(n_9534),
.A2(n_8127),
.B(n_8120),
.Y(n_11025)
);

INVx1_ASAP7_75t_L g11026 ( 
.A(n_9414),
.Y(n_11026)
);

BUFx2_ASAP7_75t_L g11027 ( 
.A(n_9439),
.Y(n_11027)
);

AOI22xp33_ASAP7_75t_L g11028 ( 
.A1(n_9685),
.A2(n_7843),
.B1(n_8657),
.B2(n_8326),
.Y(n_11028)
);

AND2x2_ASAP7_75t_L g11029 ( 
.A(n_9289),
.B(n_8758),
.Y(n_11029)
);

INVx8_ASAP7_75t_L g11030 ( 
.A(n_9130),
.Y(n_11030)
);

OAI21x1_ASAP7_75t_L g11031 ( 
.A1(n_9541),
.A2(n_8134),
.B(n_8127),
.Y(n_11031)
);

INVx2_ASAP7_75t_L g11032 ( 
.A(n_9756),
.Y(n_11032)
);

INVx1_ASAP7_75t_L g11033 ( 
.A(n_9415),
.Y(n_11033)
);

INVx2_ASAP7_75t_L g11034 ( 
.A(n_9758),
.Y(n_11034)
);

AO21x1_ASAP7_75t_SL g11035 ( 
.A1(n_9789),
.A2(n_8663),
.B(n_8125),
.Y(n_11035)
);

BUFx6f_ASAP7_75t_L g11036 ( 
.A(n_9130),
.Y(n_11036)
);

OR2x2_ASAP7_75t_L g11037 ( 
.A(n_10377),
.B(n_8519),
.Y(n_11037)
);

AND2x2_ASAP7_75t_L g11038 ( 
.A(n_9289),
.B(n_8758),
.Y(n_11038)
);

OA21x2_ASAP7_75t_L g11039 ( 
.A1(n_10149),
.A2(n_8990),
.B(n_8985),
.Y(n_11039)
);

INVx2_ASAP7_75t_L g11040 ( 
.A(n_9758),
.Y(n_11040)
);

AND2x2_ASAP7_75t_L g11041 ( 
.A(n_10271),
.B(n_8764),
.Y(n_11041)
);

INVx2_ASAP7_75t_L g11042 ( 
.A(n_9758),
.Y(n_11042)
);

INVx2_ASAP7_75t_SL g11043 ( 
.A(n_10210),
.Y(n_11043)
);

INVx2_ASAP7_75t_L g11044 ( 
.A(n_9760),
.Y(n_11044)
);

INVx2_ASAP7_75t_L g11045 ( 
.A(n_9760),
.Y(n_11045)
);

INVx2_ASAP7_75t_L g11046 ( 
.A(n_9760),
.Y(n_11046)
);

INVx2_ASAP7_75t_L g11047 ( 
.A(n_9765),
.Y(n_11047)
);

INVx1_ASAP7_75t_L g11048 ( 
.A(n_9415),
.Y(n_11048)
);

AND2x2_ASAP7_75t_L g11049 ( 
.A(n_10271),
.B(n_8764),
.Y(n_11049)
);

INVx2_ASAP7_75t_L g11050 ( 
.A(n_9765),
.Y(n_11050)
);

INVx1_ASAP7_75t_L g11051 ( 
.A(n_9417),
.Y(n_11051)
);

INVx2_ASAP7_75t_L g11052 ( 
.A(n_9765),
.Y(n_11052)
);

INVx1_ASAP7_75t_L g11053 ( 
.A(n_9417),
.Y(n_11053)
);

INVx1_ASAP7_75t_L g11054 ( 
.A(n_9420),
.Y(n_11054)
);

INVx2_ASAP7_75t_SL g11055 ( 
.A(n_10210),
.Y(n_11055)
);

INVx2_ASAP7_75t_L g11056 ( 
.A(n_9773),
.Y(n_11056)
);

INVx1_ASAP7_75t_L g11057 ( 
.A(n_9420),
.Y(n_11057)
);

NAND2xp5_ASAP7_75t_L g11058 ( 
.A(n_9907),
.B(n_8669),
.Y(n_11058)
);

INVx2_ASAP7_75t_L g11059 ( 
.A(n_9773),
.Y(n_11059)
);

INVx1_ASAP7_75t_L g11060 ( 
.A(n_9421),
.Y(n_11060)
);

INVx3_ASAP7_75t_L g11061 ( 
.A(n_10210),
.Y(n_11061)
);

INVx3_ASAP7_75t_L g11062 ( 
.A(n_10210),
.Y(n_11062)
);

INVx1_ASAP7_75t_L g11063 ( 
.A(n_9421),
.Y(n_11063)
);

INVx2_ASAP7_75t_L g11064 ( 
.A(n_9773),
.Y(n_11064)
);

INVx1_ASAP7_75t_L g11065 ( 
.A(n_9423),
.Y(n_11065)
);

INVx1_ASAP7_75t_L g11066 ( 
.A(n_9423),
.Y(n_11066)
);

OAI22xp33_ASAP7_75t_L g11067 ( 
.A1(n_10024),
.A2(n_8777),
.B1(n_8784),
.B2(n_8772),
.Y(n_11067)
);

INVx3_ASAP7_75t_L g11068 ( 
.A(n_10210),
.Y(n_11068)
);

INVx2_ASAP7_75t_SL g11069 ( 
.A(n_10268),
.Y(n_11069)
);

OAI21x1_ASAP7_75t_L g11070 ( 
.A1(n_9541),
.A2(n_8134),
.B(n_8127),
.Y(n_11070)
);

BUFx3_ASAP7_75t_L g11071 ( 
.A(n_9288),
.Y(n_11071)
);

OAI21x1_ASAP7_75t_L g11072 ( 
.A1(n_10045),
.A2(n_10125),
.B(n_9097),
.Y(n_11072)
);

OAI211xp5_ASAP7_75t_SL g11073 ( 
.A1(n_10355),
.A2(n_8642),
.B(n_8989),
.C(n_8325),
.Y(n_11073)
);

AOI21xp5_ASAP7_75t_L g11074 ( 
.A1(n_10093),
.A2(n_7912),
.B(n_8289),
.Y(n_11074)
);

HB1xp67_ASAP7_75t_L g11075 ( 
.A(n_9616),
.Y(n_11075)
);

INVx2_ASAP7_75t_SL g11076 ( 
.A(n_10268),
.Y(n_11076)
);

AND2x2_ASAP7_75t_L g11077 ( 
.A(n_10271),
.B(n_8764),
.Y(n_11077)
);

INVx1_ASAP7_75t_L g11078 ( 
.A(n_9424),
.Y(n_11078)
);

OAI21x1_ASAP7_75t_L g11079 ( 
.A1(n_10045),
.A2(n_8134),
.B(n_8985),
.Y(n_11079)
);

NOR2x1_ASAP7_75t_SL g11080 ( 
.A(n_9518),
.B(n_8766),
.Y(n_11080)
);

NAND2xp5_ASAP7_75t_L g11081 ( 
.A(n_9383),
.B(n_8669),
.Y(n_11081)
);

OR2x2_ASAP7_75t_L g11082 ( 
.A(n_10345),
.B(n_8519),
.Y(n_11082)
);

BUFx2_ASAP7_75t_L g11083 ( 
.A(n_9439),
.Y(n_11083)
);

HB1xp67_ASAP7_75t_L g11084 ( 
.A(n_9618),
.Y(n_11084)
);

INVx1_ASAP7_75t_L g11085 ( 
.A(n_9424),
.Y(n_11085)
);

INVx1_ASAP7_75t_L g11086 ( 
.A(n_9428),
.Y(n_11086)
);

INVx2_ASAP7_75t_L g11087 ( 
.A(n_9778),
.Y(n_11087)
);

AND2x2_ASAP7_75t_L g11088 ( 
.A(n_10271),
.B(n_8862),
.Y(n_11088)
);

INVx1_ASAP7_75t_L g11089 ( 
.A(n_9428),
.Y(n_11089)
);

INVx2_ASAP7_75t_L g11090 ( 
.A(n_9778),
.Y(n_11090)
);

INVx2_ASAP7_75t_SL g11091 ( 
.A(n_10268),
.Y(n_11091)
);

OA21x2_ASAP7_75t_L g11092 ( 
.A1(n_9558),
.A2(n_9941),
.B(n_9371),
.Y(n_11092)
);

INVx2_ASAP7_75t_SL g11093 ( 
.A(n_10268),
.Y(n_11093)
);

INVx2_ASAP7_75t_L g11094 ( 
.A(n_9778),
.Y(n_11094)
);

NAND2xp5_ASAP7_75t_L g11095 ( 
.A(n_9383),
.B(n_8776),
.Y(n_11095)
);

AND2x2_ASAP7_75t_L g11096 ( 
.A(n_9066),
.B(n_8862),
.Y(n_11096)
);

NOR2x1_ASAP7_75t_L g11097 ( 
.A(n_9439),
.B(n_8761),
.Y(n_11097)
);

NAND2xp5_ASAP7_75t_L g11098 ( 
.A(n_9409),
.B(n_8776),
.Y(n_11098)
);

INVx1_ASAP7_75t_L g11099 ( 
.A(n_9433),
.Y(n_11099)
);

INVx2_ASAP7_75t_L g11100 ( 
.A(n_9780),
.Y(n_11100)
);

INVx2_ASAP7_75t_L g11101 ( 
.A(n_9780),
.Y(n_11101)
);

INVx1_ASAP7_75t_L g11102 ( 
.A(n_9433),
.Y(n_11102)
);

INVx4_ASAP7_75t_SL g11103 ( 
.A(n_9130),
.Y(n_11103)
);

INVx4_ASAP7_75t_L g11104 ( 
.A(n_9167),
.Y(n_11104)
);

INVx1_ASAP7_75t_L g11105 ( 
.A(n_9447),
.Y(n_11105)
);

OR2x2_ASAP7_75t_L g11106 ( 
.A(n_10345),
.B(n_8087),
.Y(n_11106)
);

BUFx2_ASAP7_75t_L g11107 ( 
.A(n_9288),
.Y(n_11107)
);

INVx2_ASAP7_75t_L g11108 ( 
.A(n_9780),
.Y(n_11108)
);

INVx2_ASAP7_75t_L g11109 ( 
.A(n_9782),
.Y(n_11109)
);

OAI21x1_ASAP7_75t_L g11110 ( 
.A1(n_10125),
.A2(n_8990),
.B(n_8349),
.Y(n_11110)
);

AND2x2_ASAP7_75t_L g11111 ( 
.A(n_9066),
.B(n_9132),
.Y(n_11111)
);

OAI21x1_ASAP7_75t_L g11112 ( 
.A1(n_9048),
.A2(n_8349),
.B(n_8324),
.Y(n_11112)
);

HB1xp67_ASAP7_75t_L g11113 ( 
.A(n_9629),
.Y(n_11113)
);

INVx4_ASAP7_75t_L g11114 ( 
.A(n_9167),
.Y(n_11114)
);

BUFx3_ASAP7_75t_L g11115 ( 
.A(n_9288),
.Y(n_11115)
);

AOI221xp5_ASAP7_75t_L g11116 ( 
.A1(n_10355),
.A2(n_8187),
.B1(n_8222),
.B2(n_8154),
.C(n_7967),
.Y(n_11116)
);

INVx1_ASAP7_75t_L g11117 ( 
.A(n_9447),
.Y(n_11117)
);

INVx1_ASAP7_75t_L g11118 ( 
.A(n_9456),
.Y(n_11118)
);

INVx2_ASAP7_75t_L g11119 ( 
.A(n_9782),
.Y(n_11119)
);

BUFx10_ASAP7_75t_L g11120 ( 
.A(n_9167),
.Y(n_11120)
);

INVx1_ASAP7_75t_L g11121 ( 
.A(n_9456),
.Y(n_11121)
);

NAND3xp33_ASAP7_75t_SL g11122 ( 
.A(n_9162),
.B(n_8300),
.C(n_8798),
.Y(n_11122)
);

INVx1_ASAP7_75t_L g11123 ( 
.A(n_9468),
.Y(n_11123)
);

HB1xp67_ASAP7_75t_L g11124 ( 
.A(n_9662),
.Y(n_11124)
);

INVx1_ASAP7_75t_L g11125 ( 
.A(n_9468),
.Y(n_11125)
);

INVx1_ASAP7_75t_L g11126 ( 
.A(n_9470),
.Y(n_11126)
);

INVxp67_ASAP7_75t_L g11127 ( 
.A(n_10279),
.Y(n_11127)
);

NAND2xp5_ASAP7_75t_L g11128 ( 
.A(n_9409),
.B(n_8876),
.Y(n_11128)
);

INVx1_ASAP7_75t_L g11129 ( 
.A(n_9470),
.Y(n_11129)
);

INVx2_ASAP7_75t_L g11130 ( 
.A(n_9782),
.Y(n_11130)
);

INVx2_ASAP7_75t_L g11131 ( 
.A(n_9791),
.Y(n_11131)
);

AOI221xp5_ASAP7_75t_L g11132 ( 
.A1(n_10344),
.A2(n_8187),
.B1(n_8222),
.B2(n_8154),
.C(n_7967),
.Y(n_11132)
);

INVx2_ASAP7_75t_L g11133 ( 
.A(n_9791),
.Y(n_11133)
);

INVx1_ASAP7_75t_L g11134 ( 
.A(n_9477),
.Y(n_11134)
);

OR2x6_ASAP7_75t_L g11135 ( 
.A(n_9203),
.B(n_9110),
.Y(n_11135)
);

NAND2xp5_ASAP7_75t_L g11136 ( 
.A(n_10054),
.B(n_8876),
.Y(n_11136)
);

INVx2_ASAP7_75t_L g11137 ( 
.A(n_9791),
.Y(n_11137)
);

AND2x4_ASAP7_75t_L g11138 ( 
.A(n_9973),
.B(n_7905),
.Y(n_11138)
);

INVx1_ASAP7_75t_L g11139 ( 
.A(n_9477),
.Y(n_11139)
);

AND2x2_ASAP7_75t_L g11140 ( 
.A(n_9066),
.B(n_8862),
.Y(n_11140)
);

INVx1_ASAP7_75t_L g11141 ( 
.A(n_9478),
.Y(n_11141)
);

INVx1_ASAP7_75t_L g11142 ( 
.A(n_9478),
.Y(n_11142)
);

AOI21x1_ASAP7_75t_L g11143 ( 
.A1(n_10106),
.A2(n_8222),
.B(n_8187),
.Y(n_11143)
);

INVx4_ASAP7_75t_L g11144 ( 
.A(n_9167),
.Y(n_11144)
);

INVx2_ASAP7_75t_SL g11145 ( 
.A(n_10268),
.Y(n_11145)
);

AND2x2_ASAP7_75t_L g11146 ( 
.A(n_9066),
.B(n_8895),
.Y(n_11146)
);

NAND2xp5_ASAP7_75t_L g11147 ( 
.A(n_10054),
.B(n_8893),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_9802),
.Y(n_11148)
);

INVx2_ASAP7_75t_L g11149 ( 
.A(n_9802),
.Y(n_11149)
);

HB1xp67_ASAP7_75t_L g11150 ( 
.A(n_9667),
.Y(n_11150)
);

INVx2_ASAP7_75t_L g11151 ( 
.A(n_9802),
.Y(n_11151)
);

AOI21x1_ASAP7_75t_L g11152 ( 
.A1(n_10106),
.A2(n_9347),
.B(n_9350),
.Y(n_11152)
);

HB1xp67_ASAP7_75t_L g11153 ( 
.A(n_9682),
.Y(n_11153)
);

HB1xp67_ASAP7_75t_L g11154 ( 
.A(n_9719),
.Y(n_11154)
);

INVx1_ASAP7_75t_L g11155 ( 
.A(n_9479),
.Y(n_11155)
);

OA21x2_ASAP7_75t_L g11156 ( 
.A1(n_9344),
.A2(n_7818),
.B(n_7816),
.Y(n_11156)
);

INVx3_ASAP7_75t_L g11157 ( 
.A(n_10268),
.Y(n_11157)
);

HB1xp67_ASAP7_75t_L g11158 ( 
.A(n_9763),
.Y(n_11158)
);

INVx1_ASAP7_75t_L g11159 ( 
.A(n_9479),
.Y(n_11159)
);

OAI21x1_ASAP7_75t_L g11160 ( 
.A1(n_9048),
.A2(n_8349),
.B(n_8324),
.Y(n_11160)
);

INVx2_ASAP7_75t_L g11161 ( 
.A(n_9818),
.Y(n_11161)
);

BUFx4f_ASAP7_75t_L g11162 ( 
.A(n_9167),
.Y(n_11162)
);

INVx2_ASAP7_75t_SL g11163 ( 
.A(n_10373),
.Y(n_11163)
);

INVx2_ASAP7_75t_L g11164 ( 
.A(n_9818),
.Y(n_11164)
);

HB1xp67_ASAP7_75t_L g11165 ( 
.A(n_9771),
.Y(n_11165)
);

BUFx3_ASAP7_75t_L g11166 ( 
.A(n_9288),
.Y(n_11166)
);

INVx2_ASAP7_75t_L g11167 ( 
.A(n_9818),
.Y(n_11167)
);

INVx2_ASAP7_75t_L g11168 ( 
.A(n_9821),
.Y(n_11168)
);

AOI22xp33_ASAP7_75t_L g11169 ( 
.A1(n_9643),
.A2(n_7843),
.B1(n_8657),
.B2(n_8326),
.Y(n_11169)
);

INVx1_ASAP7_75t_L g11170 ( 
.A(n_9482),
.Y(n_11170)
);

INVx2_ASAP7_75t_L g11171 ( 
.A(n_9821),
.Y(n_11171)
);

INVx1_ASAP7_75t_L g11172 ( 
.A(n_9482),
.Y(n_11172)
);

INVx1_ASAP7_75t_L g11173 ( 
.A(n_9492),
.Y(n_11173)
);

AND2x2_ASAP7_75t_L g11174 ( 
.A(n_9132),
.B(n_8895),
.Y(n_11174)
);

INVx3_ASAP7_75t_L g11175 ( 
.A(n_9564),
.Y(n_11175)
);

CKINVDCx6p67_ASAP7_75t_R g11176 ( 
.A(n_10009),
.Y(n_11176)
);

INVx1_ASAP7_75t_L g11177 ( 
.A(n_9492),
.Y(n_11177)
);

NAND2xp33_ASAP7_75t_SL g11178 ( 
.A(n_9288),
.B(n_6987),
.Y(n_11178)
);

INVx2_ASAP7_75t_SL g11179 ( 
.A(n_10373),
.Y(n_11179)
);

INVx2_ASAP7_75t_L g11180 ( 
.A(n_9821),
.Y(n_11180)
);

INVx2_ASAP7_75t_L g11181 ( 
.A(n_9824),
.Y(n_11181)
);

HB1xp67_ASAP7_75t_L g11182 ( 
.A(n_9776),
.Y(n_11182)
);

INVxp67_ASAP7_75t_L g11183 ( 
.A(n_10279),
.Y(n_11183)
);

INVx3_ASAP7_75t_L g11184 ( 
.A(n_9564),
.Y(n_11184)
);

INVx1_ASAP7_75t_L g11185 ( 
.A(n_9496),
.Y(n_11185)
);

INVx1_ASAP7_75t_L g11186 ( 
.A(n_9496),
.Y(n_11186)
);

INVx1_ASAP7_75t_L g11187 ( 
.A(n_9508),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_9824),
.Y(n_11188)
);

INVx2_ASAP7_75t_L g11189 ( 
.A(n_9824),
.Y(n_11189)
);

AND2x2_ASAP7_75t_L g11190 ( 
.A(n_9132),
.B(n_9481),
.Y(n_11190)
);

INVx1_ASAP7_75t_L g11191 ( 
.A(n_9508),
.Y(n_11191)
);

AND2x2_ASAP7_75t_L g11192 ( 
.A(n_9132),
.B(n_8895),
.Y(n_11192)
);

NAND2x1p5_ASAP7_75t_L g11193 ( 
.A(n_9128),
.B(n_8805),
.Y(n_11193)
);

INVx1_ASAP7_75t_L g11194 ( 
.A(n_9509),
.Y(n_11194)
);

HB1xp67_ASAP7_75t_L g11195 ( 
.A(n_9809),
.Y(n_11195)
);

AOI21xp5_ASAP7_75t_SL g11196 ( 
.A1(n_10252),
.A2(n_8673),
.B(n_7383),
.Y(n_11196)
);

INVx3_ASAP7_75t_L g11197 ( 
.A(n_9564),
.Y(n_11197)
);

INVx2_ASAP7_75t_L g11198 ( 
.A(n_9825),
.Y(n_11198)
);

OAI21x1_ASAP7_75t_L g11199 ( 
.A1(n_9048),
.A2(n_8350),
.B(n_8324),
.Y(n_11199)
);

INVx1_ASAP7_75t_L g11200 ( 
.A(n_9509),
.Y(n_11200)
);

INVx1_ASAP7_75t_L g11201 ( 
.A(n_9524),
.Y(n_11201)
);

AOI22xp33_ASAP7_75t_L g11202 ( 
.A1(n_9643),
.A2(n_8604),
.B1(n_8590),
.B2(n_8263),
.Y(n_11202)
);

INVx4_ASAP7_75t_L g11203 ( 
.A(n_9167),
.Y(n_11203)
);

BUFx3_ASAP7_75t_L g11204 ( 
.A(n_9387),
.Y(n_11204)
);

INVx1_ASAP7_75t_L g11205 ( 
.A(n_9524),
.Y(n_11205)
);

OR2x2_ASAP7_75t_L g11206 ( 
.A(n_9828),
.B(n_8087),
.Y(n_11206)
);

INVx1_ASAP7_75t_L g11207 ( 
.A(n_9539),
.Y(n_11207)
);

OAI21x1_ASAP7_75t_L g11208 ( 
.A1(n_9097),
.A2(n_8356),
.B(n_8350),
.Y(n_11208)
);

INVx1_ASAP7_75t_L g11209 ( 
.A(n_9539),
.Y(n_11209)
);

AND2x2_ASAP7_75t_L g11210 ( 
.A(n_9481),
.B(n_8507),
.Y(n_11210)
);

INVx2_ASAP7_75t_SL g11211 ( 
.A(n_10373),
.Y(n_11211)
);

INVx1_ASAP7_75t_L g11212 ( 
.A(n_9542),
.Y(n_11212)
);

HB1xp67_ASAP7_75t_L g11213 ( 
.A(n_9819),
.Y(n_11213)
);

AND2x2_ASAP7_75t_L g11214 ( 
.A(n_9481),
.B(n_8507),
.Y(n_11214)
);

INVx1_ASAP7_75t_L g11215 ( 
.A(n_9542),
.Y(n_11215)
);

INVx2_ASAP7_75t_L g11216 ( 
.A(n_9825),
.Y(n_11216)
);

INVx1_ASAP7_75t_L g11217 ( 
.A(n_9548),
.Y(n_11217)
);

OAI21x1_ASAP7_75t_L g11218 ( 
.A1(n_9097),
.A2(n_8356),
.B(n_8350),
.Y(n_11218)
);

INVx2_ASAP7_75t_L g11219 ( 
.A(n_9825),
.Y(n_11219)
);

INVx1_ASAP7_75t_L g11220 ( 
.A(n_9548),
.Y(n_11220)
);

BUFx3_ASAP7_75t_L g11221 ( 
.A(n_9387),
.Y(n_11221)
);

INVxp67_ASAP7_75t_L g11222 ( 
.A(n_9551),
.Y(n_11222)
);

INVx1_ASAP7_75t_L g11223 ( 
.A(n_9560),
.Y(n_11223)
);

INVx2_ASAP7_75t_L g11224 ( 
.A(n_9839),
.Y(n_11224)
);

INVx2_ASAP7_75t_L g11225 ( 
.A(n_9839),
.Y(n_11225)
);

HB1xp67_ASAP7_75t_L g11226 ( 
.A(n_9822),
.Y(n_11226)
);

OA21x2_ASAP7_75t_L g11227 ( 
.A1(n_9344),
.A2(n_7818),
.B(n_7816),
.Y(n_11227)
);

HB1xp67_ASAP7_75t_L g11228 ( 
.A(n_9859),
.Y(n_11228)
);

INVx1_ASAP7_75t_L g11229 ( 
.A(n_9560),
.Y(n_11229)
);

INVx1_ASAP7_75t_SL g11230 ( 
.A(n_9690),
.Y(n_11230)
);

INVx1_ASAP7_75t_L g11231 ( 
.A(n_9566),
.Y(n_11231)
);

AND2x2_ASAP7_75t_L g11232 ( 
.A(n_9481),
.B(n_8507),
.Y(n_11232)
);

INVx2_ASAP7_75t_L g11233 ( 
.A(n_9839),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_9566),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_9573),
.Y(n_11235)
);

INVx1_ASAP7_75t_L g11236 ( 
.A(n_9573),
.Y(n_11236)
);

INVx4_ASAP7_75t_SL g11237 ( 
.A(n_9182),
.Y(n_11237)
);

INVx1_ASAP7_75t_L g11238 ( 
.A(n_9575),
.Y(n_11238)
);

INVxp67_ASAP7_75t_L g11239 ( 
.A(n_9690),
.Y(n_11239)
);

INVx1_ASAP7_75t_L g11240 ( 
.A(n_9575),
.Y(n_11240)
);

INVxp67_ASAP7_75t_L g11241 ( 
.A(n_9406),
.Y(n_11241)
);

NAND2x1_ASAP7_75t_L g11242 ( 
.A(n_9203),
.B(n_8431),
.Y(n_11242)
);

BUFx2_ASAP7_75t_SL g11243 ( 
.A(n_10101),
.Y(n_11243)
);

OAI21x1_ASAP7_75t_L g11244 ( 
.A1(n_9196),
.A2(n_8373),
.B(n_8356),
.Y(n_11244)
);

OAI21x1_ASAP7_75t_L g11245 ( 
.A1(n_9196),
.A2(n_8379),
.B(n_8373),
.Y(n_11245)
);

BUFx3_ASAP7_75t_L g11246 ( 
.A(n_9387),
.Y(n_11246)
);

AO21x2_ASAP7_75t_L g11247 ( 
.A1(n_10180),
.A2(n_8802),
.B(n_8641),
.Y(n_11247)
);

OAI22xp5_ASAP7_75t_L g11248 ( 
.A1(n_9999),
.A2(n_8937),
.B1(n_8830),
.B2(n_8784),
.Y(n_11248)
);

AND2x2_ASAP7_75t_L g11249 ( 
.A(n_9831),
.B(n_8507),
.Y(n_11249)
);

INVx2_ASAP7_75t_L g11250 ( 
.A(n_9841),
.Y(n_11250)
);

INVx1_ASAP7_75t_L g11251 ( 
.A(n_9580),
.Y(n_11251)
);

INVx2_ASAP7_75t_L g11252 ( 
.A(n_9841),
.Y(n_11252)
);

NAND2xp5_ASAP7_75t_L g11253 ( 
.A(n_9597),
.B(n_8893),
.Y(n_11253)
);

INVx2_ASAP7_75t_L g11254 ( 
.A(n_9841),
.Y(n_11254)
);

INVxp67_ASAP7_75t_L g11255 ( 
.A(n_9406),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_9580),
.Y(n_11256)
);

INVx5_ASAP7_75t_SL g11257 ( 
.A(n_9455),
.Y(n_11257)
);

INVx3_ASAP7_75t_L g11258 ( 
.A(n_9677),
.Y(n_11258)
);

AND2x4_ASAP7_75t_L g11259 ( 
.A(n_9973),
.B(n_7941),
.Y(n_11259)
);

HB1xp67_ASAP7_75t_L g11260 ( 
.A(n_9878),
.Y(n_11260)
);

OAI21xp5_ASAP7_75t_L g11261 ( 
.A1(n_10252),
.A2(n_9533),
.B(n_9104),
.Y(n_11261)
);

BUFx3_ASAP7_75t_L g11262 ( 
.A(n_9387),
.Y(n_11262)
);

AND2x4_ASAP7_75t_L g11263 ( 
.A(n_9283),
.B(n_7941),
.Y(n_11263)
);

INVx1_ASAP7_75t_L g11264 ( 
.A(n_9583),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_9583),
.Y(n_11265)
);

INVx2_ASAP7_75t_L g11266 ( 
.A(n_9849),
.Y(n_11266)
);

OA21x2_ASAP7_75t_L g11267 ( 
.A1(n_9344),
.A2(n_7818),
.B(n_7816),
.Y(n_11267)
);

INVx2_ASAP7_75t_L g11268 ( 
.A(n_9849),
.Y(n_11268)
);

AND2x2_ASAP7_75t_L g11269 ( 
.A(n_9831),
.B(n_8507),
.Y(n_11269)
);

INVx1_ASAP7_75t_L g11270 ( 
.A(n_9588),
.Y(n_11270)
);

OR2x2_ASAP7_75t_L g11271 ( 
.A(n_9695),
.B(n_7938),
.Y(n_11271)
);

INVx3_ASAP7_75t_L g11272 ( 
.A(n_9677),
.Y(n_11272)
);

AND2x2_ASAP7_75t_L g11273 ( 
.A(n_9840),
.B(n_8507),
.Y(n_11273)
);

INVx2_ASAP7_75t_L g11274 ( 
.A(n_9849),
.Y(n_11274)
);

BUFx2_ASAP7_75t_SL g11275 ( 
.A(n_9466),
.Y(n_11275)
);

INVx3_ASAP7_75t_L g11276 ( 
.A(n_9677),
.Y(n_11276)
);

BUFx3_ASAP7_75t_L g11277 ( 
.A(n_9387),
.Y(n_11277)
);

INVx1_ASAP7_75t_L g11278 ( 
.A(n_9588),
.Y(n_11278)
);

INVx1_ASAP7_75t_L g11279 ( 
.A(n_9595),
.Y(n_11279)
);

OAI21x1_ASAP7_75t_L g11280 ( 
.A1(n_9204),
.A2(n_8379),
.B(n_8373),
.Y(n_11280)
);

INVxp67_ASAP7_75t_L g11281 ( 
.A(n_9448),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_L g11282 ( 
.A(n_9597),
.B(n_8938),
.Y(n_11282)
);

INVx1_ASAP7_75t_L g11283 ( 
.A(n_9595),
.Y(n_11283)
);

INVx2_ASAP7_75t_L g11284 ( 
.A(n_9854),
.Y(n_11284)
);

INVx2_ASAP7_75t_L g11285 ( 
.A(n_9854),
.Y(n_11285)
);

INVx2_ASAP7_75t_L g11286 ( 
.A(n_9854),
.Y(n_11286)
);

INVx1_ASAP7_75t_L g11287 ( 
.A(n_9607),
.Y(n_11287)
);

OAI22xp5_ASAP7_75t_L g11288 ( 
.A1(n_9999),
.A2(n_8937),
.B1(n_8830),
.B2(n_8663),
.Y(n_11288)
);

BUFx2_ASAP7_75t_L g11289 ( 
.A(n_9387),
.Y(n_11289)
);

NAND2xp5_ASAP7_75t_L g11290 ( 
.A(n_9684),
.B(n_8938),
.Y(n_11290)
);

INVx3_ASAP7_75t_L g11291 ( 
.A(n_9814),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_9607),
.Y(n_11292)
);

NOR2xp33_ASAP7_75t_L g11293 ( 
.A(n_9042),
.B(n_8837),
.Y(n_11293)
);

INVx2_ASAP7_75t_L g11294 ( 
.A(n_9882),
.Y(n_11294)
);

INVx2_ASAP7_75t_L g11295 ( 
.A(n_9882),
.Y(n_11295)
);

INVx1_ASAP7_75t_L g11296 ( 
.A(n_9611),
.Y(n_11296)
);

AOI21xp5_ASAP7_75t_L g11297 ( 
.A1(n_9104),
.A2(n_7912),
.B(n_8289),
.Y(n_11297)
);

INVx1_ASAP7_75t_L g11298 ( 
.A(n_9611),
.Y(n_11298)
);

INVx1_ASAP7_75t_L g11299 ( 
.A(n_9617),
.Y(n_11299)
);

INVx1_ASAP7_75t_L g11300 ( 
.A(n_9617),
.Y(n_11300)
);

AO21x2_ASAP7_75t_L g11301 ( 
.A1(n_10180),
.A2(n_8802),
.B(n_8641),
.Y(n_11301)
);

OAI21x1_ASAP7_75t_L g11302 ( 
.A1(n_9204),
.A2(n_8381),
.B(n_8379),
.Y(n_11302)
);

INVx2_ASAP7_75t_L g11303 ( 
.A(n_9882),
.Y(n_11303)
);

INVx1_ASAP7_75t_L g11304 ( 
.A(n_9626),
.Y(n_11304)
);

NAND2xp5_ASAP7_75t_L g11305 ( 
.A(n_9684),
.B(n_9091),
.Y(n_11305)
);

INVx2_ASAP7_75t_L g11306 ( 
.A(n_9883),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_9840),
.B(n_9868),
.Y(n_11307)
);

INVx1_ASAP7_75t_L g11308 ( 
.A(n_9626),
.Y(n_11308)
);

INVx2_ASAP7_75t_L g11309 ( 
.A(n_9883),
.Y(n_11309)
);

AND2x2_ASAP7_75t_L g11310 ( 
.A(n_9868),
.B(n_8287),
.Y(n_11310)
);

INVx1_ASAP7_75t_L g11311 ( 
.A(n_9632),
.Y(n_11311)
);

INVx2_ASAP7_75t_L g11312 ( 
.A(n_9883),
.Y(n_11312)
);

INVx2_ASAP7_75t_L g11313 ( 
.A(n_9892),
.Y(n_11313)
);

BUFx2_ASAP7_75t_SL g11314 ( 
.A(n_9466),
.Y(n_11314)
);

AND2x2_ASAP7_75t_L g11315 ( 
.A(n_9890),
.B(n_8287),
.Y(n_11315)
);

AO21x1_ASAP7_75t_SL g11316 ( 
.A1(n_9242),
.A2(n_9245),
.B(n_9661),
.Y(n_11316)
);

OR2x2_ASAP7_75t_L g11317 ( 
.A(n_9828),
.B(n_8087),
.Y(n_11317)
);

BUFx6f_ASAP7_75t_L g11318 ( 
.A(n_9182),
.Y(n_11318)
);

HB1xp67_ASAP7_75t_L g11319 ( 
.A(n_9889),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_9632),
.Y(n_11320)
);

NAND2x1p5_ASAP7_75t_L g11321 ( 
.A(n_9128),
.B(n_8805),
.Y(n_11321)
);

INVx2_ASAP7_75t_L g11322 ( 
.A(n_9892),
.Y(n_11322)
);

INVx2_ASAP7_75t_L g11323 ( 
.A(n_9892),
.Y(n_11323)
);

OAI21x1_ASAP7_75t_L g11324 ( 
.A1(n_9226),
.A2(n_8389),
.B(n_8381),
.Y(n_11324)
);

INVx1_ASAP7_75t_L g11325 ( 
.A(n_9638),
.Y(n_11325)
);

BUFx2_ASAP7_75t_L g11326 ( 
.A(n_9296),
.Y(n_11326)
);

INVx2_ASAP7_75t_L g11327 ( 
.A(n_9894),
.Y(n_11327)
);

OR2x6_ASAP7_75t_L g11328 ( 
.A(n_9203),
.B(n_8837),
.Y(n_11328)
);

AND2x2_ASAP7_75t_L g11329 ( 
.A(n_9890),
.B(n_8287),
.Y(n_11329)
);

INVx2_ASAP7_75t_L g11330 ( 
.A(n_9894),
.Y(n_11330)
);

INVx2_ASAP7_75t_L g11331 ( 
.A(n_9894),
.Y(n_11331)
);

INVx2_ASAP7_75t_L g11332 ( 
.A(n_9896),
.Y(n_11332)
);

INVx1_ASAP7_75t_L g11333 ( 
.A(n_9638),
.Y(n_11333)
);

AND2x2_ASAP7_75t_L g11334 ( 
.A(n_9916),
.B(n_8290),
.Y(n_11334)
);

INVx1_ASAP7_75t_L g11335 ( 
.A(n_9639),
.Y(n_11335)
);

INVx2_ASAP7_75t_SL g11336 ( 
.A(n_10373),
.Y(n_11336)
);

HB1xp67_ASAP7_75t_L g11337 ( 
.A(n_9899),
.Y(n_11337)
);

HB1xp67_ASAP7_75t_L g11338 ( 
.A(n_9900),
.Y(n_11338)
);

INVx2_ASAP7_75t_L g11339 ( 
.A(n_9896),
.Y(n_11339)
);

OAI21x1_ASAP7_75t_L g11340 ( 
.A1(n_9226),
.A2(n_8389),
.B(n_8381),
.Y(n_11340)
);

INVx1_ASAP7_75t_L g11341 ( 
.A(n_9639),
.Y(n_11341)
);

INVx2_ASAP7_75t_L g11342 ( 
.A(n_9896),
.Y(n_11342)
);

INVx1_ASAP7_75t_L g11343 ( 
.A(n_9640),
.Y(n_11343)
);

INVx1_ASAP7_75t_L g11344 ( 
.A(n_9640),
.Y(n_11344)
);

AND2x2_ASAP7_75t_L g11345 ( 
.A(n_9916),
.B(n_8290),
.Y(n_11345)
);

OAI21xp5_ASAP7_75t_L g11346 ( 
.A1(n_9744),
.A2(n_7902),
.B(n_7914),
.Y(n_11346)
);

INVx3_ASAP7_75t_L g11347 ( 
.A(n_9814),
.Y(n_11347)
);

INVx1_ASAP7_75t_L g11348 ( 
.A(n_9644),
.Y(n_11348)
);

INVx3_ASAP7_75t_L g11349 ( 
.A(n_9814),
.Y(n_11349)
);

AND2x4_ASAP7_75t_L g11350 ( 
.A(n_9283),
.B(n_7941),
.Y(n_11350)
);

AOI22xp33_ASAP7_75t_L g11351 ( 
.A1(n_10299),
.A2(n_8604),
.B1(n_8590),
.B2(n_8263),
.Y(n_11351)
);

INVx2_ASAP7_75t_L g11352 ( 
.A(n_9909),
.Y(n_11352)
);

INVx2_ASAP7_75t_L g11353 ( 
.A(n_9909),
.Y(n_11353)
);

BUFx2_ASAP7_75t_L g11354 ( 
.A(n_9296),
.Y(n_11354)
);

INVx2_ASAP7_75t_L g11355 ( 
.A(n_9909),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_9644),
.Y(n_11356)
);

INVx3_ASAP7_75t_L g11357 ( 
.A(n_9877),
.Y(n_11357)
);

CKINVDCx5p33_ASAP7_75t_R g11358 ( 
.A(n_9455),
.Y(n_11358)
);

AND2x2_ASAP7_75t_L g11359 ( 
.A(n_9917),
.B(n_8290),
.Y(n_11359)
);

INVx2_ASAP7_75t_L g11360 ( 
.A(n_9912),
.Y(n_11360)
);

AND2x2_ASAP7_75t_L g11361 ( 
.A(n_9917),
.B(n_8457),
.Y(n_11361)
);

INVx1_ASAP7_75t_L g11362 ( 
.A(n_9648),
.Y(n_11362)
);

INVx1_ASAP7_75t_L g11363 ( 
.A(n_9648),
.Y(n_11363)
);

AND2x2_ASAP7_75t_L g11364 ( 
.A(n_9934),
.B(n_8457),
.Y(n_11364)
);

OA21x2_ASAP7_75t_L g11365 ( 
.A1(n_9371),
.A2(n_8457),
.B(n_7994),
.Y(n_11365)
);

OAI22xp33_ASAP7_75t_SL g11366 ( 
.A1(n_9106),
.A2(n_8798),
.B1(n_8977),
.B2(n_8762),
.Y(n_11366)
);

INVx1_ASAP7_75t_L g11367 ( 
.A(n_9654),
.Y(n_11367)
);

HB1xp67_ASAP7_75t_L g11368 ( 
.A(n_9904),
.Y(n_11368)
);

OR2x6_ASAP7_75t_L g11369 ( 
.A(n_9203),
.B(n_8837),
.Y(n_11369)
);

AND2x2_ASAP7_75t_L g11370 ( 
.A(n_9934),
.B(n_8652),
.Y(n_11370)
);

INVx1_ASAP7_75t_L g11371 ( 
.A(n_9654),
.Y(n_11371)
);

INVx2_ASAP7_75t_L g11372 ( 
.A(n_9912),
.Y(n_11372)
);

INVx1_ASAP7_75t_L g11373 ( 
.A(n_9657),
.Y(n_11373)
);

INVx1_ASAP7_75t_L g11374 ( 
.A(n_9657),
.Y(n_11374)
);

AND2x2_ASAP7_75t_L g11375 ( 
.A(n_9956),
.B(n_8652),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_9659),
.Y(n_11376)
);

INVxp67_ASAP7_75t_L g11377 ( 
.A(n_9448),
.Y(n_11377)
);

INVx2_ASAP7_75t_L g11378 ( 
.A(n_9912),
.Y(n_11378)
);

NOR2xp33_ASAP7_75t_L g11379 ( 
.A(n_9042),
.B(n_8837),
.Y(n_11379)
);

INVx1_ASAP7_75t_L g11380 ( 
.A(n_9659),
.Y(n_11380)
);

INVx2_ASAP7_75t_L g11381 ( 
.A(n_9914),
.Y(n_11381)
);

BUFx3_ASAP7_75t_L g11382 ( 
.A(n_9131),
.Y(n_11382)
);

INVx4_ASAP7_75t_SL g11383 ( 
.A(n_9182),
.Y(n_11383)
);

INVx1_ASAP7_75t_L g11384 ( 
.A(n_9666),
.Y(n_11384)
);

OA21x2_ASAP7_75t_L g11385 ( 
.A1(n_9371),
.A2(n_7994),
.B(n_7993),
.Y(n_11385)
);

INVx1_ASAP7_75t_L g11386 ( 
.A(n_9666),
.Y(n_11386)
);

BUFx3_ASAP7_75t_L g11387 ( 
.A(n_9131),
.Y(n_11387)
);

INVx1_ASAP7_75t_L g11388 ( 
.A(n_9670),
.Y(n_11388)
);

INVx4_ASAP7_75t_L g11389 ( 
.A(n_9182),
.Y(n_11389)
);

INVx1_ASAP7_75t_L g11390 ( 
.A(n_9670),
.Y(n_11390)
);

AND2x2_ASAP7_75t_L g11391 ( 
.A(n_9956),
.B(n_8658),
.Y(n_11391)
);

AND2x2_ASAP7_75t_L g11392 ( 
.A(n_10140),
.B(n_8658),
.Y(n_11392)
);

NOR2x1p5_ASAP7_75t_L g11393 ( 
.A(n_9042),
.B(n_8837),
.Y(n_11393)
);

INVx1_ASAP7_75t_L g11394 ( 
.A(n_9673),
.Y(n_11394)
);

CKINVDCx16_ASAP7_75t_R g11395 ( 
.A(n_9619),
.Y(n_11395)
);

AND2x2_ASAP7_75t_L g11396 ( 
.A(n_10140),
.B(n_7856),
.Y(n_11396)
);

NOR2xp67_ASAP7_75t_L g11397 ( 
.A(n_9042),
.B(n_8508),
.Y(n_11397)
);

INVx1_ASAP7_75t_L g11398 ( 
.A(n_9673),
.Y(n_11398)
);

INVx2_ASAP7_75t_L g11399 ( 
.A(n_9914),
.Y(n_11399)
);

BUFx2_ASAP7_75t_L g11400 ( 
.A(n_9131),
.Y(n_11400)
);

AND2x2_ASAP7_75t_L g11401 ( 
.A(n_10175),
.B(n_7856),
.Y(n_11401)
);

BUFx2_ASAP7_75t_L g11402 ( 
.A(n_9156),
.Y(n_11402)
);

INVx2_ASAP7_75t_L g11403 ( 
.A(n_9914),
.Y(n_11403)
);

INVx1_ASAP7_75t_L g11404 ( 
.A(n_9676),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_9930),
.Y(n_11405)
);

INVx2_ASAP7_75t_L g11406 ( 
.A(n_9930),
.Y(n_11406)
);

INVx1_ASAP7_75t_L g11407 ( 
.A(n_9676),
.Y(n_11407)
);

NOR2x1_ASAP7_75t_SL g11408 ( 
.A(n_9480),
.B(n_8762),
.Y(n_11408)
);

BUFx2_ASAP7_75t_L g11409 ( 
.A(n_9156),
.Y(n_11409)
);

INVx1_ASAP7_75t_L g11410 ( 
.A(n_9687),
.Y(n_11410)
);

NAND2xp5_ASAP7_75t_L g11411 ( 
.A(n_9695),
.B(n_7958),
.Y(n_11411)
);

INVx2_ASAP7_75t_SL g11412 ( 
.A(n_9718),
.Y(n_11412)
);

INVx1_ASAP7_75t_L g11413 ( 
.A(n_9687),
.Y(n_11413)
);

INVx1_ASAP7_75t_L g11414 ( 
.A(n_9692),
.Y(n_11414)
);

INVx1_ASAP7_75t_L g11415 ( 
.A(n_9692),
.Y(n_11415)
);

OAI21x1_ASAP7_75t_L g11416 ( 
.A1(n_9877),
.A2(n_8411),
.B(n_8389),
.Y(n_11416)
);

OR2x2_ASAP7_75t_L g11417 ( 
.A(n_9784),
.B(n_9805),
.Y(n_11417)
);

INVx1_ASAP7_75t_L g11418 ( 
.A(n_9696),
.Y(n_11418)
);

INVx2_ASAP7_75t_L g11419 ( 
.A(n_9930),
.Y(n_11419)
);

HB1xp67_ASAP7_75t_L g11420 ( 
.A(n_9915),
.Y(n_11420)
);

AND2x4_ASAP7_75t_L g11421 ( 
.A(n_9395),
.B(n_7941),
.Y(n_11421)
);

OAI21x1_ASAP7_75t_L g11422 ( 
.A1(n_9877),
.A2(n_8419),
.B(n_8411),
.Y(n_11422)
);

INVx3_ASAP7_75t_L g11423 ( 
.A(n_9951),
.Y(n_11423)
);

INVx2_ASAP7_75t_L g11424 ( 
.A(n_9932),
.Y(n_11424)
);

INVx2_ASAP7_75t_L g11425 ( 
.A(n_9932),
.Y(n_11425)
);

HB1xp67_ASAP7_75t_L g11426 ( 
.A(n_9992),
.Y(n_11426)
);

INVx1_ASAP7_75t_L g11427 ( 
.A(n_9696),
.Y(n_11427)
);

INVx1_ASAP7_75t_L g11428 ( 
.A(n_9701),
.Y(n_11428)
);

INVx2_ASAP7_75t_L g11429 ( 
.A(n_9932),
.Y(n_11429)
);

INVx1_ASAP7_75t_L g11430 ( 
.A(n_9701),
.Y(n_11430)
);

INVx1_ASAP7_75t_L g11431 ( 
.A(n_9705),
.Y(n_11431)
);

AND2x2_ASAP7_75t_L g11432 ( 
.A(n_10175),
.B(n_7856),
.Y(n_11432)
);

OR2x2_ASAP7_75t_L g11433 ( 
.A(n_9784),
.B(n_7938),
.Y(n_11433)
);

BUFx6f_ASAP7_75t_L g11434 ( 
.A(n_9182),
.Y(n_11434)
);

BUFx2_ASAP7_75t_L g11435 ( 
.A(n_9156),
.Y(n_11435)
);

AND2x2_ASAP7_75t_L g11436 ( 
.A(n_10224),
.B(n_7859),
.Y(n_11436)
);

BUFx2_ASAP7_75t_SL g11437 ( 
.A(n_9161),
.Y(n_11437)
);

INVx2_ASAP7_75t_L g11438 ( 
.A(n_9939),
.Y(n_11438)
);

INVx2_ASAP7_75t_L g11439 ( 
.A(n_9939),
.Y(n_11439)
);

INVx1_ASAP7_75t_L g11440 ( 
.A(n_9705),
.Y(n_11440)
);

INVx2_ASAP7_75t_L g11441 ( 
.A(n_9939),
.Y(n_11441)
);

HB1xp67_ASAP7_75t_L g11442 ( 
.A(n_9993),
.Y(n_11442)
);

CKINVDCx14_ASAP7_75t_R g11443 ( 
.A(n_9037),
.Y(n_11443)
);

BUFx2_ASAP7_75t_L g11444 ( 
.A(n_9328),
.Y(n_11444)
);

INVx2_ASAP7_75t_L g11445 ( 
.A(n_9940),
.Y(n_11445)
);

BUFx4f_ASAP7_75t_SL g11446 ( 
.A(n_9182),
.Y(n_11446)
);

AOI22xp33_ASAP7_75t_L g11447 ( 
.A1(n_10299),
.A2(n_8604),
.B1(n_8590),
.B2(n_8275),
.Y(n_11447)
);

NOR4xp25_ASAP7_75t_SL g11448 ( 
.A(n_9117),
.B(n_8420),
.C(n_7773),
.D(n_8427),
.Y(n_11448)
);

INVx1_ASAP7_75t_L g11449 ( 
.A(n_9710),
.Y(n_11449)
);

INVx1_ASAP7_75t_L g11450 ( 
.A(n_9710),
.Y(n_11450)
);

AOI21xp33_ASAP7_75t_L g11451 ( 
.A1(n_9585),
.A2(n_8212),
.B(n_8458),
.Y(n_11451)
);

INVx1_ASAP7_75t_L g11452 ( 
.A(n_9715),
.Y(n_11452)
);

CKINVDCx5p33_ASAP7_75t_R g11453 ( 
.A(n_10112),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_9715),
.Y(n_11454)
);

INVx1_ASAP7_75t_L g11455 ( 
.A(n_9716),
.Y(n_11455)
);

CKINVDCx5p33_ASAP7_75t_R g11456 ( 
.A(n_10112),
.Y(n_11456)
);

NAND2x1p5_ASAP7_75t_L g11457 ( 
.A(n_9255),
.B(n_8953),
.Y(n_11457)
);

INVx2_ASAP7_75t_L g11458 ( 
.A(n_9940),
.Y(n_11458)
);

INVx1_ASAP7_75t_L g11459 ( 
.A(n_9716),
.Y(n_11459)
);

INVx3_ASAP7_75t_L g11460 ( 
.A(n_9951),
.Y(n_11460)
);

AND2x2_ASAP7_75t_L g11461 ( 
.A(n_10224),
.B(n_7859),
.Y(n_11461)
);

INVx1_ASAP7_75t_L g11462 ( 
.A(n_9721),
.Y(n_11462)
);

AND2x2_ASAP7_75t_L g11463 ( 
.A(n_10253),
.B(n_7859),
.Y(n_11463)
);

INVx3_ASAP7_75t_L g11464 ( 
.A(n_9951),
.Y(n_11464)
);

NAND2xp5_ASAP7_75t_L g11465 ( 
.A(n_9805),
.B(n_7958),
.Y(n_11465)
);

BUFx2_ASAP7_75t_L g11466 ( 
.A(n_9561),
.Y(n_11466)
);

OAI21x1_ASAP7_75t_L g11467 ( 
.A1(n_9962),
.A2(n_8419),
.B(n_8411),
.Y(n_11467)
);

NAND2xp5_ASAP7_75t_L g11468 ( 
.A(n_10376),
.B(n_8927),
.Y(n_11468)
);

INVx2_ASAP7_75t_L g11469 ( 
.A(n_9940),
.Y(n_11469)
);

INVx1_ASAP7_75t_L g11470 ( 
.A(n_9721),
.Y(n_11470)
);

INVx2_ASAP7_75t_L g11471 ( 
.A(n_9942),
.Y(n_11471)
);

NAND2xp5_ASAP7_75t_L g11472 ( 
.A(n_10376),
.B(n_8927),
.Y(n_11472)
);

HB1xp67_ASAP7_75t_L g11473 ( 
.A(n_9255),
.Y(n_11473)
);

INVx2_ASAP7_75t_L g11474 ( 
.A(n_9942),
.Y(n_11474)
);

OR2x2_ASAP7_75t_L g11475 ( 
.A(n_9830),
.B(n_8087),
.Y(n_11475)
);

OR2x2_ASAP7_75t_L g11476 ( 
.A(n_9830),
.B(n_8087),
.Y(n_11476)
);

INVx2_ASAP7_75t_L g11477 ( 
.A(n_9942),
.Y(n_11477)
);

NAND2xp5_ASAP7_75t_L g11478 ( 
.A(n_9898),
.B(n_8958),
.Y(n_11478)
);

BUFx6f_ASAP7_75t_L g11479 ( 
.A(n_9212),
.Y(n_11479)
);

INVx1_ASAP7_75t_SL g11480 ( 
.A(n_9486),
.Y(n_11480)
);

INVx1_ASAP7_75t_L g11481 ( 
.A(n_9722),
.Y(n_11481)
);

INVx1_ASAP7_75t_L g11482 ( 
.A(n_9722),
.Y(n_11482)
);

NAND2xp5_ASAP7_75t_L g11483 ( 
.A(n_9898),
.B(n_8958),
.Y(n_11483)
);

BUFx10_ASAP7_75t_L g11484 ( 
.A(n_9212),
.Y(n_11484)
);

INVx2_ASAP7_75t_L g11485 ( 
.A(n_9944),
.Y(n_11485)
);

INVx1_ASAP7_75t_L g11486 ( 
.A(n_9726),
.Y(n_11486)
);

INVx1_ASAP7_75t_L g11487 ( 
.A(n_9726),
.Y(n_11487)
);

INVxp67_ASAP7_75t_L g11488 ( 
.A(n_9486),
.Y(n_11488)
);

INVx1_ASAP7_75t_L g11489 ( 
.A(n_9732),
.Y(n_11489)
);

AND2x2_ASAP7_75t_L g11490 ( 
.A(n_10253),
.B(n_8959),
.Y(n_11490)
);

INVx1_ASAP7_75t_L g11491 ( 
.A(n_9732),
.Y(n_11491)
);

INVx1_ASAP7_75t_L g11492 ( 
.A(n_9737),
.Y(n_11492)
);

INVx1_ASAP7_75t_L g11493 ( 
.A(n_9737),
.Y(n_11493)
);

OAI21x1_ASAP7_75t_L g11494 ( 
.A1(n_9962),
.A2(n_8422),
.B(n_8419),
.Y(n_11494)
);

AOI222xp33_ASAP7_75t_L g11495 ( 
.A1(n_9585),
.A2(n_9020),
.B1(n_8984),
.B2(n_8980),
.C1(n_8407),
.C2(n_8699),
.Y(n_11495)
);

INVx1_ASAP7_75t_L g11496 ( 
.A(n_9738),
.Y(n_11496)
);

BUFx3_ASAP7_75t_L g11497 ( 
.A(n_9105),
.Y(n_11497)
);

INVx2_ASAP7_75t_L g11498 ( 
.A(n_9944),
.Y(n_11498)
);

INVx1_ASAP7_75t_L g11499 ( 
.A(n_9738),
.Y(n_11499)
);

NAND2xp5_ASAP7_75t_L g11500 ( 
.A(n_9092),
.B(n_8202),
.Y(n_11500)
);

INVx1_ASAP7_75t_L g11501 ( 
.A(n_9740),
.Y(n_11501)
);

INVx1_ASAP7_75t_L g11502 ( 
.A(n_9740),
.Y(n_11502)
);

BUFx2_ASAP7_75t_L g11503 ( 
.A(n_9046),
.Y(n_11503)
);

NAND2xp5_ASAP7_75t_L g11504 ( 
.A(n_9968),
.B(n_8202),
.Y(n_11504)
);

OA21x2_ASAP7_75t_L g11505 ( 
.A1(n_9398),
.A2(n_7994),
.B(n_7993),
.Y(n_11505)
);

INVx1_ASAP7_75t_L g11506 ( 
.A(n_9746),
.Y(n_11506)
);

OAI21x1_ASAP7_75t_L g11507 ( 
.A1(n_9962),
.A2(n_8425),
.B(n_8422),
.Y(n_11507)
);

INVx2_ASAP7_75t_L g11508 ( 
.A(n_9944),
.Y(n_11508)
);

OR2x2_ASAP7_75t_L g11509 ( 
.A(n_9416),
.B(n_8087),
.Y(n_11509)
);

INVx2_ASAP7_75t_L g11510 ( 
.A(n_9953),
.Y(n_11510)
);

BUFx3_ASAP7_75t_L g11511 ( 
.A(n_9105),
.Y(n_11511)
);

INVx1_ASAP7_75t_L g11512 ( 
.A(n_9746),
.Y(n_11512)
);

INVx1_ASAP7_75t_L g11513 ( 
.A(n_9762),
.Y(n_11513)
);

INVx2_ASAP7_75t_SL g11514 ( 
.A(n_9718),
.Y(n_11514)
);

INVx2_ASAP7_75t_L g11515 ( 
.A(n_9953),
.Y(n_11515)
);

BUFx2_ASAP7_75t_L g11516 ( 
.A(n_9046),
.Y(n_11516)
);

INVx1_ASAP7_75t_L g11517 ( 
.A(n_9762),
.Y(n_11517)
);

NAND2x1p5_ASAP7_75t_L g11518 ( 
.A(n_9446),
.B(n_8953),
.Y(n_11518)
);

HB1xp67_ASAP7_75t_L g11519 ( 
.A(n_9446),
.Y(n_11519)
);

INVx1_ASAP7_75t_L g11520 ( 
.A(n_9772),
.Y(n_11520)
);

AOI21xp5_ASAP7_75t_L g11521 ( 
.A1(n_9115),
.A2(n_8035),
.B(n_8163),
.Y(n_11521)
);

CKINVDCx5p33_ASAP7_75t_R g11522 ( 
.A(n_9586),
.Y(n_11522)
);

INVx1_ASAP7_75t_L g11523 ( 
.A(n_9772),
.Y(n_11523)
);

INVx2_ASAP7_75t_L g11524 ( 
.A(n_9953),
.Y(n_11524)
);

INVx1_ASAP7_75t_L g11525 ( 
.A(n_9775),
.Y(n_11525)
);

OAI21x1_ASAP7_75t_L g11526 ( 
.A1(n_10233),
.A2(n_8425),
.B(n_8422),
.Y(n_11526)
);

AOI22xp5_ASAP7_75t_L g11527 ( 
.A1(n_9795),
.A2(n_8192),
.B1(n_8576),
.B2(n_8505),
.Y(n_11527)
);

AOI21x1_ASAP7_75t_L g11528 ( 
.A1(n_9347),
.A2(n_8001),
.B(n_7951),
.Y(n_11528)
);

OR2x2_ASAP7_75t_L g11529 ( 
.A(n_9416),
.B(n_8087),
.Y(n_11529)
);

INVx2_ASAP7_75t_L g11530 ( 
.A(n_9964),
.Y(n_11530)
);

BUFx3_ASAP7_75t_L g11531 ( 
.A(n_9105),
.Y(n_11531)
);

BUFx2_ASAP7_75t_L g11532 ( 
.A(n_9046),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_9775),
.Y(n_11533)
);

HB1xp67_ASAP7_75t_L g11534 ( 
.A(n_9493),
.Y(n_11534)
);

OR2x6_ASAP7_75t_L g11535 ( 
.A(n_9203),
.B(n_7766),
.Y(n_11535)
);

OAI21x1_ASAP7_75t_L g11536 ( 
.A1(n_10233),
.A2(n_8456),
.B(n_8425),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_9783),
.Y(n_11537)
);

INVx3_ASAP7_75t_L g11538 ( 
.A(n_10233),
.Y(n_11538)
);

INVx2_ASAP7_75t_SL g11539 ( 
.A(n_9718),
.Y(n_11539)
);

INVxp67_ASAP7_75t_L g11540 ( 
.A(n_9502),
.Y(n_11540)
);

INVx2_ASAP7_75t_L g11541 ( 
.A(n_9964),
.Y(n_11541)
);

HB1xp67_ASAP7_75t_L g11542 ( 
.A(n_11473),
.Y(n_11542)
);

AOI22xp33_ASAP7_75t_L g11543 ( 
.A1(n_10433),
.A2(n_9162),
.B1(n_9893),
.B2(n_9115),
.Y(n_11543)
);

INVx1_ASAP7_75t_L g11544 ( 
.A(n_10391),
.Y(n_11544)
);

INVx2_ASAP7_75t_L g11545 ( 
.A(n_11071),
.Y(n_11545)
);

NAND2xp5_ASAP7_75t_L g11546 ( 
.A(n_10555),
.B(n_9619),
.Y(n_11546)
);

OAI21xp33_ASAP7_75t_L g11547 ( 
.A1(n_10856),
.A2(n_10240),
.B(n_10304),
.Y(n_11547)
);

OAI22xp33_ASAP7_75t_SL g11548 ( 
.A1(n_10856),
.A2(n_9106),
.B1(n_10078),
.B2(n_10131),
.Y(n_11548)
);

INVx1_ASAP7_75t_L g11549 ( 
.A(n_10397),
.Y(n_11549)
);

AOI22xp33_ASAP7_75t_L g11550 ( 
.A1(n_10855),
.A2(n_9403),
.B1(n_9945),
.B2(n_9035),
.Y(n_11550)
);

NAND2xp5_ASAP7_75t_L g11551 ( 
.A(n_10555),
.B(n_9459),
.Y(n_11551)
);

AND2x2_ASAP7_75t_L g11552 ( 
.A(n_11395),
.B(n_9935),
.Y(n_11552)
);

INVx1_ASAP7_75t_L g11553 ( 
.A(n_10432),
.Y(n_11553)
);

BUFx6f_ASAP7_75t_L g11554 ( 
.A(n_10422),
.Y(n_11554)
);

AOI22xp33_ASAP7_75t_L g11555 ( 
.A1(n_10855),
.A2(n_9403),
.B1(n_9035),
.B2(n_9229),
.Y(n_11555)
);

AOI22xp33_ASAP7_75t_L g11556 ( 
.A1(n_10855),
.A2(n_9229),
.B1(n_9186),
.B2(n_10078),
.Y(n_11556)
);

OAI221xp5_ASAP7_75t_L g11557 ( 
.A1(n_10528),
.A2(n_10240),
.B1(n_9106),
.B2(n_9544),
.C(n_10078),
.Y(n_11557)
);

AOI22xp33_ASAP7_75t_SL g11558 ( 
.A1(n_11261),
.A2(n_9235),
.B1(n_9460),
.B2(n_10289),
.Y(n_11558)
);

BUFx2_ASAP7_75t_L g11559 ( 
.A(n_11326),
.Y(n_11559)
);

AOI22xp33_ASAP7_75t_SL g11560 ( 
.A1(n_10436),
.A2(n_9235),
.B1(n_9460),
.B2(n_10289),
.Y(n_11560)
);

OAI211xp5_ASAP7_75t_SL g11561 ( 
.A1(n_10480),
.A2(n_10368),
.B(n_9432),
.C(n_10181),
.Y(n_11561)
);

NAND3xp33_ASAP7_75t_L g11562 ( 
.A(n_10467),
.B(n_10273),
.C(n_9186),
.Y(n_11562)
);

AOI22xp33_ASAP7_75t_SL g11563 ( 
.A1(n_10538),
.A2(n_10352),
.B1(n_9360),
.B2(n_10131),
.Y(n_11563)
);

OAI211xp5_ASAP7_75t_L g11564 ( 
.A1(n_10708),
.A2(n_10181),
.B(n_9252),
.C(n_10209),
.Y(n_11564)
);

INVx2_ASAP7_75t_L g11565 ( 
.A(n_11071),
.Y(n_11565)
);

AOI21xp5_ASAP7_75t_L g11566 ( 
.A1(n_11074),
.A2(n_10352),
.B(n_10086),
.Y(n_11566)
);

NAND2xp5_ASAP7_75t_L g11567 ( 
.A(n_10387),
.B(n_9968),
.Y(n_11567)
);

OR2x2_ASAP7_75t_SL g11568 ( 
.A(n_10734),
.B(n_9212),
.Y(n_11568)
);

INVx5_ASAP7_75t_L g11569 ( 
.A(n_10632),
.Y(n_11569)
);

BUFx6f_ASAP7_75t_L g11570 ( 
.A(n_10422),
.Y(n_11570)
);

OAI211xp5_ASAP7_75t_L g11571 ( 
.A1(n_11122),
.A2(n_9252),
.B(n_9794),
.C(n_9652),
.Y(n_11571)
);

INVx1_ASAP7_75t_L g11572 ( 
.A(n_10455),
.Y(n_11572)
);

INVx1_ASAP7_75t_L g11573 ( 
.A(n_10456),
.Y(n_11573)
);

AOI22xp33_ASAP7_75t_L g11574 ( 
.A1(n_11451),
.A2(n_9480),
.B1(n_9489),
.B2(n_10038),
.Y(n_11574)
);

OAI221xp5_ASAP7_75t_L g11575 ( 
.A1(n_11028),
.A2(n_9485),
.B1(n_10364),
.B2(n_10086),
.C(n_9234),
.Y(n_11575)
);

AOI211xp5_ASAP7_75t_L g11576 ( 
.A1(n_10999),
.A2(n_9735),
.B(n_9231),
.C(n_10067),
.Y(n_11576)
);

OAI22xp33_ASAP7_75t_L g11577 ( 
.A1(n_10870),
.A2(n_9500),
.B1(n_9652),
.B2(n_9360),
.Y(n_11577)
);

AOI22xp33_ASAP7_75t_L g11578 ( 
.A1(n_11495),
.A2(n_9489),
.B1(n_10038),
.B2(n_9231),
.Y(n_11578)
);

AND2x2_ASAP7_75t_L g11579 ( 
.A(n_10470),
.B(n_10325),
.Y(n_11579)
);

AND2x2_ASAP7_75t_L g11580 ( 
.A(n_10470),
.B(n_9395),
.Y(n_11580)
);

BUFx6f_ASAP7_75t_L g11581 ( 
.A(n_10632),
.Y(n_11581)
);

AOI21xp5_ASAP7_75t_L g11582 ( 
.A1(n_11521),
.A2(n_9523),
.B(n_10067),
.Y(n_11582)
);

AOI221xp5_ASAP7_75t_L g11583 ( 
.A1(n_10467),
.A2(n_9795),
.B1(n_9807),
.B2(n_9579),
.C(n_9803),
.Y(n_11583)
);

AOI22xp33_ASAP7_75t_L g11584 ( 
.A1(n_10418),
.A2(n_9261),
.B1(n_9735),
.B2(n_9279),
.Y(n_11584)
);

AOI22xp33_ASAP7_75t_L g11585 ( 
.A1(n_11028),
.A2(n_9261),
.B1(n_9279),
.B2(n_9206),
.Y(n_11585)
);

OAI22xp33_ASAP7_75t_L g11586 ( 
.A1(n_10833),
.A2(n_9500),
.B1(n_9661),
.B2(n_9794),
.Y(n_11586)
);

OAI221xp5_ASAP7_75t_L g11587 ( 
.A1(n_11169),
.A2(n_9402),
.B1(n_9578),
.B2(n_10360),
.C(n_10301),
.Y(n_11587)
);

AOI22xp33_ASAP7_75t_L g11588 ( 
.A1(n_11169),
.A2(n_9206),
.B1(n_9750),
.B2(n_9056),
.Y(n_11588)
);

AOI22xp33_ASAP7_75t_SL g11589 ( 
.A1(n_11408),
.A2(n_9750),
.B1(n_9987),
.B2(n_9954),
.Y(n_11589)
);

AOI22xp33_ASAP7_75t_L g11590 ( 
.A1(n_11035),
.A2(n_9199),
.B1(n_9193),
.B2(n_9987),
.Y(n_11590)
);

AOI22xp33_ASAP7_75t_L g11591 ( 
.A1(n_11248),
.A2(n_9647),
.B1(n_9062),
.B2(n_9954),
.Y(n_11591)
);

AOI22xp33_ASAP7_75t_L g11592 ( 
.A1(n_11067),
.A2(n_9647),
.B1(n_9364),
.B2(n_9032),
.Y(n_11592)
);

NOR3xp33_ASAP7_75t_L g11593 ( 
.A(n_11152),
.B(n_9055),
.C(n_9046),
.Y(n_11593)
);

OAI22xp5_ASAP7_75t_L g11594 ( 
.A1(n_10586),
.A2(n_9051),
.B1(n_9073),
.B2(n_10165),
.Y(n_11594)
);

AOI22xp33_ASAP7_75t_L g11595 ( 
.A1(n_11316),
.A2(n_9103),
.B1(n_9137),
.B2(n_9077),
.Y(n_11595)
);

AOI222xp33_ASAP7_75t_L g11596 ( 
.A1(n_11136),
.A2(n_9807),
.B1(n_9700),
.B2(n_9668),
.C1(n_9997),
.C2(n_10033),
.Y(n_11596)
);

AOI22xp5_ASAP7_75t_L g11597 ( 
.A1(n_10930),
.A2(n_10316),
.B1(n_9700),
.B2(n_9937),
.Y(n_11597)
);

INVx1_ASAP7_75t_L g11598 ( 
.A(n_10521),
.Y(n_11598)
);

AOI22xp33_ASAP7_75t_L g11599 ( 
.A1(n_11288),
.A2(n_9668),
.B1(n_9308),
.B2(n_9837),
.Y(n_11599)
);

AOI22xp33_ASAP7_75t_L g11600 ( 
.A1(n_10983),
.A2(n_9149),
.B1(n_9997),
.B2(n_9265),
.Y(n_11600)
);

OR2x2_ASAP7_75t_L g11601 ( 
.A(n_10415),
.B(n_10076),
.Y(n_11601)
);

BUFx2_ASAP7_75t_L g11602 ( 
.A(n_11354),
.Y(n_11602)
);

AND2x2_ASAP7_75t_L g11603 ( 
.A(n_11444),
.B(n_9396),
.Y(n_11603)
);

OAI22xp33_ASAP7_75t_L g11604 ( 
.A1(n_10999),
.A2(n_9453),
.B1(n_9329),
.B2(n_10339),
.Y(n_11604)
);

AOI22xp33_ASAP7_75t_L g11605 ( 
.A1(n_10983),
.A2(n_10033),
.B1(n_9307),
.B2(n_9381),
.Y(n_11605)
);

OAI21xp33_ASAP7_75t_L g11606 ( 
.A1(n_10523),
.A2(n_11202),
.B(n_10675),
.Y(n_11606)
);

NAND2xp5_ASAP7_75t_L g11607 ( 
.A(n_10387),
.B(n_9978),
.Y(n_11607)
);

AOI221xp5_ASAP7_75t_L g11608 ( 
.A1(n_11202),
.A2(n_10008),
.B1(n_9117),
.B2(n_9232),
.C(n_9159),
.Y(n_11608)
);

AOI22xp33_ASAP7_75t_L g11609 ( 
.A1(n_10813),
.A2(n_9267),
.B1(n_9326),
.B2(n_10176),
.Y(n_11609)
);

AOI21xp5_ASAP7_75t_L g11610 ( 
.A1(n_11297),
.A2(n_10586),
.B(n_11147),
.Y(n_11610)
);

AOI22xp33_ASAP7_75t_L g11611 ( 
.A1(n_11073),
.A2(n_9258),
.B1(n_9733),
.B2(n_9431),
.Y(n_11611)
);

NAND2xp5_ASAP7_75t_SL g11612 ( 
.A(n_11366),
.B(n_9490),
.Y(n_11612)
);

AOI22xp33_ASAP7_75t_L g11613 ( 
.A1(n_10641),
.A2(n_9450),
.B1(n_9538),
.B2(n_9761),
.Y(n_11613)
);

AOI33xp33_ASAP7_75t_L g11614 ( 
.A1(n_10948),
.A2(n_9510),
.A3(n_9507),
.B1(n_10272),
.B2(n_10288),
.B3(n_9513),
.Y(n_11614)
);

AOI21xp5_ASAP7_75t_L g11615 ( 
.A1(n_10984),
.A2(n_9523),
.B(n_9241),
.Y(n_11615)
);

INVx1_ASAP7_75t_L g11616 ( 
.A(n_10546),
.Y(n_11616)
);

OAI22xp5_ASAP7_75t_L g11617 ( 
.A1(n_10641),
.A2(n_10177),
.B1(n_10219),
.B2(n_10165),
.Y(n_11617)
);

INVx2_ASAP7_75t_SL g11618 ( 
.A(n_10632),
.Y(n_11618)
);

AOI211xp5_ASAP7_75t_L g11619 ( 
.A1(n_10980),
.A2(n_10206),
.B(n_9453),
.C(n_10050),
.Y(n_11619)
);

AO21x2_ASAP7_75t_L g11620 ( 
.A1(n_10478),
.A2(n_9350),
.B(n_9370),
.Y(n_11620)
);

INVx2_ASAP7_75t_L g11621 ( 
.A(n_11115),
.Y(n_11621)
);

OAI221xp5_ASAP7_75t_L g11622 ( 
.A1(n_10523),
.A2(n_10644),
.B1(n_10675),
.B2(n_10624),
.C(n_10642),
.Y(n_11622)
);

OAI22xp5_ASAP7_75t_L g11623 ( 
.A1(n_11351),
.A2(n_10219),
.B1(n_10177),
.B2(n_9790),
.Y(n_11623)
);

INVx2_ASAP7_75t_L g11624 ( 
.A(n_11115),
.Y(n_11624)
);

AND2x4_ASAP7_75t_L g11625 ( 
.A(n_11097),
.B(n_9114),
.Y(n_11625)
);

OR2x2_ASAP7_75t_L g11626 ( 
.A(n_10839),
.B(n_10076),
.Y(n_11626)
);

AOI22xp33_ASAP7_75t_L g11627 ( 
.A1(n_10617),
.A2(n_9538),
.B1(n_9769),
.B2(n_9334),
.Y(n_11627)
);

AOI221xp5_ASAP7_75t_L g11628 ( 
.A1(n_10948),
.A2(n_9145),
.B1(n_9273),
.B2(n_9232),
.C(n_9159),
.Y(n_11628)
);

INVx1_ASAP7_75t_L g11629 ( 
.A(n_10608),
.Y(n_11629)
);

AOI221xp5_ASAP7_75t_L g11630 ( 
.A1(n_10978),
.A2(n_9145),
.B1(n_9342),
.B2(n_9273),
.C(n_9241),
.Y(n_11630)
);

INVx2_ASAP7_75t_L g11631 ( 
.A(n_11166),
.Y(n_11631)
);

AOI22xp33_ASAP7_75t_L g11632 ( 
.A1(n_11020),
.A2(n_9823),
.B1(n_9869),
.B2(n_9329),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_10616),
.Y(n_11633)
);

AOI22xp33_ASAP7_75t_SL g11634 ( 
.A1(n_10781),
.A2(n_9342),
.B1(n_9770),
.B2(n_7815),
.Y(n_11634)
);

OAI22xp5_ASAP7_75t_L g11635 ( 
.A1(n_11351),
.A2(n_9790),
.B1(n_9977),
.B2(n_9262),
.Y(n_11635)
);

OAI22xp33_ASAP7_75t_L g11636 ( 
.A1(n_11527),
.A2(n_9488),
.B1(n_9567),
.B2(n_9454),
.Y(n_11636)
);

AOI22xp33_ASAP7_75t_L g11637 ( 
.A1(n_11466),
.A2(n_10649),
.B1(n_11500),
.B2(n_10598),
.Y(n_11637)
);

AOI22xp33_ASAP7_75t_SL g11638 ( 
.A1(n_10757),
.A2(n_9770),
.B1(n_7815),
.B2(n_10295),
.Y(n_11638)
);

AOI22xp33_ASAP7_75t_L g11639 ( 
.A1(n_11305),
.A2(n_9369),
.B1(n_9457),
.B2(n_9918),
.Y(n_11639)
);

AOI22xp33_ASAP7_75t_L g11640 ( 
.A1(n_11176),
.A2(n_9127),
.B1(n_9834),
.B2(n_9584),
.Y(n_11640)
);

INVx1_ASAP7_75t_L g11641 ( 
.A(n_10658),
.Y(n_11641)
);

AOI22xp33_ASAP7_75t_L g11642 ( 
.A1(n_11176),
.A2(n_9410),
.B1(n_9672),
.B2(n_9584),
.Y(n_11642)
);

AOI21xp5_ASAP7_75t_SL g11643 ( 
.A1(n_10567),
.A2(n_10043),
.B(n_9080),
.Y(n_11643)
);

AOI22xp33_ASAP7_75t_L g11644 ( 
.A1(n_10575),
.A2(n_9410),
.B1(n_9672),
.B2(n_9584),
.Y(n_11644)
);

AOI22xp33_ASAP7_75t_L g11645 ( 
.A1(n_11132),
.A2(n_11483),
.B1(n_11478),
.B2(n_10670),
.Y(n_11645)
);

AOI221xp5_ASAP7_75t_L g11646 ( 
.A1(n_10978),
.A2(n_9748),
.B1(n_9332),
.B2(n_9337),
.C(n_9546),
.Y(n_11646)
);

OAI22xp5_ASAP7_75t_L g11647 ( 
.A1(n_11447),
.A2(n_9977),
.B1(n_9118),
.B2(n_9563),
.Y(n_11647)
);

AOI22xp33_ASAP7_75t_L g11648 ( 
.A1(n_10905),
.A2(n_9410),
.B1(n_9672),
.B2(n_9584),
.Y(n_11648)
);

INVx2_ASAP7_75t_SL g11649 ( 
.A(n_10632),
.Y(n_11649)
);

AND2x2_ASAP7_75t_L g11650 ( 
.A(n_11111),
.B(n_9396),
.Y(n_11650)
);

AND2x2_ASAP7_75t_SL g11651 ( 
.A(n_10940),
.B(n_9055),
.Y(n_11651)
);

AND2x2_ASAP7_75t_L g11652 ( 
.A(n_11111),
.B(n_9516),
.Y(n_11652)
);

AOI22xp5_ASAP7_75t_L g11653 ( 
.A1(n_10520),
.A2(n_10375),
.B1(n_9759),
.B2(n_9569),
.Y(n_11653)
);

AOI22xp33_ASAP7_75t_L g11654 ( 
.A1(n_11468),
.A2(n_9410),
.B1(n_9672),
.B2(n_9584),
.Y(n_11654)
);

OAI22xp33_ASAP7_75t_L g11655 ( 
.A1(n_10926),
.A2(n_9567),
.B1(n_9702),
.B2(n_9488),
.Y(n_11655)
);

INVx2_ASAP7_75t_L g11656 ( 
.A(n_11166),
.Y(n_11656)
);

OAI22xp5_ASAP7_75t_L g11657 ( 
.A1(n_11447),
.A2(n_9356),
.B1(n_9645),
.B2(n_9599),
.Y(n_11657)
);

AND2x2_ASAP7_75t_L g11658 ( 
.A(n_11190),
.B(n_9516),
.Y(n_11658)
);

NAND2xp5_ASAP7_75t_L g11659 ( 
.A(n_10869),
.B(n_9978),
.Y(n_11659)
);

INVx6_ASAP7_75t_L g11660 ( 
.A(n_10425),
.Y(n_11660)
);

OR2x2_ASAP7_75t_L g11661 ( 
.A(n_11417),
.B(n_10085),
.Y(n_11661)
);

INVx2_ASAP7_75t_L g11662 ( 
.A(n_11204),
.Y(n_11662)
);

BUFx6f_ASAP7_75t_L g11663 ( 
.A(n_10425),
.Y(n_11663)
);

OAI22xp5_ASAP7_75t_SL g11664 ( 
.A1(n_11443),
.A2(n_9080),
.B1(n_9281),
.B2(n_9055),
.Y(n_11664)
);

NAND2xp5_ASAP7_75t_L g11665 ( 
.A(n_10520),
.B(n_10000),
.Y(n_11665)
);

AOI22xp33_ASAP7_75t_L g11666 ( 
.A1(n_11472),
.A2(n_9410),
.B1(n_9675),
.B2(n_9672),
.Y(n_11666)
);

OAI33xp33_ASAP7_75t_L g11667 ( 
.A1(n_10423),
.A2(n_9332),
.A3(n_9337),
.B1(n_7951),
.B2(n_8001),
.B3(n_7923),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_10382),
.Y(n_11668)
);

CKINVDCx20_ASAP7_75t_R g11669 ( 
.A(n_10702),
.Y(n_11669)
);

OAI22xp33_ASAP7_75t_L g11670 ( 
.A1(n_11397),
.A2(n_9702),
.B1(n_10006),
.B2(n_9986),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_SL g11671 ( 
.A(n_11178),
.B(n_9490),
.Y(n_11671)
);

AOI21xp5_ASAP7_75t_L g11672 ( 
.A1(n_11196),
.A2(n_9490),
.B(n_9080),
.Y(n_11672)
);

OAI22xp5_ASAP7_75t_L g11673 ( 
.A1(n_11448),
.A2(n_9568),
.B1(n_9314),
.B2(n_9340),
.Y(n_11673)
);

OAI21xp33_ASAP7_75t_L g11674 ( 
.A1(n_10733),
.A2(n_9759),
.B(n_9390),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_11204),
.Y(n_11675)
);

BUFx4f_ASAP7_75t_L g11676 ( 
.A(n_10454),
.Y(n_11676)
);

AND2x4_ASAP7_75t_L g11677 ( 
.A(n_10915),
.B(n_9114),
.Y(n_11677)
);

BUFx3_ASAP7_75t_L g11678 ( 
.A(n_10702),
.Y(n_11678)
);

NOR2xp33_ASAP7_75t_L g11679 ( 
.A(n_10886),
.B(n_9055),
.Y(n_11679)
);

AOI22xp33_ASAP7_75t_L g11680 ( 
.A1(n_10602),
.A2(n_9928),
.B1(n_10174),
.B2(n_9675),
.Y(n_11680)
);

BUFx12f_ASAP7_75t_L g11681 ( 
.A(n_11011),
.Y(n_11681)
);

OAI211xp5_ASAP7_75t_L g11682 ( 
.A1(n_10733),
.A2(n_10290),
.B(n_9099),
.C(n_9497),
.Y(n_11682)
);

INVx1_ASAP7_75t_L g11683 ( 
.A(n_10384),
.Y(n_11683)
);

INVx3_ASAP7_75t_L g11684 ( 
.A(n_10558),
.Y(n_11684)
);

AOI21xp5_ASAP7_75t_L g11685 ( 
.A1(n_11196),
.A2(n_9490),
.B(n_9281),
.Y(n_11685)
);

INVx2_ASAP7_75t_L g11686 ( 
.A(n_11221),
.Y(n_11686)
);

INVxp67_ASAP7_75t_L g11687 ( 
.A(n_10977),
.Y(n_11687)
);

NAND2xp5_ASAP7_75t_L g11688 ( 
.A(n_10697),
.B(n_10000),
.Y(n_11688)
);

AOI22xp33_ASAP7_75t_SL g11689 ( 
.A1(n_11080),
.A2(n_7815),
.B1(n_9723),
.B2(n_9157),
.Y(n_11689)
);

AND2x2_ASAP7_75t_L g11690 ( 
.A(n_11190),
.B(n_10499),
.Y(n_11690)
);

OAI22xp5_ASAP7_75t_L g11691 ( 
.A1(n_10825),
.A2(n_9201),
.B1(n_9240),
.B2(n_9649),
.Y(n_11691)
);

NOR2xp33_ASAP7_75t_L g11692 ( 
.A(n_10886),
.B(n_9080),
.Y(n_11692)
);

OAI211xp5_ASAP7_75t_L g11693 ( 
.A1(n_10825),
.A2(n_9491),
.B(n_9829),
.C(n_9731),
.Y(n_11693)
);

OAI22xp33_ASAP7_75t_L g11694 ( 
.A1(n_10402),
.A2(n_10006),
.B1(n_10030),
.B2(n_9986),
.Y(n_11694)
);

INVx2_ASAP7_75t_L g11695 ( 
.A(n_11221),
.Y(n_11695)
);

AOI22xp33_ASAP7_75t_SL g11696 ( 
.A1(n_10667),
.A2(n_7815),
.B1(n_9157),
.B2(n_9110),
.Y(n_11696)
);

AOI21xp33_ASAP7_75t_L g11697 ( 
.A1(n_11017),
.A2(n_9748),
.B(n_9086),
.Y(n_11697)
);

AOI22xp33_ASAP7_75t_L g11698 ( 
.A1(n_10602),
.A2(n_9928),
.B1(n_10174),
.B2(n_9675),
.Y(n_11698)
);

OA21x2_ASAP7_75t_L g11699 ( 
.A1(n_11116),
.A2(n_9399),
.B(n_9398),
.Y(n_11699)
);

OR2x6_ASAP7_75t_L g11700 ( 
.A(n_11243),
.B(n_9212),
.Y(n_11700)
);

AOI22xp33_ASAP7_75t_L g11701 ( 
.A1(n_10421),
.A2(n_9928),
.B1(n_10174),
.B2(n_9675),
.Y(n_11701)
);

NAND2xp5_ASAP7_75t_L g11702 ( 
.A(n_10717),
.B(n_10046),
.Y(n_11702)
);

OAI22xp5_ASAP7_75t_L g11703 ( 
.A1(n_11017),
.A2(n_9938),
.B1(n_9971),
.B2(n_9946),
.Y(n_11703)
);

A2O1A1Ixp33_ASAP7_75t_L g11704 ( 
.A1(n_11443),
.A2(n_10178),
.B(n_10146),
.C(n_8686),
.Y(n_11704)
);

AND2x2_ASAP7_75t_L g11705 ( 
.A(n_10499),
.B(n_9555),
.Y(n_11705)
);

AND2x2_ASAP7_75t_L g11706 ( 
.A(n_10512),
.B(n_9555),
.Y(n_11706)
);

HB1xp67_ASAP7_75t_L g11707 ( 
.A(n_11519),
.Y(n_11707)
);

AND2x4_ASAP7_75t_L g11708 ( 
.A(n_10934),
.B(n_9114),
.Y(n_11708)
);

INVx2_ASAP7_75t_L g11709 ( 
.A(n_11246),
.Y(n_11709)
);

OAI22xp5_ASAP7_75t_L g11710 ( 
.A1(n_10622),
.A2(n_9848),
.B1(n_9853),
.B2(n_9936),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_10388),
.Y(n_11711)
);

OR2x2_ASAP7_75t_L g11712 ( 
.A(n_10389),
.B(n_11271),
.Y(n_11712)
);

AND2x2_ASAP7_75t_L g11713 ( 
.A(n_10512),
.B(n_10515),
.Y(n_11713)
);

AOI22xp33_ASAP7_75t_L g11714 ( 
.A1(n_10481),
.A2(n_9928),
.B1(n_10174),
.B2(n_9675),
.Y(n_11714)
);

OAI22xp33_ASAP7_75t_L g11715 ( 
.A1(n_10402),
.A2(n_10006),
.B1(n_10030),
.B2(n_9986),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_10515),
.B(n_9623),
.Y(n_11716)
);

OAI211xp5_ASAP7_75t_L g11717 ( 
.A1(n_11346),
.A2(n_9908),
.B(n_9906),
.C(n_9527),
.Y(n_11717)
);

INVx1_ASAP7_75t_L g11718 ( 
.A(n_10394),
.Y(n_11718)
);

AOI22xp33_ASAP7_75t_L g11719 ( 
.A1(n_10482),
.A2(n_10174),
.B1(n_10220),
.B2(n_9928),
.Y(n_11719)
);

AOI22xp33_ASAP7_75t_L g11720 ( 
.A1(n_10490),
.A2(n_10220),
.B1(n_10312),
.B2(n_9739),
.Y(n_11720)
);

AOI22xp33_ASAP7_75t_L g11721 ( 
.A1(n_10532),
.A2(n_10220),
.B1(n_10312),
.B2(n_9736),
.Y(n_11721)
);

OA21x2_ASAP7_75t_L g11722 ( 
.A1(n_10924),
.A2(n_10958),
.B(n_10914),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_10399),
.Y(n_11723)
);

OAI21x1_ASAP7_75t_L g11724 ( 
.A1(n_10451),
.A2(n_10353),
.B(n_10328),
.Y(n_11724)
);

HB1xp67_ASAP7_75t_L g11725 ( 
.A(n_11534),
.Y(n_11725)
);

AND2x2_ASAP7_75t_L g11726 ( 
.A(n_10518),
.B(n_9623),
.Y(n_11726)
);

OAI22xp33_ASAP7_75t_L g11727 ( 
.A1(n_10402),
.A2(n_10031),
.B1(n_10064),
.B2(n_10030),
.Y(n_11727)
);

OA21x2_ASAP7_75t_L g11728 ( 
.A1(n_10924),
.A2(n_9399),
.B(n_9398),
.Y(n_11728)
);

AOI21xp33_ASAP7_75t_L g11729 ( 
.A1(n_10478),
.A2(n_9748),
.B(n_10196),
.Y(n_11729)
);

BUFx2_ASAP7_75t_L g11730 ( 
.A(n_11178),
.Y(n_11730)
);

AOI22xp33_ASAP7_75t_SL g11731 ( 
.A1(n_10410),
.A2(n_7815),
.B1(n_9157),
.B2(n_9110),
.Y(n_11731)
);

AOI221xp5_ASAP7_75t_L g11732 ( 
.A1(n_10549),
.A2(n_9748),
.B1(n_9332),
.B2(n_9337),
.C(n_9546),
.Y(n_11732)
);

NOR2xp33_ASAP7_75t_L g11733 ( 
.A(n_10900),
.B(n_9281),
.Y(n_11733)
);

INVx2_ASAP7_75t_SL g11734 ( 
.A(n_10599),
.Y(n_11734)
);

AOI222xp33_ASAP7_75t_L g11735 ( 
.A1(n_10530),
.A2(n_8508),
.B1(n_9020),
.B2(n_9281),
.C1(n_9285),
.C2(n_8980),
.Y(n_11735)
);

AOI22xp33_ASAP7_75t_L g11736 ( 
.A1(n_10566),
.A2(n_10220),
.B1(n_9110),
.B2(n_9173),
.Y(n_11736)
);

NAND3xp33_ASAP7_75t_L g11737 ( 
.A(n_11092),
.B(n_10245),
.C(n_10196),
.Y(n_11737)
);

AOI22xp33_ASAP7_75t_SL g11738 ( 
.A1(n_10410),
.A2(n_7815),
.B1(n_9157),
.B2(n_9110),
.Y(n_11738)
);

AND2x4_ASAP7_75t_L g11739 ( 
.A(n_10974),
.B(n_11027),
.Y(n_11739)
);

AOI22xp33_ASAP7_75t_L g11740 ( 
.A1(n_10604),
.A2(n_10220),
.B1(n_9157),
.B2(n_9188),
.Y(n_11740)
);

AOI22xp33_ASAP7_75t_SL g11741 ( 
.A1(n_10410),
.A2(n_10562),
.B1(n_11289),
.B2(n_11107),
.Y(n_11741)
);

CKINVDCx5p33_ASAP7_75t_R g11742 ( 
.A(n_11011),
.Y(n_11742)
);

AOI221xp5_ASAP7_75t_L g11743 ( 
.A1(n_10524),
.A2(n_9527),
.B1(n_9725),
.B2(n_9609),
.C(n_9552),
.Y(n_11743)
);

INVx1_ASAP7_75t_L g11744 ( 
.A(n_10400),
.Y(n_11744)
);

AOI21xp33_ASAP7_75t_L g11745 ( 
.A1(n_11127),
.A2(n_10245),
.B(n_10196),
.Y(n_11745)
);

OR2x2_ASAP7_75t_L g11746 ( 
.A(n_11433),
.B(n_10085),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_10409),
.Y(n_11747)
);

INVx2_ASAP7_75t_L g11748 ( 
.A(n_11246),
.Y(n_11748)
);

OAI22xp5_ASAP7_75t_L g11749 ( 
.A1(n_10727),
.A2(n_8673),
.B1(n_9948),
.B2(n_10040),
.Y(n_11749)
);

NAND3xp33_ASAP7_75t_L g11750 ( 
.A(n_11092),
.B(n_10245),
.C(n_10196),
.Y(n_11750)
);

CKINVDCx11_ASAP7_75t_R g11751 ( 
.A(n_10454),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_10413),
.Y(n_11752)
);

AOI22xp33_ASAP7_75t_L g11753 ( 
.A1(n_10614),
.A2(n_9173),
.B1(n_9190),
.B2(n_9188),
.Y(n_11753)
);

CKINVDCx20_ASAP7_75t_R g11754 ( 
.A(n_10900),
.Y(n_11754)
);

OAI21xp5_ASAP7_75t_SL g11755 ( 
.A1(n_10940),
.A2(n_10972),
.B(n_11222),
.Y(n_11755)
);

OAI21x1_ASAP7_75t_L g11756 ( 
.A1(n_10464),
.A2(n_10353),
.B(n_10328),
.Y(n_11756)
);

AOI22xp33_ASAP7_75t_L g11757 ( 
.A1(n_10615),
.A2(n_9173),
.B1(n_9190),
.B2(n_9188),
.Y(n_11757)
);

BUFx6f_ASAP7_75t_L g11758 ( 
.A(n_10613),
.Y(n_11758)
);

INVx3_ASAP7_75t_L g11759 ( 
.A(n_10558),
.Y(n_11759)
);

AOI22xp33_ASAP7_75t_L g11760 ( 
.A1(n_11083),
.A2(n_9173),
.B1(n_9190),
.B2(n_9188),
.Y(n_11760)
);

INVx1_ASAP7_75t_L g11761 ( 
.A(n_10414),
.Y(n_11761)
);

AOI22xp33_ASAP7_75t_L g11762 ( 
.A1(n_10972),
.A2(n_11262),
.B1(n_11277),
.B2(n_11275),
.Y(n_11762)
);

INVx1_ASAP7_75t_L g11763 ( 
.A(n_10419),
.Y(n_11763)
);

AO31x2_ASAP7_75t_L g11764 ( 
.A1(n_11503),
.A2(n_9285),
.A3(n_10245),
.B(n_9335),
.Y(n_11764)
);

OAI22xp5_ASAP7_75t_L g11765 ( 
.A1(n_11183),
.A2(n_10136),
.B1(n_10070),
.B2(n_9989),
.Y(n_11765)
);

BUFx4f_ASAP7_75t_L g11766 ( 
.A(n_10599),
.Y(n_11766)
);

AOI22xp5_ASAP7_75t_L g11767 ( 
.A1(n_11262),
.A2(n_10347),
.B1(n_9173),
.B2(n_9190),
.Y(n_11767)
);

OAI22xp5_ASAP7_75t_L g11768 ( 
.A1(n_11239),
.A2(n_11241),
.B1(n_11281),
.B2(n_11255),
.Y(n_11768)
);

NAND2xp5_ASAP7_75t_L g11769 ( 
.A(n_10921),
.B(n_10046),
.Y(n_11769)
);

INVx2_ASAP7_75t_L g11770 ( 
.A(n_11277),
.Y(n_11770)
);

INVx1_ASAP7_75t_L g11771 ( 
.A(n_10427),
.Y(n_11771)
);

AOI221xp5_ASAP7_75t_L g11772 ( 
.A1(n_10581),
.A2(n_9552),
.B1(n_9812),
.B2(n_9725),
.C(n_9609),
.Y(n_11772)
);

AND2x4_ASAP7_75t_SL g11773 ( 
.A(n_11120),
.B(n_9718),
.Y(n_11773)
);

AOI22xp33_ASAP7_75t_SL g11774 ( 
.A1(n_10920),
.A2(n_10859),
.B1(n_10599),
.B2(n_11314),
.Y(n_11774)
);

INVx2_ASAP7_75t_L g11775 ( 
.A(n_11382),
.Y(n_11775)
);

A2O1A1Ixp33_ASAP7_75t_L g11776 ( 
.A1(n_11377),
.A2(n_11540),
.B(n_11488),
.C(n_11162),
.Y(n_11776)
);

AO21x2_ASAP7_75t_L g11777 ( 
.A1(n_11143),
.A2(n_9864),
.B(n_10292),
.Y(n_11777)
);

INVx1_ASAP7_75t_L g11778 ( 
.A(n_10428),
.Y(n_11778)
);

AND2x4_ASAP7_75t_L g11779 ( 
.A(n_11412),
.B(n_9290),
.Y(n_11779)
);

INVx1_ASAP7_75t_SL g11780 ( 
.A(n_10803),
.Y(n_11780)
);

AOI22xp33_ASAP7_75t_L g11781 ( 
.A1(n_11532),
.A2(n_9188),
.B1(n_9216),
.B2(n_9190),
.Y(n_11781)
);

OAI22xp5_ASAP7_75t_L g11782 ( 
.A1(n_11135),
.A2(n_9192),
.B1(n_9171),
.B2(n_9000),
.Y(n_11782)
);

INVx2_ASAP7_75t_L g11783 ( 
.A(n_11382),
.Y(n_11783)
);

AOI221xp5_ASAP7_75t_L g11784 ( 
.A1(n_10640),
.A2(n_9812),
.B1(n_9864),
.B2(n_8642),
.C(n_8686),
.Y(n_11784)
);

AOI22xp5_ASAP7_75t_L g11785 ( 
.A1(n_11412),
.A2(n_9216),
.B1(n_9302),
.B2(n_9263),
.Y(n_11785)
);

NAND2xp5_ASAP7_75t_L g11786 ( 
.A(n_10996),
.B(n_10159),
.Y(n_11786)
);

INVxp67_ASAP7_75t_SL g11787 ( 
.A(n_11457),
.Y(n_11787)
);

INVx1_ASAP7_75t_L g11788 ( 
.A(n_10430),
.Y(n_11788)
);

OAI221xp5_ASAP7_75t_L g11789 ( 
.A1(n_11516),
.A2(n_9913),
.B1(n_9766),
.B2(n_9624),
.C(n_9285),
.Y(n_11789)
);

OAI22xp33_ASAP7_75t_L g11790 ( 
.A1(n_11135),
.A2(n_10031),
.B1(n_10064),
.B2(n_8942),
.Y(n_11790)
);

AOI22xp33_ASAP7_75t_SL g11791 ( 
.A1(n_10920),
.A2(n_9263),
.B1(n_9302),
.B2(n_9216),
.Y(n_11791)
);

INVx1_ASAP7_75t_L g11792 ( 
.A(n_10431),
.Y(n_11792)
);

OAI22xp5_ASAP7_75t_L g11793 ( 
.A1(n_11135),
.A2(n_9000),
.B1(n_8997),
.B2(n_9357),
.Y(n_11793)
);

OAI21xp5_ASAP7_75t_L g11794 ( 
.A1(n_11528),
.A2(n_7902),
.B(n_9844),
.Y(n_11794)
);

AOI22xp33_ASAP7_75t_L g11795 ( 
.A1(n_11387),
.A2(n_9263),
.B1(n_9302),
.B2(n_9216),
.Y(n_11795)
);

BUFx4f_ASAP7_75t_SL g11796 ( 
.A(n_10390),
.Y(n_11796)
);

AOI222xp33_ASAP7_75t_L g11797 ( 
.A1(n_11230),
.A2(n_8508),
.B1(n_9285),
.B2(n_8407),
.C1(n_8984),
.C2(n_8781),
.Y(n_11797)
);

OA21x2_ASAP7_75t_L g11798 ( 
.A1(n_10426),
.A2(n_9401),
.B(n_9399),
.Y(n_11798)
);

AND2x2_ASAP7_75t_L g11799 ( 
.A(n_10518),
.B(n_9656),
.Y(n_11799)
);

NAND2xp5_ASAP7_75t_L g11800 ( 
.A(n_11015),
.B(n_10159),
.Y(n_11800)
);

INVx1_ASAP7_75t_L g11801 ( 
.A(n_10439),
.Y(n_11801)
);

HB1xp67_ASAP7_75t_L g11802 ( 
.A(n_10674),
.Y(n_11802)
);

NOR2x1_ASAP7_75t_SL g11803 ( 
.A(n_11135),
.B(n_9713),
.Y(n_11803)
);

INVx4_ASAP7_75t_L g11804 ( 
.A(n_10398),
.Y(n_11804)
);

AOI22xp33_ASAP7_75t_L g11805 ( 
.A1(n_11387),
.A2(n_9263),
.B1(n_9302),
.B2(n_9216),
.Y(n_11805)
);

AOI22xp33_ASAP7_75t_L g11806 ( 
.A1(n_11400),
.A2(n_9302),
.B1(n_9313),
.B2(n_9263),
.Y(n_11806)
);

OAI21x1_ASAP7_75t_L g11807 ( 
.A1(n_10570),
.A2(n_10353),
.B(n_10328),
.Y(n_11807)
);

OAI22xp33_ASAP7_75t_L g11808 ( 
.A1(n_11535),
.A2(n_10031),
.B1(n_10064),
.B2(n_8942),
.Y(n_11808)
);

AND2x2_ASAP7_75t_L g11809 ( 
.A(n_10542),
.B(n_9656),
.Y(n_11809)
);

OAI22xp33_ASAP7_75t_SL g11810 ( 
.A1(n_10691),
.A2(n_9827),
.B1(n_9313),
.B2(n_10126),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_10440),
.Y(n_11811)
);

AOI221xp5_ASAP7_75t_L g11812 ( 
.A1(n_11058),
.A2(n_9864),
.B1(n_9230),
.B2(n_8904),
.C(n_8911),
.Y(n_11812)
);

AOI22xp5_ASAP7_75t_L g11813 ( 
.A1(n_11514),
.A2(n_9313),
.B1(n_8192),
.B2(n_10043),
.Y(n_11813)
);

AOI221xp5_ASAP7_75t_L g11814 ( 
.A1(n_11081),
.A2(n_9864),
.B1(n_9230),
.B2(n_8904),
.C(n_8911),
.Y(n_11814)
);

OAI211xp5_ASAP7_75t_L g11815 ( 
.A1(n_10826),
.A2(n_7832),
.B(n_7747),
.C(n_10207),
.Y(n_11815)
);

AOI222xp33_ASAP7_75t_L g11816 ( 
.A1(n_11480),
.A2(n_8699),
.B1(n_8781),
.B2(n_8729),
.C1(n_8505),
.C2(n_8576),
.Y(n_11816)
);

INVx1_ASAP7_75t_SL g11817 ( 
.A(n_10548),
.Y(n_11817)
);

OAI211xp5_ASAP7_75t_SL g11818 ( 
.A1(n_11106),
.A2(n_11206),
.B(n_11475),
.C(n_11317),
.Y(n_11818)
);

INVx1_ASAP7_75t_L g11819 ( 
.A(n_10443),
.Y(n_11819)
);

OAI22xp33_ASAP7_75t_L g11820 ( 
.A1(n_11535),
.A2(n_9022),
.B1(n_8275),
.B2(n_9449),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_10444),
.Y(n_11821)
);

AO21x2_ASAP7_75t_L g11822 ( 
.A1(n_10956),
.A2(n_10835),
.B(n_10859),
.Y(n_11822)
);

INVx2_ASAP7_75t_L g11823 ( 
.A(n_10420),
.Y(n_11823)
);

OAI322xp33_ASAP7_75t_L g11824 ( 
.A1(n_11106),
.A2(n_11317),
.A3(n_11475),
.B1(n_11476),
.B2(n_11206),
.C1(n_11529),
.C2(n_11509),
.Y(n_11824)
);

AOI22xp33_ASAP7_75t_L g11825 ( 
.A1(n_11402),
.A2(n_11435),
.B1(n_11409),
.B2(n_10676),
.Y(n_11825)
);

INVx1_ASAP7_75t_L g11826 ( 
.A(n_10447),
.Y(n_11826)
);

AOI22xp33_ASAP7_75t_L g11827 ( 
.A1(n_10628),
.A2(n_9313),
.B1(n_10137),
.B2(n_10126),
.Y(n_11827)
);

OAI21x1_ASAP7_75t_L g11828 ( 
.A1(n_10570),
.A2(n_9461),
.B(n_9388),
.Y(n_11828)
);

OAI22xp33_ASAP7_75t_L g11829 ( 
.A1(n_11535),
.A2(n_10691),
.B1(n_10765),
.B2(n_11328),
.Y(n_11829)
);

AOI22xp33_ASAP7_75t_L g11830 ( 
.A1(n_10680),
.A2(n_9313),
.B1(n_10137),
.B2(n_10126),
.Y(n_11830)
);

CKINVDCx5p33_ASAP7_75t_R g11831 ( 
.A(n_11522),
.Y(n_11831)
);

AOI22xp33_ASAP7_75t_SL g11832 ( 
.A1(n_10767),
.A2(n_9212),
.B1(n_9210),
.B2(n_8590),
.Y(n_11832)
);

AOI22xp33_ASAP7_75t_SL g11833 ( 
.A1(n_10767),
.A2(n_10719),
.B1(n_10386),
.B2(n_10395),
.Y(n_11833)
);

INVx5_ASAP7_75t_SL g11834 ( 
.A(n_10613),
.Y(n_11834)
);

AOI222xp33_ASAP7_75t_L g11835 ( 
.A1(n_11411),
.A2(n_8729),
.B1(n_8533),
.B2(n_9693),
.C1(n_8517),
.C2(n_9212),
.Y(n_11835)
);

AOI22xp33_ASAP7_75t_L g11836 ( 
.A1(n_10808),
.A2(n_10137),
.B1(n_10200),
.B2(n_10167),
.Y(n_11836)
);

AOI21xp33_ASAP7_75t_L g11837 ( 
.A1(n_10691),
.A2(n_10200),
.B(n_10167),
.Y(n_11837)
);

AOI22xp33_ASAP7_75t_L g11838 ( 
.A1(n_10851),
.A2(n_10167),
.B1(n_10200),
.B2(n_10043),
.Y(n_11838)
);

OAI22xp33_ASAP7_75t_L g11839 ( 
.A1(n_11535),
.A2(n_9022),
.B1(n_9449),
.B2(n_9764),
.Y(n_11839)
);

INVx3_ASAP7_75t_L g11840 ( 
.A(n_10715),
.Y(n_11840)
);

INVx1_ASAP7_75t_L g11841 ( 
.A(n_10448),
.Y(n_11841)
);

OAI221xp5_ASAP7_75t_L g11842 ( 
.A1(n_11293),
.A2(n_9631),
.B1(n_9689),
.B2(n_9683),
.C(n_9377),
.Y(n_11842)
);

OAI22xp33_ASAP7_75t_L g11843 ( 
.A1(n_10691),
.A2(n_9449),
.B1(n_9984),
.B2(n_9764),
.Y(n_11843)
);

INVx1_ASAP7_75t_L g11844 ( 
.A(n_10463),
.Y(n_11844)
);

AOI22xp33_ASAP7_75t_SL g11845 ( 
.A1(n_10719),
.A2(n_8590),
.B1(n_8604),
.B2(n_7957),
.Y(n_11845)
);

OAI22xp33_ASAP7_75t_SL g11846 ( 
.A1(n_10765),
.A2(n_9827),
.B1(n_9751),
.B2(n_9745),
.Y(n_11846)
);

AOI221xp5_ASAP7_75t_SL g11847 ( 
.A1(n_10403),
.A2(n_8447),
.B1(n_8617),
.B2(n_8476),
.C(n_8428),
.Y(n_11847)
);

AND2x2_ASAP7_75t_L g11848 ( 
.A(n_10542),
.B(n_9745),
.Y(n_11848)
);

OR2x2_ASAP7_75t_L g11849 ( 
.A(n_10552),
.B(n_9462),
.Y(n_11849)
);

INVx3_ASAP7_75t_L g11850 ( 
.A(n_10715),
.Y(n_11850)
);

OAI22xp5_ASAP7_75t_L g11851 ( 
.A1(n_11514),
.A2(n_11539),
.B1(n_10765),
.B2(n_8997),
.Y(n_11851)
);

OAI221xp5_ASAP7_75t_L g11852 ( 
.A1(n_11293),
.A2(n_9786),
.B1(n_9355),
.B2(n_10204),
.C(n_10315),
.Y(n_11852)
);

OAI22xp33_ASAP7_75t_L g11853 ( 
.A1(n_10765),
.A2(n_9449),
.B1(n_9984),
.B2(n_9764),
.Y(n_11853)
);

INVx1_ASAP7_75t_L g11854 ( 
.A(n_10466),
.Y(n_11854)
);

AOI221xp5_ASAP7_75t_L g11855 ( 
.A1(n_11095),
.A2(n_9230),
.B1(n_8928),
.B2(n_8344),
.C(n_8947),
.Y(n_11855)
);

BUFx6f_ASAP7_75t_L g11856 ( 
.A(n_10613),
.Y(n_11856)
);

OA21x2_ASAP7_75t_L g11857 ( 
.A1(n_10426),
.A2(n_9411),
.B(n_9401),
.Y(n_11857)
);

INVx2_ASAP7_75t_L g11858 ( 
.A(n_10420),
.Y(n_11858)
);

AOI221xp5_ASAP7_75t_L g11859 ( 
.A1(n_11098),
.A2(n_9230),
.B1(n_8928),
.B2(n_8344),
.C(n_8947),
.Y(n_11859)
);

INVx2_ASAP7_75t_L g11860 ( 
.A(n_10420),
.Y(n_11860)
);

AND2x2_ASAP7_75t_L g11861 ( 
.A(n_10544),
.B(n_9751),
.Y(n_11861)
);

AO21x1_ASAP7_75t_SL g11862 ( 
.A1(n_10725),
.A2(n_10237),
.B(n_10235),
.Y(n_11862)
);

INVx1_ASAP7_75t_L g11863 ( 
.A(n_10475),
.Y(n_11863)
);

AOI22xp33_ASAP7_75t_SL g11864 ( 
.A1(n_10386),
.A2(n_8604),
.B1(n_7957),
.B2(n_8977),
.Y(n_11864)
);

OAI21x1_ASAP7_75t_L g11865 ( 
.A1(n_10811),
.A2(n_9461),
.B(n_9388),
.Y(n_11865)
);

INVx1_ASAP7_75t_L g11866 ( 
.A(n_10476),
.Y(n_11866)
);

OAI211xp5_ASAP7_75t_L g11867 ( 
.A1(n_11092),
.A2(n_7832),
.B(n_7747),
.C(n_10241),
.Y(n_11867)
);

OR2x2_ASAP7_75t_L g11868 ( 
.A(n_10784),
.B(n_9462),
.Y(n_11868)
);

OAI22xp5_ASAP7_75t_L g11869 ( 
.A1(n_11539),
.A2(n_10250),
.B1(n_10139),
.B2(n_10069),
.Y(n_11869)
);

AOI22xp33_ASAP7_75t_L g11870 ( 
.A1(n_10853),
.A2(n_10043),
.B1(n_10108),
.B2(n_9996),
.Y(n_11870)
);

AND2x2_ASAP7_75t_L g11871 ( 
.A(n_10544),
.B(n_9911),
.Y(n_11871)
);

OR2x6_ASAP7_75t_L g11872 ( 
.A(n_11030),
.B(n_9290),
.Y(n_11872)
);

OAI22xp5_ASAP7_75t_L g11873 ( 
.A1(n_11128),
.A2(n_10139),
.B1(n_10069),
.B2(n_10133),
.Y(n_11873)
);

INVx4_ASAP7_75t_L g11874 ( 
.A(n_10398),
.Y(n_11874)
);

BUFx12f_ASAP7_75t_L g11875 ( 
.A(n_11522),
.Y(n_11875)
);

OAI22xp33_ASAP7_75t_L g11876 ( 
.A1(n_11328),
.A2(n_9449),
.B1(n_9984),
.B2(n_9764),
.Y(n_11876)
);

AOI211xp5_ASAP7_75t_L g11877 ( 
.A1(n_11379),
.A2(n_8427),
.B(n_8063),
.C(n_7979),
.Y(n_11877)
);

AND2x2_ASAP7_75t_L g11878 ( 
.A(n_10554),
.B(n_9911),
.Y(n_11878)
);

AND2x2_ASAP7_75t_SL g11879 ( 
.A(n_10898),
.B(n_9706),
.Y(n_11879)
);

AOI22xp33_ASAP7_75t_L g11880 ( 
.A1(n_10904),
.A2(n_10108),
.B1(n_10184),
.B2(n_9996),
.Y(n_11880)
);

NAND2xp5_ASAP7_75t_L g11881 ( 
.A(n_11253),
.B(n_10221),
.Y(n_11881)
);

OAI221xp5_ASAP7_75t_L g11882 ( 
.A1(n_11379),
.A2(n_9121),
.B1(n_9274),
.B2(n_9045),
.C(n_10121),
.Y(n_11882)
);

OAI22xp5_ASAP7_75t_L g11883 ( 
.A1(n_11290),
.A2(n_11282),
.B1(n_11465),
.B2(n_10416),
.Y(n_11883)
);

AOI21xp33_ASAP7_75t_SL g11884 ( 
.A1(n_10548),
.A2(n_9223),
.B(n_9140),
.Y(n_11884)
);

AOI22xp33_ASAP7_75t_L g11885 ( 
.A1(n_10613),
.A2(n_10108),
.B1(n_10184),
.B2(n_9996),
.Y(n_11885)
);

OAI211xp5_ASAP7_75t_SL g11886 ( 
.A1(n_11476),
.A2(n_9467),
.B(n_9820),
.C(n_9674),
.Y(n_11886)
);

BUFx2_ASAP7_75t_L g11887 ( 
.A(n_10390),
.Y(n_11887)
);

AND2x2_ASAP7_75t_L g11888 ( 
.A(n_10554),
.B(n_9952),
.Y(n_11888)
);

OAI21x1_ASAP7_75t_L g11889 ( 
.A1(n_10811),
.A2(n_9543),
.B(n_9506),
.Y(n_11889)
);

INVx3_ASAP7_75t_L g11890 ( 
.A(n_11001),
.Y(n_11890)
);

OAI21x1_ASAP7_75t_L g11891 ( 
.A1(n_11001),
.A2(n_9543),
.B(n_9506),
.Y(n_11891)
);

OAI22xp5_ASAP7_75t_L g11892 ( 
.A1(n_10408),
.A2(n_10160),
.B1(n_10158),
.B2(n_8843),
.Y(n_11892)
);

AND2x2_ASAP7_75t_L g11893 ( 
.A(n_10557),
.B(n_9952),
.Y(n_11893)
);

AOI22xp33_ASAP7_75t_SL g11894 ( 
.A1(n_10395),
.A2(n_7957),
.B1(n_7747),
.B2(n_7832),
.Y(n_11894)
);

OAI22xp5_ASAP7_75t_L g11895 ( 
.A1(n_10408),
.A2(n_8843),
.B1(n_8892),
.B2(n_8878),
.Y(n_11895)
);

BUFx3_ASAP7_75t_L g11896 ( 
.A(n_10461),
.Y(n_11896)
);

AOI211x1_ASAP7_75t_L g11897 ( 
.A1(n_10785),
.A2(n_8706),
.B(n_9891),
.C(n_9844),
.Y(n_11897)
);

INVx1_ASAP7_75t_L g11898 ( 
.A(n_10479),
.Y(n_11898)
);

INVx3_ASAP7_75t_L g11899 ( 
.A(n_11457),
.Y(n_11899)
);

AOI22xp33_ASAP7_75t_L g11900 ( 
.A1(n_10623),
.A2(n_10239),
.B1(n_10369),
.B2(n_10184),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_10483),
.Y(n_11901)
);

INVx1_ASAP7_75t_L g11902 ( 
.A(n_10489),
.Y(n_11902)
);

OAI22xp33_ASAP7_75t_L g11903 ( 
.A1(n_11328),
.A2(n_9984),
.B1(n_10117),
.B2(n_9764),
.Y(n_11903)
);

OAI22xp5_ASAP7_75t_L g11904 ( 
.A1(n_10416),
.A2(n_8878),
.B1(n_8892),
.B2(n_10225),
.Y(n_11904)
);

AOI221xp5_ASAP7_75t_L g11905 ( 
.A1(n_11509),
.A2(n_8869),
.B1(n_8807),
.B2(n_9836),
.C(n_9835),
.Y(n_11905)
);

AND2x2_ASAP7_75t_L g11906 ( 
.A(n_10557),
.B(n_9957),
.Y(n_11906)
);

HB1xp67_ASAP7_75t_L g11907 ( 
.A(n_10751),
.Y(n_11907)
);

OR2x2_ASAP7_75t_L g11908 ( 
.A(n_10793),
.B(n_9505),
.Y(n_11908)
);

INVx2_ASAP7_75t_L g11909 ( 
.A(n_10424),
.Y(n_11909)
);

OAI22xp5_ASAP7_75t_L g11910 ( 
.A1(n_10417),
.A2(n_10214),
.B1(n_8880),
.B2(n_8325),
.Y(n_11910)
);

NAND2xp5_ASAP7_75t_L g11911 ( 
.A(n_11504),
.B(n_10221),
.Y(n_11911)
);

AOI22xp33_ASAP7_75t_L g11912 ( 
.A1(n_10623),
.A2(n_10369),
.B1(n_10239),
.B2(n_9498),
.Y(n_11912)
);

AOI22xp33_ASAP7_75t_L g11913 ( 
.A1(n_10623),
.A2(n_10369),
.B1(n_10239),
.B2(n_9498),
.Y(n_11913)
);

AOI22xp33_ASAP7_75t_L g11914 ( 
.A1(n_10623),
.A2(n_9498),
.B1(n_9574),
.B2(n_9571),
.Y(n_11914)
);

OR2x2_ASAP7_75t_SL g11915 ( 
.A(n_10703),
.B(n_8961),
.Y(n_11915)
);

AOI22xp5_ASAP7_75t_L g11916 ( 
.A1(n_11446),
.A2(n_9969),
.B1(n_10052),
.B2(n_9957),
.Y(n_11916)
);

AOI22xp33_ASAP7_75t_L g11917 ( 
.A1(n_10703),
.A2(n_9571),
.B1(n_9587),
.B2(n_9574),
.Y(n_11917)
);

HB1xp67_ASAP7_75t_L g11918 ( 
.A(n_10786),
.Y(n_11918)
);

AOI22xp5_ASAP7_75t_L g11919 ( 
.A1(n_11446),
.A2(n_10052),
.B1(n_10063),
.B2(n_9969),
.Y(n_11919)
);

INVx1_ASAP7_75t_L g11920 ( 
.A(n_10500),
.Y(n_11920)
);

INVx2_ASAP7_75t_L g11921 ( 
.A(n_10424),
.Y(n_11921)
);

AOI22xp33_ASAP7_75t_L g11922 ( 
.A1(n_10703),
.A2(n_9571),
.B1(n_9587),
.B2(n_9574),
.Y(n_11922)
);

AOI22xp33_ASAP7_75t_L g11923 ( 
.A1(n_10703),
.A2(n_9587),
.B1(n_9650),
.B2(n_9628),
.Y(n_11923)
);

OAI221xp5_ASAP7_75t_L g11924 ( 
.A1(n_11162),
.A2(n_9755),
.B1(n_9711),
.B2(n_9365),
.C(n_9469),
.Y(n_11924)
);

OAI22xp33_ASAP7_75t_L g11925 ( 
.A1(n_11328),
.A2(n_10117),
.B1(n_10190),
.B2(n_9984),
.Y(n_11925)
);

AOI22xp33_ASAP7_75t_L g11926 ( 
.A1(n_10830),
.A2(n_9628),
.B1(n_9669),
.B2(n_9650),
.Y(n_11926)
);

OAI21x1_ASAP7_75t_L g11927 ( 
.A1(n_11518),
.A2(n_9554),
.B(n_9277),
.Y(n_11927)
);

AOI22xp33_ASAP7_75t_L g11928 ( 
.A1(n_10830),
.A2(n_9628),
.B1(n_9669),
.B2(n_9650),
.Y(n_11928)
);

AOI22xp33_ASAP7_75t_L g11929 ( 
.A1(n_10830),
.A2(n_9680),
.B1(n_9686),
.B2(n_9669),
.Y(n_11929)
);

OAI22xp5_ASAP7_75t_L g11930 ( 
.A1(n_10417),
.A2(n_8880),
.B1(n_8989),
.B2(n_9290),
.Y(n_11930)
);

OAI211xp5_ASAP7_75t_L g11931 ( 
.A1(n_10473),
.A2(n_7832),
.B(n_7747),
.C(n_7841),
.Y(n_11931)
);

INVx2_ASAP7_75t_L g11932 ( 
.A(n_10424),
.Y(n_11932)
);

AOI22xp5_ASAP7_75t_L g11933 ( 
.A1(n_10435),
.A2(n_10081),
.B1(n_10095),
.B2(n_10063),
.Y(n_11933)
);

AOI22xp33_ASAP7_75t_SL g11934 ( 
.A1(n_10888),
.A2(n_7957),
.B1(n_7747),
.B2(n_7832),
.Y(n_11934)
);

AOI221xp5_ASAP7_75t_L g11935 ( 
.A1(n_11529),
.A2(n_8869),
.B1(n_8807),
.B2(n_9836),
.C(n_9835),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_10501),
.Y(n_11936)
);

CKINVDCx5p33_ASAP7_75t_R g11937 ( 
.A(n_10404),
.Y(n_11937)
);

AOI22xp33_ASAP7_75t_L g11938 ( 
.A1(n_10830),
.A2(n_9686),
.B1(n_9712),
.B2(n_9680),
.Y(n_11938)
);

OAI22xp5_ASAP7_75t_L g11939 ( 
.A1(n_10435),
.A2(n_10446),
.B1(n_10612),
.B2(n_10474),
.Y(n_11939)
);

AOI22xp33_ASAP7_75t_L g11940 ( 
.A1(n_10861),
.A2(n_9686),
.B1(n_9712),
.B2(n_9680),
.Y(n_11940)
);

AND2x4_ASAP7_75t_L g11941 ( 
.A(n_10835),
.B(n_9290),
.Y(n_11941)
);

AOI22xp33_ASAP7_75t_L g11942 ( 
.A1(n_10861),
.A2(n_9779),
.B1(n_9797),
.B2(n_9712),
.Y(n_11942)
);

HB1xp67_ASAP7_75t_L g11943 ( 
.A(n_10790),
.Y(n_11943)
);

INVx2_ASAP7_75t_SL g11944 ( 
.A(n_10398),
.Y(n_11944)
);

CKINVDCx5p33_ASAP7_75t_R g11945 ( 
.A(n_10404),
.Y(n_11945)
);

AND2x2_ASAP7_75t_L g11946 ( 
.A(n_10838),
.B(n_10081),
.Y(n_11946)
);

AO31x2_ASAP7_75t_L g11947 ( 
.A1(n_10473),
.A2(n_9365),
.A3(n_9469),
.B(n_9335),
.Y(n_11947)
);

AOI221xp5_ASAP7_75t_L g11948 ( 
.A1(n_10473),
.A2(n_9835),
.B1(n_9836),
.B2(n_10306),
.C(n_10294),
.Y(n_11948)
);

OAI21xp5_ASAP7_75t_SL g11949 ( 
.A1(n_10565),
.A2(n_8473),
.B(n_8458),
.Y(n_11949)
);

AND2x2_ASAP7_75t_L g11950 ( 
.A(n_10838),
.B(n_10095),
.Y(n_11950)
);

AOI22xp5_ASAP7_75t_L g11951 ( 
.A1(n_10446),
.A2(n_10166),
.B1(n_10170),
.B2(n_10097),
.Y(n_11951)
);

INVx1_ASAP7_75t_L g11952 ( 
.A(n_10502),
.Y(n_11952)
);

AOI22xp33_ASAP7_75t_L g11953 ( 
.A1(n_10861),
.A2(n_9797),
.B1(n_9816),
.B2(n_9779),
.Y(n_11953)
);

NOR2x1_ASAP7_75t_R g11954 ( 
.A(n_10612),
.B(n_9847),
.Y(n_11954)
);

AND2x2_ASAP7_75t_L g11955 ( 
.A(n_10468),
.B(n_10097),
.Y(n_11955)
);

OAI221xp5_ASAP7_75t_L g11956 ( 
.A1(n_11162),
.A2(n_9469),
.B1(n_9501),
.B2(n_9365),
.C(n_9335),
.Y(n_11956)
);

AOI221xp5_ASAP7_75t_L g11957 ( 
.A1(n_10592),
.A2(n_9835),
.B1(n_9836),
.B2(n_10365),
.C(n_10340),
.Y(n_11957)
);

AND2x4_ASAP7_75t_L g11958 ( 
.A(n_10835),
.B(n_11497),
.Y(n_11958)
);

INVx2_ASAP7_75t_L g11959 ( 
.A(n_10486),
.Y(n_11959)
);

NOR2xp33_ASAP7_75t_L g11960 ( 
.A(n_10461),
.B(n_9502),
.Y(n_11960)
);

INVx1_ASAP7_75t_L g11961 ( 
.A(n_10503),
.Y(n_11961)
);

AOI22xp5_ASAP7_75t_L g11962 ( 
.A1(n_11497),
.A2(n_10170),
.B1(n_10192),
.B2(n_10166),
.Y(n_11962)
);

BUFx2_ASAP7_75t_L g11963 ( 
.A(n_10474),
.Y(n_11963)
);

INVxp67_ASAP7_75t_SL g11964 ( 
.A(n_11518),
.Y(n_11964)
);

AOI22xp33_ASAP7_75t_L g11965 ( 
.A1(n_10861),
.A2(n_10883),
.B1(n_11024),
.B2(n_10864),
.Y(n_11965)
);

OAI22xp5_ASAP7_75t_L g11966 ( 
.A1(n_10497),
.A2(n_9365),
.B1(n_9469),
.B2(n_9335),
.Y(n_11966)
);

OAI22xp33_ASAP7_75t_SL g11967 ( 
.A1(n_11193),
.A2(n_10211),
.B1(n_10222),
.B2(n_10192),
.Y(n_11967)
);

NAND2xp5_ASAP7_75t_L g11968 ( 
.A(n_10792),
.B(n_10350),
.Y(n_11968)
);

AOI221xp5_ASAP7_75t_L g11969 ( 
.A1(n_10592),
.A2(n_8706),
.B1(n_8840),
.B2(n_8610),
.C(n_8516),
.Y(n_11969)
);

OAI211xp5_ASAP7_75t_L g11970 ( 
.A1(n_10592),
.A2(n_7832),
.B(n_7747),
.C(n_7841),
.Y(n_11970)
);

OAI22xp33_ASAP7_75t_L g11971 ( 
.A1(n_11369),
.A2(n_10190),
.B1(n_10117),
.B2(n_9660),
.Y(n_11971)
);

OAI21x1_ASAP7_75t_L g11972 ( 
.A1(n_10509),
.A2(n_9554),
.B(n_9277),
.Y(n_11972)
);

BUFx2_ASAP7_75t_L g11973 ( 
.A(n_10497),
.Y(n_11973)
);

BUFx3_ASAP7_75t_L g11974 ( 
.A(n_10560),
.Y(n_11974)
);

A2O1A1Ixp33_ASAP7_75t_L g11975 ( 
.A1(n_10560),
.A2(n_9891),
.B(n_8645),
.C(n_8476),
.Y(n_11975)
);

OAI22xp5_ASAP7_75t_L g11976 ( 
.A1(n_10600),
.A2(n_9602),
.B1(n_9637),
.B2(n_9501),
.Y(n_11976)
);

AND2x4_ASAP7_75t_L g11977 ( 
.A(n_11511),
.B(n_9501),
.Y(n_11977)
);

AOI221xp5_ASAP7_75t_L g11978 ( 
.A1(n_10694),
.A2(n_8840),
.B1(n_8610),
.B2(n_8516),
.C(n_8473),
.Y(n_11978)
);

AOI221xp5_ASAP7_75t_L g11979 ( 
.A1(n_10694),
.A2(n_8533),
.B1(n_7923),
.B2(n_8966),
.C(n_8617),
.Y(n_11979)
);

INVx3_ASAP7_75t_L g11980 ( 
.A(n_11120),
.Y(n_11980)
);

INVx1_ASAP7_75t_L g11981 ( 
.A(n_10506),
.Y(n_11981)
);

OAI211xp5_ASAP7_75t_SL g11982 ( 
.A1(n_10656),
.A2(n_9860),
.B(n_10194),
.C(n_10162),
.Y(n_11982)
);

OAI22xp5_ASAP7_75t_L g11983 ( 
.A1(n_10600),
.A2(n_9602),
.B1(n_9637),
.B2(n_9501),
.Y(n_11983)
);

OAI22xp5_ASAP7_75t_L g11984 ( 
.A1(n_10634),
.A2(n_9637),
.B1(n_9602),
.B2(n_10117),
.Y(n_11984)
);

AOI22xp33_ASAP7_75t_L g11985 ( 
.A1(n_10864),
.A2(n_9797),
.B1(n_9816),
.B2(n_9779),
.Y(n_11985)
);

AOI22xp33_ASAP7_75t_L g11986 ( 
.A1(n_10864),
.A2(n_9851),
.B1(n_9902),
.B2(n_9816),
.Y(n_11986)
);

AOI22xp33_ASAP7_75t_L g11987 ( 
.A1(n_10864),
.A2(n_9902),
.B1(n_9851),
.B2(n_9660),
.Y(n_11987)
);

AND2x2_ASAP7_75t_L g11988 ( 
.A(n_10468),
.B(n_10211),
.Y(n_11988)
);

AOI22xp33_ASAP7_75t_L g11989 ( 
.A1(n_10883),
.A2(n_9902),
.B1(n_9851),
.B2(n_9660),
.Y(n_11989)
);

BUFx3_ASAP7_75t_L g11990 ( 
.A(n_10634),
.Y(n_11990)
);

AOI22xp33_ASAP7_75t_L g11991 ( 
.A1(n_10883),
.A2(n_9660),
.B1(n_9813),
.B2(n_9801),
.Y(n_11991)
);

INVx1_ASAP7_75t_L g11992 ( 
.A(n_10510),
.Y(n_11992)
);

AOI22xp33_ASAP7_75t_L g11993 ( 
.A1(n_10883),
.A2(n_9801),
.B1(n_9903),
.B2(n_9813),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_10514),
.Y(n_11994)
);

AOI22xp33_ASAP7_75t_SL g11995 ( 
.A1(n_10888),
.A2(n_10403),
.B1(n_10565),
.B2(n_10441),
.Y(n_11995)
);

BUFx2_ASAP7_75t_L g11996 ( 
.A(n_10635),
.Y(n_11996)
);

AOI21xp33_ASAP7_75t_L g11997 ( 
.A1(n_11369),
.A2(n_10222),
.B(n_7751),
.Y(n_11997)
);

INVx1_ASAP7_75t_SL g11998 ( 
.A(n_11358),
.Y(n_11998)
);

AND2x2_ASAP7_75t_L g11999 ( 
.A(n_10496),
.B(n_9038),
.Y(n_11999)
);

INVx1_ASAP7_75t_L g12000 ( 
.A(n_10519),
.Y(n_12000)
);

AOI22xp33_ASAP7_75t_SL g12001 ( 
.A1(n_10441),
.A2(n_7957),
.B1(n_7841),
.B2(n_8488),
.Y(n_12001)
);

OAI221xp5_ASAP7_75t_L g12002 ( 
.A1(n_11369),
.A2(n_9637),
.B1(n_9602),
.B2(n_10317),
.C(n_9160),
.Y(n_12002)
);

AND2x2_ASAP7_75t_L g12003 ( 
.A(n_10496),
.B(n_9038),
.Y(n_12003)
);

BUFx6f_ASAP7_75t_L g12004 ( 
.A(n_11024),
.Y(n_12004)
);

OR2x2_ASAP7_75t_L g12005 ( 
.A(n_10429),
.B(n_9505),
.Y(n_12005)
);

AOI22xp33_ASAP7_75t_L g12006 ( 
.A1(n_11024),
.A2(n_9801),
.B1(n_9903),
.B2(n_9813),
.Y(n_12006)
);

OR2x2_ASAP7_75t_L g12007 ( 
.A(n_11082),
.B(n_9549),
.Y(n_12007)
);

AOI22xp33_ASAP7_75t_L g12008 ( 
.A1(n_11024),
.A2(n_11318),
.B1(n_11434),
.B2(n_11036),
.Y(n_12008)
);

OAI221xp5_ASAP7_75t_L g12009 ( 
.A1(n_11369),
.A2(n_9160),
.B1(n_8447),
.B2(n_8736),
.C(n_8181),
.Y(n_12009)
);

OAI22xp33_ASAP7_75t_L g12010 ( 
.A1(n_11242),
.A2(n_10190),
.B1(n_10117),
.B2(n_9801),
.Y(n_12010)
);

AOI222xp33_ASAP7_75t_L g12011 ( 
.A1(n_10635),
.A2(n_8517),
.B1(n_8921),
.B2(n_8499),
.C1(n_8485),
.C2(n_8707),
.Y(n_12011)
);

AOI22xp5_ASAP7_75t_SL g12012 ( 
.A1(n_10652),
.A2(n_9282),
.B1(n_9353),
.B2(n_9343),
.Y(n_12012)
);

INVx3_ASAP7_75t_L g12013 ( 
.A(n_11120),
.Y(n_12013)
);

NAND4xp25_ASAP7_75t_L g12014 ( 
.A(n_10652),
.B(n_8181),
.C(n_8471),
.D(n_8225),
.Y(n_12014)
);

OR2x2_ASAP7_75t_L g12015 ( 
.A(n_11082),
.B(n_9549),
.Y(n_12015)
);

OAI22xp33_ASAP7_75t_L g12016 ( 
.A1(n_11193),
.A2(n_10190),
.B1(n_11321),
.B2(n_9813),
.Y(n_12016)
);

AOI22xp33_ASAP7_75t_L g12017 ( 
.A1(n_11036),
.A2(n_9903),
.B1(n_8225),
.B2(n_10005),
.Y(n_12017)
);

AOI21xp5_ASAP7_75t_L g12018 ( 
.A1(n_11030),
.A2(n_8035),
.B(n_8690),
.Y(n_12018)
);

CKINVDCx11_ASAP7_75t_R g12019 ( 
.A(n_10655),
.Y(n_12019)
);

NAND2xp5_ASAP7_75t_SL g12020 ( 
.A(n_11511),
.B(n_9678),
.Y(n_12020)
);

OAI211xp5_ASAP7_75t_L g12021 ( 
.A1(n_10694),
.A2(n_7841),
.B(n_7751),
.C(n_9926),
.Y(n_12021)
);

AOI22xp33_ASAP7_75t_L g12022 ( 
.A1(n_11036),
.A2(n_9903),
.B1(n_10263),
.B2(n_9028),
.Y(n_12022)
);

OAI221xp5_ASAP7_75t_L g12023 ( 
.A1(n_10840),
.A2(n_8736),
.B1(n_8707),
.B2(n_7960),
.C(n_8074),
.Y(n_12023)
);

INVx4_ASAP7_75t_L g12024 ( 
.A(n_10398),
.Y(n_12024)
);

INVx3_ASAP7_75t_L g12025 ( 
.A(n_11484),
.Y(n_12025)
);

AOI22xp33_ASAP7_75t_SL g12026 ( 
.A1(n_10438),
.A2(n_7841),
.B1(n_8506),
.B2(n_8488),
.Y(n_12026)
);

AOI22xp33_ASAP7_75t_SL g12027 ( 
.A1(n_10438),
.A2(n_8488),
.B1(n_8506),
.B2(n_8787),
.Y(n_12027)
);

INVx1_ASAP7_75t_L g12028 ( 
.A(n_10525),
.Y(n_12028)
);

O2A1O1Ixp33_ASAP7_75t_SL g12029 ( 
.A1(n_10449),
.A2(n_10511),
.B(n_10529),
.C(n_10492),
.Y(n_12029)
);

AOI32xp33_ASAP7_75t_L g12030 ( 
.A1(n_10840),
.A2(n_8063),
.A3(n_7979),
.B1(n_8471),
.B2(n_7920),
.Y(n_12030)
);

AOI22xp33_ASAP7_75t_L g12031 ( 
.A1(n_11036),
.A2(n_9028),
.B1(n_10372),
.B2(n_9777),
.Y(n_12031)
);

INVx1_ASAP7_75t_L g12032 ( 
.A(n_10527),
.Y(n_12032)
);

AOI221xp5_ASAP7_75t_L g12033 ( 
.A1(n_10840),
.A2(n_8966),
.B1(n_8212),
.B2(n_9445),
.C(n_8690),
.Y(n_12033)
);

OAI211xp5_ASAP7_75t_SL g12034 ( 
.A1(n_10656),
.A2(n_9165),
.B(n_9363),
.C(n_9278),
.Y(n_12034)
);

AOI22xp33_ASAP7_75t_SL g12035 ( 
.A1(n_10442),
.A2(n_8488),
.B1(n_8506),
.B2(n_8787),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_10533),
.Y(n_12036)
);

AOI22xp33_ASAP7_75t_SL g12037 ( 
.A1(n_10442),
.A2(n_8488),
.B1(n_8506),
.B2(n_8787),
.Y(n_12037)
);

OAI22xp5_ASAP7_75t_L g12038 ( 
.A1(n_10655),
.A2(n_10190),
.B1(n_10372),
.B2(n_8105),
.Y(n_12038)
);

AOI22xp33_ASAP7_75t_L g12039 ( 
.A1(n_11318),
.A2(n_9777),
.B1(n_9679),
.B2(n_8441),
.Y(n_12039)
);

OAI22xp33_ASAP7_75t_L g12040 ( 
.A1(n_11321),
.A2(n_8645),
.B1(n_8354),
.B2(n_8400),
.Y(n_12040)
);

AOI22xp33_ASAP7_75t_L g12041 ( 
.A1(n_11318),
.A2(n_9777),
.B1(n_9679),
.B2(n_8441),
.Y(n_12041)
);

INVx1_ASAP7_75t_L g12042 ( 
.A(n_10535),
.Y(n_12042)
);

OAI221xp5_ASAP7_75t_L g12043 ( 
.A1(n_11104),
.A2(n_7866),
.B1(n_8074),
.B2(n_7960),
.C(n_7820),
.Y(n_12043)
);

AOI221xp5_ASAP7_75t_L g12044 ( 
.A1(n_11104),
.A2(n_9445),
.B1(n_9425),
.B2(n_8499),
.C(n_8433),
.Y(n_12044)
);

OAI22xp33_ASAP7_75t_L g12045 ( 
.A1(n_11163),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12045)
);

AOI22xp33_ASAP7_75t_SL g12046 ( 
.A1(n_11531),
.A2(n_8488),
.B1(n_8506),
.B2(n_8787),
.Y(n_12046)
);

AOI22xp5_ASAP7_75t_L g12047 ( 
.A1(n_11531),
.A2(n_11114),
.B1(n_11144),
.B2(n_11104),
.Y(n_12047)
);

INVx2_ASAP7_75t_L g12048 ( 
.A(n_10486),
.Y(n_12048)
);

OAI221xp5_ASAP7_75t_L g12049 ( 
.A1(n_11114),
.A2(n_7866),
.B1(n_8179),
.B2(n_7820),
.C(n_8921),
.Y(n_12049)
);

OR2x2_ASAP7_75t_L g12050 ( 
.A(n_10771),
.B(n_10350),
.Y(n_12050)
);

INVx1_ASAP7_75t_L g12051 ( 
.A(n_10537),
.Y(n_12051)
);

INVx1_ASAP7_75t_L g12052 ( 
.A(n_10551),
.Y(n_12052)
);

BUFx6f_ASAP7_75t_L g12053 ( 
.A(n_11318),
.Y(n_12053)
);

AOI22xp33_ASAP7_75t_L g12054 ( 
.A1(n_11434),
.A2(n_11479),
.B1(n_10716),
.B2(n_10745),
.Y(n_12054)
);

INVx1_ASAP7_75t_L g12055 ( 
.A(n_10553),
.Y(n_12055)
);

OAI221xp5_ASAP7_75t_L g12056 ( 
.A1(n_11114),
.A2(n_8179),
.B1(n_10361),
.B2(n_10354),
.C(n_9713),
.Y(n_12056)
);

BUFx2_ASAP7_75t_L g12057 ( 
.A(n_10661),
.Y(n_12057)
);

AO31x2_ASAP7_75t_L g12058 ( 
.A1(n_11144),
.A2(n_9411),
.A3(n_9412),
.B(n_9401),
.Y(n_12058)
);

AOI22xp33_ASAP7_75t_L g12059 ( 
.A1(n_11434),
.A2(n_9777),
.B1(n_9679),
.B2(n_8441),
.Y(n_12059)
);

NAND4xp25_ASAP7_75t_SL g12060 ( 
.A(n_10411),
.B(n_8622),
.C(n_8296),
.D(n_8428),
.Y(n_12060)
);

CKINVDCx5p33_ASAP7_75t_R g12061 ( 
.A(n_11358),
.Y(n_12061)
);

OAI22xp33_ASAP7_75t_L g12062 ( 
.A1(n_11163),
.A2(n_11179),
.B1(n_11336),
.B2(n_11211),
.Y(n_12062)
);

AOI22xp33_ASAP7_75t_L g12063 ( 
.A1(n_11434),
.A2(n_9777),
.B1(n_9679),
.B2(n_8441),
.Y(n_12063)
);

NAND2xp5_ASAP7_75t_L g12064 ( 
.A(n_10797),
.B(n_8251),
.Y(n_12064)
);

INVxp67_ASAP7_75t_L g12065 ( 
.A(n_10661),
.Y(n_12065)
);

INVx1_ASAP7_75t_SL g12066 ( 
.A(n_11453),
.Y(n_12066)
);

AOI22xp33_ASAP7_75t_L g12067 ( 
.A1(n_11479),
.A2(n_9679),
.B1(n_8441),
.B2(n_8752),
.Y(n_12067)
);

INVx2_ASAP7_75t_L g12068 ( 
.A(n_10486),
.Y(n_12068)
);

AOI221xp5_ASAP7_75t_L g12069 ( 
.A1(n_11144),
.A2(n_9445),
.B1(n_9425),
.B2(n_8433),
.C(n_8365),
.Y(n_12069)
);

AOI21xp5_ASAP7_75t_L g12070 ( 
.A1(n_11030),
.A2(n_8163),
.B(n_9276),
.Y(n_12070)
);

OAI22xp33_ASAP7_75t_L g12071 ( 
.A1(n_11179),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12071)
);

INVx4_ASAP7_75t_L g12072 ( 
.A(n_10398),
.Y(n_12072)
);

AOI22xp33_ASAP7_75t_L g12073 ( 
.A1(n_11479),
.A2(n_8441),
.B1(n_8752),
.B2(n_8565),
.Y(n_12073)
);

AOI22xp33_ASAP7_75t_L g12074 ( 
.A1(n_11479),
.A2(n_10745),
.B1(n_10809),
.B2(n_10716),
.Y(n_12074)
);

AND2x4_ASAP7_75t_L g12075 ( 
.A(n_11393),
.B(n_9933),
.Y(n_12075)
);

OAI22xp33_ASAP7_75t_L g12076 ( 
.A1(n_11211),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12076)
);

OAI22xp5_ASAP7_75t_L g12077 ( 
.A1(n_10809),
.A2(n_8105),
.B1(n_9359),
.B2(n_8969),
.Y(n_12077)
);

AND2x2_ASAP7_75t_L g12078 ( 
.A(n_10902),
.B(n_10964),
.Y(n_12078)
);

AOI22xp33_ASAP7_75t_L g12079 ( 
.A1(n_10885),
.A2(n_8441),
.B1(n_8752),
.B2(n_8565),
.Y(n_12079)
);

NAND2xp5_ASAP7_75t_L g12080 ( 
.A(n_10798),
.B(n_8251),
.Y(n_12080)
);

OR2x2_ASAP7_75t_L g12081 ( 
.A(n_10771),
.B(n_8872),
.Y(n_12081)
);

OAI22xp5_ASAP7_75t_L g12082 ( 
.A1(n_10885),
.A2(n_9359),
.B1(n_8969),
.B2(n_9029),
.Y(n_12082)
);

INVx2_ASAP7_75t_L g12083 ( 
.A(n_10495),
.Y(n_12083)
);

INVx2_ASAP7_75t_L g12084 ( 
.A(n_10495),
.Y(n_12084)
);

HB1xp67_ASAP7_75t_L g12085 ( 
.A(n_10815),
.Y(n_12085)
);

AOI22xp33_ASAP7_75t_L g12086 ( 
.A1(n_10917),
.A2(n_8565),
.B1(n_8753),
.B2(n_8752),
.Y(n_12086)
);

AOI22xp33_ASAP7_75t_L g12087 ( 
.A1(n_10917),
.A2(n_8565),
.B1(n_8753),
.B2(n_8752),
.Y(n_12087)
);

AOI22xp33_ASAP7_75t_L g12088 ( 
.A1(n_10955),
.A2(n_8565),
.B1(n_8753),
.B2(n_8752),
.Y(n_12088)
);

INVx3_ASAP7_75t_L g12089 ( 
.A(n_11484),
.Y(n_12089)
);

OAI221xp5_ASAP7_75t_L g12090 ( 
.A1(n_11203),
.A2(n_10361),
.B1(n_10354),
.B2(n_8741),
.C(n_8838),
.Y(n_12090)
);

AOI22xp33_ASAP7_75t_L g12091 ( 
.A1(n_10955),
.A2(n_8565),
.B1(n_8753),
.B2(n_8752),
.Y(n_12091)
);

AO21x2_ASAP7_75t_L g12092 ( 
.A1(n_10385),
.A2(n_9412),
.B(n_9411),
.Y(n_12092)
);

NAND2xp5_ASAP7_75t_L g12093 ( 
.A(n_10824),
.B(n_10829),
.Y(n_12093)
);

AND2x4_ASAP7_75t_L g12094 ( 
.A(n_10648),
.B(n_9933),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_10561),
.Y(n_12095)
);

AND2x2_ASAP7_75t_L g12096 ( 
.A(n_10902),
.B(n_10964),
.Y(n_12096)
);

BUFx4f_ASAP7_75t_L g12097 ( 
.A(n_11030),
.Y(n_12097)
);

BUFx4f_ASAP7_75t_L g12098 ( 
.A(n_10805),
.Y(n_12098)
);

OA21x2_ASAP7_75t_L g12099 ( 
.A1(n_10437),
.A2(n_9427),
.B(n_9412),
.Y(n_12099)
);

OAI21x1_ASAP7_75t_L g12100 ( 
.A1(n_10484),
.A2(n_11072),
.B(n_10477),
.Y(n_12100)
);

NOR2xp33_ASAP7_75t_L g12101 ( 
.A(n_10960),
.B(n_9767),
.Y(n_12101)
);

AOI21xp5_ASAP7_75t_L g12102 ( 
.A1(n_10960),
.A2(n_8553),
.B(n_9361),
.Y(n_12102)
);

OAI22xp33_ASAP7_75t_L g12103 ( 
.A1(n_11336),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12103)
);

AOI22xp33_ASAP7_75t_L g12104 ( 
.A1(n_10981),
.A2(n_8565),
.B1(n_8753),
.B2(n_8622),
.Y(n_12104)
);

INVx3_ASAP7_75t_L g12105 ( 
.A(n_11484),
.Y(n_12105)
);

OAI22xp33_ASAP7_75t_L g12106 ( 
.A1(n_10805),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12106)
);

AOI22xp33_ASAP7_75t_L g12107 ( 
.A1(n_10981),
.A2(n_8753),
.B1(n_8296),
.B2(n_8598),
.Y(n_12107)
);

NOR2xp33_ASAP7_75t_L g12108 ( 
.A(n_10985),
.B(n_9105),
.Y(n_12108)
);

AOI22xp33_ASAP7_75t_L g12109 ( 
.A1(n_10985),
.A2(n_11389),
.B1(n_11203),
.B2(n_11490),
.Y(n_12109)
);

AOI22xp33_ASAP7_75t_L g12110 ( 
.A1(n_11203),
.A2(n_11389),
.B1(n_11490),
.B2(n_10805),
.Y(n_12110)
);

AOI22xp33_ASAP7_75t_L g12111 ( 
.A1(n_11389),
.A2(n_8753),
.B1(n_8598),
.B2(n_8587),
.Y(n_12111)
);

OAI22xp5_ASAP7_75t_L g12112 ( 
.A1(n_11257),
.A2(n_9029),
.B1(n_7921),
.B2(n_7766),
.Y(n_12112)
);

CKINVDCx5p33_ASAP7_75t_R g12113 ( 
.A(n_11453),
.Y(n_12113)
);

AOI22xp5_ASAP7_75t_L g12114 ( 
.A1(n_10791),
.A2(n_8994),
.B1(n_8833),
.B2(n_9163),
.Y(n_12114)
);

CKINVDCx5p33_ASAP7_75t_R g12115 ( 
.A(n_11456),
.Y(n_12115)
);

AND2x4_ASAP7_75t_L g12116 ( 
.A(n_10648),
.B(n_10806),
.Y(n_12116)
);

INVx1_ASAP7_75t_L g12117 ( 
.A(n_10568),
.Y(n_12117)
);

OAI221xp5_ASAP7_75t_L g12118 ( 
.A1(n_10805),
.A2(n_8827),
.B1(n_8838),
.B2(n_8741),
.C(n_8934),
.Y(n_12118)
);

AOI221xp5_ASAP7_75t_L g12119 ( 
.A1(n_10845),
.A2(n_9445),
.B1(n_9425),
.B2(n_8365),
.C(n_8378),
.Y(n_12119)
);

BUFx12f_ASAP7_75t_L g12120 ( 
.A(n_11456),
.Y(n_12120)
);

OAI211xp5_ASAP7_75t_SL g12121 ( 
.A1(n_10495),
.A2(n_9278),
.B(n_9363),
.C(n_9165),
.Y(n_12121)
);

AND2x6_ASAP7_75t_L g12122 ( 
.A(n_11257),
.B(n_9526),
.Y(n_12122)
);

AOI221xp5_ASAP7_75t_L g12123 ( 
.A1(n_10846),
.A2(n_9425),
.B1(n_8378),
.B2(n_8322),
.C(n_8302),
.Y(n_12123)
);

HB1xp67_ASAP7_75t_L g12124 ( 
.A(n_10847),
.Y(n_12124)
);

INVx2_ASAP7_75t_L g12125 ( 
.A(n_10534),
.Y(n_12125)
);

AOI22xp33_ASAP7_75t_L g12126 ( 
.A1(n_10872),
.A2(n_8598),
.B1(n_8587),
.B2(n_10370),
.Y(n_12126)
);

AOI22xp33_ASAP7_75t_L g12127 ( 
.A1(n_10872),
.A2(n_8587),
.B1(n_10370),
.B2(n_9174),
.Y(n_12127)
);

BUFx2_ASAP7_75t_R g12128 ( 
.A(n_10459),
.Y(n_12128)
);

INVx2_ASAP7_75t_L g12129 ( 
.A(n_10534),
.Y(n_12129)
);

AND2x2_ASAP7_75t_L g12130 ( 
.A(n_10902),
.B(n_9642),
.Y(n_12130)
);

OAI22xp5_ASAP7_75t_L g12131 ( 
.A1(n_11257),
.A2(n_7921),
.B1(n_7766),
.B2(n_8934),
.Y(n_12131)
);

BUFx3_ASAP7_75t_L g12132 ( 
.A(n_10791),
.Y(n_12132)
);

INVx1_ASAP7_75t_L g12133 ( 
.A(n_10571),
.Y(n_12133)
);

OAI222xp33_ASAP7_75t_L g12134 ( 
.A1(n_10872),
.A2(n_8399),
.B1(n_8208),
.B2(n_8160),
.C1(n_8962),
.C2(n_8959),
.Y(n_12134)
);

OAI22xp33_ASAP7_75t_L g12135 ( 
.A1(n_10872),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12135)
);

OAI22xp5_ASAP7_75t_L g12136 ( 
.A1(n_10964),
.A2(n_7921),
.B1(n_7766),
.B2(n_9389),
.Y(n_12136)
);

OAI21x1_ASAP7_75t_L g12137 ( 
.A1(n_10484),
.A2(n_9278),
.B(n_9165),
.Y(n_12137)
);

INVx2_ASAP7_75t_L g12138 ( 
.A(n_10534),
.Y(n_12138)
);

AND2x4_ASAP7_75t_L g12139 ( 
.A(n_10648),
.B(n_9933),
.Y(n_12139)
);

OAI22xp33_ASAP7_75t_L g12140 ( 
.A1(n_10849),
.A2(n_8354),
.B1(n_8400),
.B2(n_7948),
.Y(n_12140)
);

AOI22xp33_ASAP7_75t_L g12141 ( 
.A1(n_11023),
.A2(n_10370),
.B1(n_9174),
.B2(n_9198),
.Y(n_12141)
);

OAI22xp33_ASAP7_75t_L g12142 ( 
.A1(n_10880),
.A2(n_8593),
.B1(n_7948),
.B2(n_7921),
.Y(n_12142)
);

AND2x2_ASAP7_75t_L g12143 ( 
.A(n_11023),
.B(n_9642),
.Y(n_12143)
);

NAND2xp5_ASAP7_75t_L g12144 ( 
.A(n_10881),
.B(n_8302),
.Y(n_12144)
);

AOI221xp5_ASAP7_75t_L g12145 ( 
.A1(n_10892),
.A2(n_8322),
.B1(n_8398),
.B2(n_8485),
.C(n_9345),
.Y(n_12145)
);

AOI22xp33_ASAP7_75t_L g12146 ( 
.A1(n_11023),
.A2(n_10370),
.B1(n_9174),
.B2(n_9198),
.Y(n_12146)
);

AND2x2_ASAP7_75t_L g12147 ( 
.A(n_11138),
.B(n_9646),
.Y(n_12147)
);

AOI22xp33_ASAP7_75t_L g12148 ( 
.A1(n_11138),
.A2(n_9174),
.B1(n_9198),
.B2(n_9163),
.Y(n_12148)
);

OAI22xp5_ASAP7_75t_L g12149 ( 
.A1(n_11138),
.A2(n_9392),
.B1(n_9430),
.B2(n_9393),
.Y(n_12149)
);

AOI22xp33_ASAP7_75t_L g12150 ( 
.A1(n_11259),
.A2(n_10791),
.B1(n_10620),
.B2(n_10657),
.Y(n_12150)
);

AND2x2_ASAP7_75t_L g12151 ( 
.A(n_11259),
.B(n_9646),
.Y(n_12151)
);

AOI22xp33_ASAP7_75t_L g12152 ( 
.A1(n_11259),
.A2(n_9198),
.B1(n_9219),
.B2(n_9163),
.Y(n_12152)
);

AOI21xp5_ASAP7_75t_L g12153 ( 
.A1(n_11247),
.A2(n_8553),
.B(n_9474),
.Y(n_12153)
);

AND2x2_ASAP7_75t_L g12154 ( 
.A(n_10547),
.B(n_10620),
.Y(n_12154)
);

INVx1_ASAP7_75t_L g12155 ( 
.A(n_10572),
.Y(n_12155)
);

OR2x6_ASAP7_75t_L g12156 ( 
.A(n_11437),
.B(n_7396),
.Y(n_12156)
);

OAI22xp5_ASAP7_75t_L g12157 ( 
.A1(n_10411),
.A2(n_9537),
.B1(n_9634),
.B2(n_9621),
.Y(n_12157)
);

AOI221xp5_ASAP7_75t_L g12158 ( 
.A1(n_10893),
.A2(n_8398),
.B1(n_9345),
.B2(n_9352),
.C(n_8527),
.Y(n_12158)
);

INVx1_ASAP7_75t_L g12159 ( 
.A(n_10573),
.Y(n_12159)
);

INVx1_ASAP7_75t_L g12160 ( 
.A(n_10576),
.Y(n_12160)
);

AOI22xp33_ASAP7_75t_L g12161 ( 
.A1(n_10791),
.A2(n_9219),
.B1(n_9297),
.B2(n_9163),
.Y(n_12161)
);

AOI22xp33_ASAP7_75t_L g12162 ( 
.A1(n_10791),
.A2(n_9297),
.B1(n_9362),
.B2(n_9219),
.Y(n_12162)
);

OAI22xp33_ASAP7_75t_L g12163 ( 
.A1(n_10942),
.A2(n_8593),
.B1(n_10953),
.B2(n_10947),
.Y(n_12163)
);

INVx1_ASAP7_75t_SL g12164 ( 
.A(n_10806),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_10577),
.Y(n_12165)
);

AOI22xp33_ASAP7_75t_L g12166 ( 
.A1(n_10547),
.A2(n_10620),
.B1(n_10660),
.B2(n_10657),
.Y(n_12166)
);

OAI22xp5_ASAP7_75t_L g12167 ( 
.A1(n_10434),
.A2(n_9703),
.B1(n_9774),
.B2(n_9714),
.Y(n_12167)
);

NAND3xp33_ASAP7_75t_L g12168 ( 
.A(n_11154),
.B(n_7751),
.C(n_8787),
.Y(n_12168)
);

OAI21xp5_ASAP7_75t_L g12169 ( 
.A1(n_10450),
.A2(n_7914),
.B(n_8025),
.Y(n_12169)
);

OAI22xp33_ASAP7_75t_L g12170 ( 
.A1(n_10954),
.A2(n_8593),
.B1(n_8018),
.B2(n_8119),
.Y(n_12170)
);

AOI22xp33_ASAP7_75t_L g12171 ( 
.A1(n_10547),
.A2(n_9297),
.B1(n_9362),
.B2(n_9219),
.Y(n_12171)
);

AOI22xp5_ASAP7_75t_L g12172 ( 
.A1(n_10657),
.A2(n_8994),
.B1(n_8833),
.B2(n_9297),
.Y(n_12172)
);

AND2x2_ASAP7_75t_L g12173 ( 
.A(n_10660),
.B(n_9671),
.Y(n_12173)
);

AND2x4_ASAP7_75t_L g12174 ( 
.A(n_10806),
.B(n_9933),
.Y(n_12174)
);

AND2x2_ASAP7_75t_L g12175 ( 
.A(n_10660),
.B(n_10671),
.Y(n_12175)
);

AOI22xp33_ASAP7_75t_L g12176 ( 
.A1(n_10671),
.A2(n_9590),
.B1(n_9625),
.B2(n_9362),
.Y(n_12176)
);

AOI221xp5_ASAP7_75t_L g12177 ( 
.A1(n_10993),
.A2(n_9352),
.B1(n_9345),
.B2(n_8527),
.C(n_8868),
.Y(n_12177)
);

AOI22xp33_ASAP7_75t_L g12178 ( 
.A1(n_10671),
.A2(n_9590),
.B1(n_9625),
.B2(n_9362),
.Y(n_12178)
);

AOI22xp33_ASAP7_75t_L g12179 ( 
.A1(n_10672),
.A2(n_9625),
.B1(n_9863),
.B2(n_9590),
.Y(n_12179)
);

AOI22xp33_ASAP7_75t_SL g12180 ( 
.A1(n_10434),
.A2(n_8506),
.B1(n_8817),
.B2(n_8813),
.Y(n_12180)
);

BUFx4f_ASAP7_75t_SL g12181 ( 
.A(n_10672),
.Y(n_12181)
);

INVx1_ASAP7_75t_L g12182 ( 
.A(n_10578),
.Y(n_12182)
);

AOI22xp33_ASAP7_75t_L g12183 ( 
.A1(n_10672),
.A2(n_9625),
.B1(n_9863),
.B2(n_9590),
.Y(n_12183)
);

AOI22xp33_ASAP7_75t_L g12184 ( 
.A1(n_10742),
.A2(n_9895),
.B1(n_9897),
.B2(n_9863),
.Y(n_12184)
);

OAI21xp5_ASAP7_75t_SL g12185 ( 
.A1(n_11370),
.A2(n_8370),
.B(n_8827),
.Y(n_12185)
);

AND2x2_ASAP7_75t_L g12186 ( 
.A(n_10742),
.B(n_9671),
.Y(n_12186)
);

INVx1_ASAP7_75t_L g12187 ( 
.A(n_10579),
.Y(n_12187)
);

AOI22xp33_ASAP7_75t_L g12188 ( 
.A1(n_10742),
.A2(n_9895),
.B1(n_9897),
.B2(n_9863),
.Y(n_12188)
);

INVx1_ASAP7_75t_L g12189 ( 
.A(n_10582),
.Y(n_12189)
);

AOI22xp33_ASAP7_75t_L g12190 ( 
.A1(n_10879),
.A2(n_9897),
.B1(n_9895),
.B2(n_8046),
.Y(n_12190)
);

BUFx3_ASAP7_75t_L g12191 ( 
.A(n_10879),
.Y(n_12191)
);

INVx1_ASAP7_75t_L g12192 ( 
.A(n_10584),
.Y(n_12192)
);

OAI22xp5_ASAP7_75t_L g12193 ( 
.A1(n_11075),
.A2(n_9873),
.B1(n_8593),
.B2(n_8046),
.Y(n_12193)
);

OAI221xp5_ASAP7_75t_L g12194 ( 
.A1(n_10780),
.A2(n_9363),
.B1(n_9378),
.B2(n_9278),
.C(n_9165),
.Y(n_12194)
);

INVx1_ASAP7_75t_L g12195 ( 
.A(n_10588),
.Y(n_12195)
);

AOI22xp33_ASAP7_75t_L g12196 ( 
.A1(n_10879),
.A2(n_9897),
.B1(n_9895),
.B2(n_8046),
.Y(n_12196)
);

BUFx3_ASAP7_75t_L g12197 ( 
.A(n_10775),
.Y(n_12197)
);

CKINVDCx5p33_ASAP7_75t_R g12198 ( 
.A(n_11103),
.Y(n_12198)
);

INVx1_ASAP7_75t_L g12199 ( 
.A(n_10590),
.Y(n_12199)
);

AOI221xp5_ASAP7_75t_L g12200 ( 
.A1(n_11084),
.A2(n_9352),
.B1(n_9345),
.B2(n_8868),
.C(n_9985),
.Y(n_12200)
);

OAI221xp5_ASAP7_75t_L g12201 ( 
.A1(n_10780),
.A2(n_9438),
.B1(n_9472),
.B2(n_9378),
.C(n_9363),
.Y(n_12201)
);

AOI22xp33_ASAP7_75t_L g12202 ( 
.A1(n_11263),
.A2(n_8046),
.B1(n_8119),
.B2(n_8018),
.Y(n_12202)
);

OAI222xp33_ASAP7_75t_L g12203 ( 
.A1(n_11307),
.A2(n_8399),
.B1(n_8208),
.B2(n_8160),
.C1(n_8962),
.C2(n_8959),
.Y(n_12203)
);

AOI22xp33_ASAP7_75t_L g12204 ( 
.A1(n_11263),
.A2(n_8119),
.B1(n_8133),
.B2(n_8018),
.Y(n_12204)
);

AOI22xp33_ASAP7_75t_L g12205 ( 
.A1(n_11263),
.A2(n_8119),
.B1(n_8133),
.B2(n_8018),
.Y(n_12205)
);

NAND2xp5_ASAP7_75t_L g12206 ( 
.A(n_11113),
.B(n_9493),
.Y(n_12206)
);

BUFx3_ASAP7_75t_L g12207 ( 
.A(n_10775),
.Y(n_12207)
);

INVx1_ASAP7_75t_L g12208 ( 
.A(n_10591),
.Y(n_12208)
);

AOI22xp33_ASAP7_75t_L g12209 ( 
.A1(n_11350),
.A2(n_8189),
.B1(n_8197),
.B2(n_8133),
.Y(n_12209)
);

INVx1_ASAP7_75t_L g12210 ( 
.A(n_10597),
.Y(n_12210)
);

INVx1_ASAP7_75t_L g12211 ( 
.A(n_10603),
.Y(n_12211)
);

OAI22xp5_ASAP7_75t_L g12212 ( 
.A1(n_11124),
.A2(n_8593),
.B1(n_8189),
.B2(n_8197),
.Y(n_12212)
);

INVx1_ASAP7_75t_L g12213 ( 
.A(n_10605),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_10607),
.Y(n_12214)
);

OAI322xp33_ASAP7_75t_L g12215 ( 
.A1(n_10677),
.A2(n_9699),
.A3(n_9633),
.B1(n_10071),
.B2(n_10099),
.C1(n_9709),
.C2(n_9553),
.Y(n_12215)
);

AO31x2_ASAP7_75t_L g12216 ( 
.A1(n_10385),
.A2(n_9435),
.A3(n_9437),
.B(n_9427),
.Y(n_12216)
);

CKINVDCx5p33_ASAP7_75t_R g12217 ( 
.A(n_11103),
.Y(n_12217)
);

INVx11_ASAP7_75t_L g12218 ( 
.A(n_11103),
.Y(n_12218)
);

OAI22xp5_ASAP7_75t_L g12219 ( 
.A1(n_11150),
.A2(n_8593),
.B1(n_8189),
.B2(n_8197),
.Y(n_12219)
);

AOI221xp5_ASAP7_75t_L g12220 ( 
.A1(n_11153),
.A2(n_9352),
.B1(n_8868),
.B2(n_9985),
.C(n_7892),
.Y(n_12220)
);

AOI22xp5_ASAP7_75t_L g12221 ( 
.A1(n_11350),
.A2(n_9965),
.B1(n_10168),
.B2(n_10044),
.Y(n_12221)
);

INVx1_ASAP7_75t_L g12222 ( 
.A(n_10609),
.Y(n_12222)
);

OA21x2_ASAP7_75t_L g12223 ( 
.A1(n_10437),
.A2(n_9435),
.B(n_9427),
.Y(n_12223)
);

OA21x2_ASAP7_75t_L g12224 ( 
.A1(n_11072),
.A2(n_9437),
.B(n_9435),
.Y(n_12224)
);

OAI22xp5_ASAP7_75t_L g12225 ( 
.A1(n_11158),
.A2(n_8593),
.B1(n_8189),
.B2(n_8197),
.Y(n_12225)
);

BUFx8_ASAP7_75t_L g12226 ( 
.A(n_11237),
.Y(n_12226)
);

AOI222xp33_ASAP7_75t_L g12227 ( 
.A1(n_11165),
.A2(n_7848),
.B1(n_7920),
.B2(n_7954),
.C1(n_9633),
.C2(n_9553),
.Y(n_12227)
);

INVx2_ASAP7_75t_L g12228 ( 
.A(n_10536),
.Y(n_12228)
);

OAI22xp33_ASAP7_75t_SL g12229 ( 
.A1(n_10449),
.A2(n_9378),
.B1(n_9472),
.B2(n_9438),
.Y(n_12229)
);

OAI22xp5_ASAP7_75t_L g12230 ( 
.A1(n_11182),
.A2(n_8593),
.B1(n_8230),
.B2(n_8243),
.Y(n_12230)
);

AOI22xp33_ASAP7_75t_SL g12231 ( 
.A1(n_10596),
.A2(n_8817),
.B1(n_8813),
.B2(n_7914),
.Y(n_12231)
);

OAI22xp5_ASAP7_75t_L g12232 ( 
.A1(n_11195),
.A2(n_8230),
.B1(n_8243),
.B2(n_8133),
.Y(n_12232)
);

OR2x2_ASAP7_75t_L g12233 ( 
.A(n_10913),
.B(n_8872),
.Y(n_12233)
);

CKINVDCx11_ASAP7_75t_R g12234 ( 
.A(n_11237),
.Y(n_12234)
);

AOI221xp5_ASAP7_75t_SL g12235 ( 
.A1(n_11249),
.A2(n_8785),
.B1(n_8794),
.B2(n_9709),
.C(n_9699),
.Y(n_12235)
);

INVx11_ASAP7_75t_L g12236 ( 
.A(n_11237),
.Y(n_12236)
);

NOR2xp33_ASAP7_75t_L g12237 ( 
.A(n_11383),
.B(n_9487),
.Y(n_12237)
);

AOI322xp5_ASAP7_75t_L g12238 ( 
.A1(n_11310),
.A2(n_7920),
.A3(n_7954),
.B1(n_7848),
.B2(n_7826),
.C1(n_7765),
.C2(n_7752),
.Y(n_12238)
);

OAI21x1_ASAP7_75t_SL g12239 ( 
.A1(n_10492),
.A2(n_8918),
.B(n_8873),
.Y(n_12239)
);

BUFx6f_ASAP7_75t_L g12240 ( 
.A(n_10536),
.Y(n_12240)
);

OAI221xp5_ASAP7_75t_L g12241 ( 
.A1(n_11213),
.A2(n_9472),
.B1(n_9476),
.B2(n_9438),
.C(n_9378),
.Y(n_12241)
);

AOI211xp5_ASAP7_75t_L g12242 ( 
.A1(n_11370),
.A2(n_11375),
.B(n_11392),
.C(n_11391),
.Y(n_12242)
);

NAND2xp5_ASAP7_75t_L g12243 ( 
.A(n_11226),
.B(n_10071),
.Y(n_12243)
);

BUFx2_ASAP7_75t_L g12244 ( 
.A(n_11383),
.Y(n_12244)
);

AOI22xp33_ASAP7_75t_L g12245 ( 
.A1(n_11350),
.A2(n_8243),
.B1(n_8249),
.B2(n_8230),
.Y(n_12245)
);

AO21x2_ASAP7_75t_L g12246 ( 
.A1(n_10396),
.A2(n_9440),
.B(n_9437),
.Y(n_12246)
);

AOI22xp33_ASAP7_75t_L g12247 ( 
.A1(n_11421),
.A2(n_8243),
.B1(n_8249),
.B2(n_8230),
.Y(n_12247)
);

INVx1_ASAP7_75t_L g12248 ( 
.A(n_10618),
.Y(n_12248)
);

AOI221xp5_ASAP7_75t_L g12249 ( 
.A1(n_11228),
.A2(n_8868),
.B1(n_9985),
.B2(n_7892),
.C(n_8497),
.Y(n_12249)
);

AOI221xp5_ASAP7_75t_L g12250 ( 
.A1(n_11260),
.A2(n_8868),
.B1(n_9985),
.B2(n_7892),
.C(n_8497),
.Y(n_12250)
);

INVx2_ASAP7_75t_L g12251 ( 
.A(n_10536),
.Y(n_12251)
);

AOI22xp5_ASAP7_75t_L g12252 ( 
.A1(n_11421),
.A2(n_9965),
.B1(n_10168),
.B2(n_10044),
.Y(n_12252)
);

AOI22xp33_ASAP7_75t_L g12253 ( 
.A1(n_11421),
.A2(n_8424),
.B1(n_8442),
.B2(n_8249),
.Y(n_12253)
);

INVx4_ASAP7_75t_L g12254 ( 
.A(n_11383),
.Y(n_12254)
);

OA21x2_ASAP7_75t_L g12255 ( 
.A1(n_10396),
.A2(n_9441),
.B(n_9440),
.Y(n_12255)
);

AOI22xp33_ASAP7_75t_L g12256 ( 
.A1(n_11307),
.A2(n_8424),
.B1(n_8442),
.B2(n_8249),
.Y(n_12256)
);

AOI221xp5_ASAP7_75t_L g12257 ( 
.A1(n_11319),
.A2(n_7892),
.B1(n_8462),
.B2(n_8461),
.C(n_8261),
.Y(n_12257)
);

AND2x2_ASAP7_75t_L g12258 ( 
.A(n_10891),
.B(n_9688),
.Y(n_12258)
);

OAI21x1_ASAP7_75t_L g12259 ( 
.A1(n_10450),
.A2(n_10477),
.B(n_10735),
.Y(n_12259)
);

OAI22xp5_ASAP7_75t_L g12260 ( 
.A1(n_11337),
.A2(n_8424),
.B1(n_8580),
.B2(n_8442),
.Y(n_12260)
);

OAI221xp5_ASAP7_75t_L g12261 ( 
.A1(n_11338),
.A2(n_9476),
.B1(n_9612),
.B2(n_9472),
.C(n_9438),
.Y(n_12261)
);

AOI22xp33_ASAP7_75t_L g12262 ( 
.A1(n_11375),
.A2(n_8424),
.B1(n_8580),
.B2(n_8442),
.Y(n_12262)
);

AOI22xp33_ASAP7_75t_L g12263 ( 
.A1(n_11391),
.A2(n_8580),
.B1(n_8630),
.B2(n_8603),
.Y(n_12263)
);

OA21x2_ASAP7_75t_L g12264 ( 
.A1(n_10401),
.A2(n_9441),
.B(n_9440),
.Y(n_12264)
);

OAI21xp5_ASAP7_75t_L g12265 ( 
.A1(n_11368),
.A2(n_8025),
.B(n_7966),
.Y(n_12265)
);

AO21x2_ASAP7_75t_L g12266 ( 
.A1(n_10401),
.A2(n_9443),
.B(n_9441),
.Y(n_12266)
);

AO21x2_ASAP7_75t_L g12267 ( 
.A1(n_10406),
.A2(n_9511),
.B(n_9443),
.Y(n_12267)
);

BUFx6f_ASAP7_75t_L g12268 ( 
.A(n_10663),
.Y(n_12268)
);

AOI21xp33_ASAP7_75t_L g12269 ( 
.A1(n_11426),
.A2(n_7751),
.B(n_9526),
.Y(n_12269)
);

OAI221xp5_ASAP7_75t_L g12270 ( 
.A1(n_11420),
.A2(n_9630),
.B1(n_9804),
.B2(n_9612),
.C(n_9476),
.Y(n_12270)
);

OAI22xp5_ASAP7_75t_L g12271 ( 
.A1(n_11442),
.A2(n_8580),
.B1(n_8630),
.B2(n_8603),
.Y(n_12271)
);

OAI22xp5_ASAP7_75t_L g12272 ( 
.A1(n_10891),
.A2(n_8603),
.B1(n_8637),
.B2(n_8630),
.Y(n_12272)
);

OAI21x1_ASAP7_75t_L g12273 ( 
.A1(n_10735),
.A2(n_9612),
.B(n_9476),
.Y(n_12273)
);

INVx2_ASAP7_75t_L g12274 ( 
.A(n_10663),
.Y(n_12274)
);

AOI22xp33_ASAP7_75t_SL g12275 ( 
.A1(n_10596),
.A2(n_8813),
.B1(n_8817),
.B2(n_7751),
.Y(n_12275)
);

AND2x2_ASAP7_75t_L g12276 ( 
.A(n_10919),
.B(n_9688),
.Y(n_12276)
);

AOI22xp33_ASAP7_75t_SL g12277 ( 
.A1(n_10621),
.A2(n_8813),
.B1(n_8817),
.B2(n_7751),
.Y(n_12277)
);

INVx1_ASAP7_75t_L g12278 ( 
.A(n_10619),
.Y(n_12278)
);

OAI221xp5_ASAP7_75t_L g12279 ( 
.A1(n_11392),
.A2(n_9804),
.B1(n_9884),
.B2(n_9630),
.C(n_9612),
.Y(n_12279)
);

AOI22xp33_ASAP7_75t_SL g12280 ( 
.A1(n_10621),
.A2(n_8813),
.B1(n_8817),
.B2(n_10651),
.Y(n_12280)
);

NOR2x1_ASAP7_75t_SL g12281 ( 
.A(n_11010),
.B(n_9134),
.Y(n_12281)
);

AOI22xp5_ASAP7_75t_L g12282 ( 
.A1(n_10651),
.A2(n_9965),
.B1(n_10168),
.B2(n_10044),
.Y(n_12282)
);

AOI22xp33_ASAP7_75t_L g12283 ( 
.A1(n_10919),
.A2(n_8603),
.B1(n_8637),
.B2(n_8630),
.Y(n_12283)
);

INVx2_ASAP7_75t_L g12284 ( 
.A(n_10663),
.Y(n_12284)
);

OR2x6_ASAP7_75t_L g12285 ( 
.A(n_10511),
.B(n_9227),
.Y(n_12285)
);

AOI22xp33_ASAP7_75t_L g12286 ( 
.A1(n_10943),
.A2(n_8637),
.B1(n_8399),
.B2(n_7877),
.Y(n_12286)
);

OAI22xp33_ASAP7_75t_L g12287 ( 
.A1(n_10529),
.A2(n_8637),
.B1(n_10201),
.B2(n_10099),
.Y(n_12287)
);

AOI22xp33_ASAP7_75t_L g12288 ( 
.A1(n_10943),
.A2(n_8399),
.B1(n_7877),
.B2(n_7947),
.Y(n_12288)
);

OAI22xp33_ASAP7_75t_L g12289 ( 
.A1(n_10580),
.A2(n_10768),
.B1(n_10795),
.B2(n_10760),
.Y(n_12289)
);

OAI21xp5_ASAP7_75t_L g12290 ( 
.A1(n_10580),
.A2(n_8025),
.B(n_7966),
.Y(n_12290)
);

NOR2xp33_ASAP7_75t_L g12291 ( 
.A(n_10913),
.B(n_9487),
.Y(n_12291)
);

AOI21xp5_ASAP7_75t_L g12292 ( 
.A1(n_11247),
.A2(n_11301),
.B(n_9581),
.Y(n_12292)
);

OAI221xp5_ASAP7_75t_L g12293 ( 
.A1(n_10760),
.A2(n_9884),
.B1(n_9887),
.B2(n_9804),
.C(n_9630),
.Y(n_12293)
);

OAI322xp33_ASAP7_75t_L g12294 ( 
.A1(n_10677),
.A2(n_10238),
.A3(n_10341),
.B1(n_10201),
.B2(n_8845),
.C1(n_8594),
.C2(n_10363),
.Y(n_12294)
);

AOI22xp33_ASAP7_75t_L g12295 ( 
.A1(n_10966),
.A2(n_8399),
.B1(n_7877),
.B2(n_7947),
.Y(n_12295)
);

OR2x2_ASAP7_75t_L g12296 ( 
.A(n_10938),
.B(n_8872),
.Y(n_12296)
);

AOI22xp5_ASAP7_75t_L g12297 ( 
.A1(n_10966),
.A2(n_9965),
.B1(n_10168),
.B2(n_10044),
.Y(n_12297)
);

AOI21xp33_ASAP7_75t_SL g12298 ( 
.A1(n_11010),
.A2(n_9603),
.B(n_9499),
.Y(n_12298)
);

AOI22xp33_ASAP7_75t_SL g12299 ( 
.A1(n_10971),
.A2(n_7892),
.B1(n_8095),
.B2(n_7861),
.Y(n_12299)
);

AND2x2_ASAP7_75t_L g12300 ( 
.A(n_10971),
.B(n_9291),
.Y(n_12300)
);

INVx5_ASAP7_75t_L g12301 ( 
.A(n_10683),
.Y(n_12301)
);

AOI21xp5_ASAP7_75t_L g12302 ( 
.A1(n_11301),
.A2(n_9796),
.B(n_8370),
.Y(n_12302)
);

OAI22xp33_ASAP7_75t_L g12303 ( 
.A1(n_10768),
.A2(n_10238),
.B1(n_10341),
.B2(n_8399),
.Y(n_12303)
);

AOI211xp5_ASAP7_75t_L g12304 ( 
.A1(n_10795),
.A2(n_9526),
.B(n_9681),
.C(n_9604),
.Y(n_12304)
);

OAI221xp5_ASAP7_75t_L g12305 ( 
.A1(n_10857),
.A2(n_9804),
.B1(n_9887),
.B2(n_9884),
.C(n_9630),
.Y(n_12305)
);

AOI22xp33_ASAP7_75t_L g12306 ( 
.A1(n_10991),
.A2(n_8399),
.B1(n_7877),
.B2(n_7947),
.Y(n_12306)
);

OAI22xp5_ASAP7_75t_L g12307 ( 
.A1(n_10991),
.A2(n_8962),
.B1(n_8959),
.B2(n_6982),
.Y(n_12307)
);

AND2x2_ASAP7_75t_L g12308 ( 
.A(n_11003),
.B(n_11004),
.Y(n_12308)
);

A2O1A1Ixp33_ASAP7_75t_L g12309 ( 
.A1(n_10516),
.A2(n_8785),
.B(n_8665),
.C(n_7915),
.Y(n_12309)
);

AOI22xp33_ASAP7_75t_L g12310 ( 
.A1(n_11003),
.A2(n_7877),
.B1(n_7947),
.B2(n_7712),
.Y(n_12310)
);

NAND3xp33_ASAP7_75t_L g12311 ( 
.A(n_10696),
.B(n_7741),
.C(n_9526),
.Y(n_12311)
);

AOI22xp33_ASAP7_75t_L g12312 ( 
.A1(n_11004),
.A2(n_7877),
.B1(n_7947),
.B2(n_7712),
.Y(n_12312)
);

OAI221xp5_ASAP7_75t_L g12313 ( 
.A1(n_10857),
.A2(n_9887),
.B1(n_9960),
.B2(n_9919),
.C(n_9884),
.Y(n_12313)
);

AOI22xp33_ASAP7_75t_L g12314 ( 
.A1(n_11008),
.A2(n_7877),
.B1(n_7947),
.B2(n_7712),
.Y(n_12314)
);

AND2x2_ASAP7_75t_L g12315 ( 
.A(n_11008),
.B(n_9291),
.Y(n_12315)
);

HB1xp67_ASAP7_75t_L g12316 ( 
.A(n_11310),
.Y(n_12316)
);

AND2x2_ASAP7_75t_SL g12317 ( 
.A(n_11029),
.B(n_8896),
.Y(n_12317)
);

OAI22xp5_ASAP7_75t_SL g12318 ( 
.A1(n_10858),
.A2(n_7690),
.B1(n_7684),
.B2(n_7472),
.Y(n_12318)
);

AOI22xp33_ASAP7_75t_L g12319 ( 
.A1(n_11029),
.A2(n_7947),
.B1(n_8059),
.B2(n_7712),
.Y(n_12319)
);

INVx1_ASAP7_75t_L g12320 ( 
.A(n_10626),
.Y(n_12320)
);

AOI22xp33_ASAP7_75t_SL g12321 ( 
.A1(n_11038),
.A2(n_8095),
.B1(n_7861),
.B2(n_8166),
.Y(n_12321)
);

AOI22xp33_ASAP7_75t_L g12322 ( 
.A1(n_11038),
.A2(n_8059),
.B1(n_8162),
.B2(n_7712),
.Y(n_12322)
);

AOI21xp33_ASAP7_75t_L g12323 ( 
.A1(n_10858),
.A2(n_9604),
.B(n_9526),
.Y(n_12323)
);

INVx2_ASAP7_75t_L g12324 ( 
.A(n_10683),
.Y(n_12324)
);

OAI22xp33_ASAP7_75t_L g12325 ( 
.A1(n_10862),
.A2(n_8962),
.B1(n_8959),
.B2(n_8954),
.Y(n_12325)
);

INVx1_ASAP7_75t_L g12326 ( 
.A(n_10627),
.Y(n_12326)
);

CKINVDCx5p33_ASAP7_75t_R g12327 ( 
.A(n_10685),
.Y(n_12327)
);

AOI22xp33_ASAP7_75t_SL g12328 ( 
.A1(n_11315),
.A2(n_8095),
.B1(n_7861),
.B2(n_8166),
.Y(n_12328)
);

OAI221xp5_ASAP7_75t_L g12329 ( 
.A1(n_10862),
.A2(n_9919),
.B1(n_10051),
.B2(n_9960),
.C(n_9887),
.Y(n_12329)
);

AND2x4_ASAP7_75t_L g12330 ( 
.A(n_10683),
.B(n_10169),
.Y(n_12330)
);

CKINVDCx5p33_ASAP7_75t_R g12331 ( 
.A(n_11006),
.Y(n_12331)
);

AOI22xp33_ASAP7_75t_L g12332 ( 
.A1(n_11096),
.A2(n_8059),
.B1(n_8162),
.B2(n_7712),
.Y(n_12332)
);

AOI21xp33_ASAP7_75t_SL g12333 ( 
.A1(n_10906),
.A2(n_9976),
.B(n_9880),
.Y(n_12333)
);

INVx2_ASAP7_75t_L g12334 ( 
.A(n_10685),
.Y(n_12334)
);

AOI21xp33_ASAP7_75t_R g12335 ( 
.A1(n_10685),
.A2(n_9960),
.B(n_9919),
.Y(n_12335)
);

OAI211xp5_ASAP7_75t_L g12336 ( 
.A1(n_10687),
.A2(n_9655),
.B(n_9517),
.C(n_9426),
.Y(n_12336)
);

OAI21xp5_ASAP7_75t_L g12337 ( 
.A1(n_10906),
.A2(n_7966),
.B(n_7965),
.Y(n_12337)
);

NAND2xp5_ASAP7_75t_L g12338 ( 
.A(n_11016),
.B(n_8461),
.Y(n_12338)
);

INVx1_ASAP7_75t_L g12339 ( 
.A(n_10629),
.Y(n_12339)
);

OAI22xp5_ASAP7_75t_L g12340 ( 
.A1(n_10938),
.A2(n_8962),
.B1(n_6982),
.B2(n_7140),
.Y(n_12340)
);

AND2x2_ASAP7_75t_L g12341 ( 
.A(n_11096),
.B(n_9318),
.Y(n_12341)
);

INVxp67_ASAP7_75t_L g12342 ( 
.A(n_11043),
.Y(n_12342)
);

OAI211xp5_ASAP7_75t_L g12343 ( 
.A1(n_10687),
.A2(n_9655),
.B(n_9517),
.C(n_9426),
.Y(n_12343)
);

AOI22xp5_ASAP7_75t_L g12344 ( 
.A1(n_11140),
.A2(n_10198),
.B1(n_10169),
.B2(n_7964),
.Y(n_12344)
);

AOI221xp5_ASAP7_75t_L g12345 ( 
.A1(n_11315),
.A2(n_8462),
.B1(n_8259),
.B2(n_8261),
.C(n_9083),
.Y(n_12345)
);

OAI221xp5_ASAP7_75t_L g12346 ( 
.A1(n_11043),
.A2(n_9960),
.B1(n_10057),
.B2(n_10051),
.C(n_9919),
.Y(n_12346)
);

AOI22xp33_ASAP7_75t_L g12347 ( 
.A1(n_11140),
.A2(n_8059),
.B1(n_8162),
.B2(n_7712),
.Y(n_12347)
);

AND2x4_ASAP7_75t_L g12348 ( 
.A(n_10687),
.B(n_10169),
.Y(n_12348)
);

NAND2xp5_ASAP7_75t_SL g12349 ( 
.A(n_11016),
.B(n_9678),
.Y(n_12349)
);

INVx1_ASAP7_75t_L g12350 ( 
.A(n_10636),
.Y(n_12350)
);

AND2x4_ASAP7_75t_L g12351 ( 
.A(n_10692),
.B(n_10169),
.Y(n_12351)
);

AOI22xp33_ASAP7_75t_SL g12352 ( 
.A1(n_11329),
.A2(n_8095),
.B1(n_7861),
.B2(n_8166),
.Y(n_12352)
);

INVx1_ASAP7_75t_L g12353 ( 
.A(n_10637),
.Y(n_12353)
);

AOI22xp33_ASAP7_75t_SL g12354 ( 
.A1(n_11329),
.A2(n_8095),
.B1(n_7861),
.B2(n_8166),
.Y(n_12354)
);

AOI211xp5_ASAP7_75t_L g12355 ( 
.A1(n_11055),
.A2(n_9526),
.B(n_9681),
.C(n_9604),
.Y(n_12355)
);

INVx1_ASAP7_75t_L g12356 ( 
.A(n_10639),
.Y(n_12356)
);

INVx4_ASAP7_75t_L g12357 ( 
.A(n_10692),
.Y(n_12357)
);

OAI22xp5_ASAP7_75t_L g12358 ( 
.A1(n_11022),
.A2(n_8962),
.B1(n_6982),
.B2(n_7140),
.Y(n_12358)
);

INVx1_ASAP7_75t_L g12359 ( 
.A(n_10646),
.Y(n_12359)
);

NAND2xp5_ASAP7_75t_L g12360 ( 
.A(n_11022),
.B(n_10129),
.Y(n_12360)
);

AOI22xp33_ASAP7_75t_L g12361 ( 
.A1(n_11146),
.A2(n_8059),
.B1(n_8162),
.B2(n_10198),
.Y(n_12361)
);

AOI22xp33_ASAP7_75t_L g12362 ( 
.A1(n_11146),
.A2(n_8059),
.B1(n_8162),
.B2(n_10198),
.Y(n_12362)
);

INVx1_ASAP7_75t_L g12363 ( 
.A(n_10650),
.Y(n_12363)
);

AOI22xp33_ASAP7_75t_L g12364 ( 
.A1(n_11174),
.A2(n_8059),
.B1(n_8162),
.B2(n_10198),
.Y(n_12364)
);

AOI22xp33_ASAP7_75t_L g12365 ( 
.A1(n_11174),
.A2(n_8162),
.B1(n_8208),
.B2(n_8160),
.Y(n_12365)
);

HB1xp67_ASAP7_75t_L g12366 ( 
.A(n_11334),
.Y(n_12366)
);

AOI22xp33_ASAP7_75t_L g12367 ( 
.A1(n_11192),
.A2(n_8160),
.B1(n_8208),
.B2(n_8166),
.Y(n_12367)
);

AOI211xp5_ASAP7_75t_L g12368 ( 
.A1(n_11055),
.A2(n_9604),
.B(n_9708),
.C(n_9681),
.Y(n_12368)
);

INVx2_ASAP7_75t_L g12369 ( 
.A(n_10692),
.Y(n_12369)
);

AOI22xp33_ASAP7_75t_L g12370 ( 
.A1(n_11192),
.A2(n_8962),
.B1(n_7828),
.B2(n_7761),
.Y(n_12370)
);

BUFx3_ASAP7_75t_L g12371 ( 
.A(n_10701),
.Y(n_12371)
);

AOI22xp33_ASAP7_75t_L g12372 ( 
.A1(n_11041),
.A2(n_7828),
.B1(n_7761),
.B2(n_7778),
.Y(n_12372)
);

INVx2_ASAP7_75t_SL g12373 ( 
.A(n_10701),
.Y(n_12373)
);

AOI22xp33_ASAP7_75t_L g12374 ( 
.A1(n_11041),
.A2(n_7828),
.B1(n_7761),
.B2(n_7778),
.Y(n_12374)
);

INVx1_ASAP7_75t_L g12375 ( 
.A(n_10653),
.Y(n_12375)
);

INVx2_ASAP7_75t_L g12376 ( 
.A(n_10701),
.Y(n_12376)
);

BUFx3_ASAP7_75t_L g12377 ( 
.A(n_10731),
.Y(n_12377)
);

AOI221xp5_ASAP7_75t_L g12378 ( 
.A1(n_11334),
.A2(n_8259),
.B1(n_9089),
.B2(n_9084),
.C(n_9083),
.Y(n_12378)
);

AOI22xp33_ASAP7_75t_L g12379 ( 
.A1(n_11049),
.A2(n_7828),
.B1(n_7761),
.B2(n_7778),
.Y(n_12379)
);

OAI211xp5_ASAP7_75t_L g12380 ( 
.A1(n_10731),
.A2(n_9655),
.B(n_9517),
.C(n_9426),
.Y(n_12380)
);

AND2x2_ASAP7_75t_L g12381 ( 
.A(n_11049),
.B(n_9318),
.Y(n_12381)
);

INVx2_ASAP7_75t_L g12382 ( 
.A(n_10731),
.Y(n_12382)
);

AOI22xp33_ASAP7_75t_L g12383 ( 
.A1(n_11077),
.A2(n_7828),
.B1(n_7761),
.B2(n_7778),
.Y(n_12383)
);

INVx1_ASAP7_75t_L g12384 ( 
.A(n_10659),
.Y(n_12384)
);

AOI22xp33_ASAP7_75t_L g12385 ( 
.A1(n_11077),
.A2(n_7778),
.B1(n_7755),
.B2(n_7992),
.Y(n_12385)
);

BUFx12f_ASAP7_75t_L g12386 ( 
.A(n_11069),
.Y(n_12386)
);

AOI221xp5_ASAP7_75t_L g12387 ( 
.A1(n_11345),
.A2(n_9084),
.B1(n_9096),
.B2(n_9089),
.C(n_9083),
.Y(n_12387)
);

NAND3xp33_ASAP7_75t_L g12388 ( 
.A(n_10696),
.B(n_7741),
.C(n_9604),
.Y(n_12388)
);

AOI222xp33_ASAP7_75t_L g12389 ( 
.A1(n_11345),
.A2(n_7848),
.B1(n_7954),
.B2(n_10363),
.C1(n_8701),
.C2(n_8518),
.Y(n_12389)
);

INVx1_ASAP7_75t_L g12390 ( 
.A(n_10662),
.Y(n_12390)
);

INVx1_ASAP7_75t_L g12391 ( 
.A(n_10664),
.Y(n_12391)
);

HB1xp67_ASAP7_75t_L g12392 ( 
.A(n_11359),
.Y(n_12392)
);

OAI22xp5_ASAP7_75t_L g12393 ( 
.A1(n_11069),
.A2(n_6982),
.B1(n_7140),
.B2(n_7426),
.Y(n_12393)
);

OAI21xp33_ASAP7_75t_L g12394 ( 
.A1(n_10392),
.A2(n_8328),
.B(n_8316),
.Y(n_12394)
);

AOI22xp5_ASAP7_75t_L g12395 ( 
.A1(n_11396),
.A2(n_7964),
.B1(n_8870),
.B2(n_8841),
.Y(n_12395)
);

AOI22xp33_ASAP7_75t_L g12396 ( 
.A1(n_11088),
.A2(n_7755),
.B1(n_8415),
.B2(n_7992),
.Y(n_12396)
);

OAI21x1_ASAP7_75t_L g12397 ( 
.A1(n_10770),
.A2(n_10689),
.B(n_10595),
.Y(n_12397)
);

OAI22xp33_ASAP7_75t_L g12398 ( 
.A1(n_11076),
.A2(n_8954),
.B1(n_8896),
.B2(n_8952),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_11088),
.A2(n_7755),
.B1(n_8415),
.B2(n_7992),
.Y(n_12399)
);

AND2x2_ASAP7_75t_L g12400 ( 
.A(n_11396),
.B(n_9341),
.Y(n_12400)
);

NAND3xp33_ASAP7_75t_L g12401 ( 
.A(n_10750),
.B(n_7741),
.C(n_9604),
.Y(n_12401)
);

INVx2_ASAP7_75t_L g12402 ( 
.A(n_10744),
.Y(n_12402)
);

OAI22xp5_ASAP7_75t_L g12403 ( 
.A1(n_11076),
.A2(n_6982),
.B1(n_7140),
.B2(n_7426),
.Y(n_12403)
);

NAND2xp5_ASAP7_75t_SL g12404 ( 
.A(n_11037),
.B(n_9678),
.Y(n_12404)
);

NAND3xp33_ASAP7_75t_L g12405 ( 
.A(n_10750),
.B(n_7741),
.C(n_9681),
.Y(n_12405)
);

AOI221xp5_ASAP7_75t_L g12406 ( 
.A1(n_11359),
.A2(n_9089),
.B1(n_9122),
.B2(n_9096),
.C(n_9084),
.Y(n_12406)
);

INVx1_ASAP7_75t_L g12407 ( 
.A(n_10665),
.Y(n_12407)
);

INVx1_ASAP7_75t_L g12408 ( 
.A(n_10666),
.Y(n_12408)
);

OAI22xp33_ASAP7_75t_L g12409 ( 
.A1(n_11091),
.A2(n_8954),
.B1(n_8896),
.B2(n_8952),
.Y(n_12409)
);

OR2x2_ASAP7_75t_L g12410 ( 
.A(n_10392),
.B(n_8872),
.Y(n_12410)
);

AO21x2_ASAP7_75t_L g12411 ( 
.A1(n_10406),
.A2(n_9511),
.B(n_9443),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_10668),
.Y(n_12412)
);

AOI22xp33_ASAP7_75t_L g12413 ( 
.A1(n_11210),
.A2(n_7755),
.B1(n_8415),
.B2(n_7992),
.Y(n_12413)
);

INVx1_ASAP7_75t_L g12414 ( 
.A(n_10669),
.Y(n_12414)
);

AOI221xp5_ASAP7_75t_L g12415 ( 
.A1(n_11361),
.A2(n_11364),
.B1(n_10412),
.B2(n_10407),
.C(n_11401),
.Y(n_12415)
);

AOI22xp33_ASAP7_75t_L g12416 ( 
.A1(n_11210),
.A2(n_7755),
.B1(n_8415),
.B2(n_7992),
.Y(n_12416)
);

OAI22xp5_ASAP7_75t_L g12417 ( 
.A1(n_11091),
.A2(n_7140),
.B1(n_7465),
.B2(n_7464),
.Y(n_12417)
);

AOI21xp5_ASAP7_75t_L g12418 ( 
.A1(n_10589),
.A2(n_8961),
.B(n_9655),
.Y(n_12418)
);

AND2x2_ASAP7_75t_L g12419 ( 
.A(n_11401),
.B(n_9341),
.Y(n_12419)
);

NAND2xp5_ASAP7_75t_L g12420 ( 
.A(n_11432),
.B(n_10129),
.Y(n_12420)
);

INVx2_ASAP7_75t_L g12421 ( 
.A(n_10744),
.Y(n_12421)
);

INVx2_ASAP7_75t_L g12422 ( 
.A(n_10744),
.Y(n_12422)
);

INVx2_ASAP7_75t_L g12423 ( 
.A(n_10769),
.Y(n_12423)
);

A2O1A1Ixp33_ASAP7_75t_L g12424 ( 
.A1(n_10516),
.A2(n_8665),
.B(n_7915),
.C(n_7965),
.Y(n_12424)
);

INVx2_ASAP7_75t_SL g12425 ( 
.A(n_10769),
.Y(n_12425)
);

BUFx6f_ASAP7_75t_L g12426 ( 
.A(n_10769),
.Y(n_12426)
);

OAI22xp33_ASAP7_75t_L g12427 ( 
.A1(n_11093),
.A2(n_8954),
.B1(n_8896),
.B2(n_8952),
.Y(n_12427)
);

A2O1A1Ixp33_ASAP7_75t_L g12428 ( 
.A1(n_10543),
.A2(n_8665),
.B(n_7915),
.C(n_7965),
.Y(n_12428)
);

HB1xp67_ASAP7_75t_L g12429 ( 
.A(n_11361),
.Y(n_12429)
);

BUFx4f_ASAP7_75t_SL g12430 ( 
.A(n_10823),
.Y(n_12430)
);

INVx2_ASAP7_75t_L g12431 ( 
.A(n_10823),
.Y(n_12431)
);

AOI21xp33_ASAP7_75t_L g12432 ( 
.A1(n_11093),
.A2(n_9708),
.B(n_9681),
.Y(n_12432)
);

AOI31xp33_ASAP7_75t_SL g12433 ( 
.A1(n_11037),
.A2(n_8794),
.A3(n_7717),
.B(n_7872),
.Y(n_12433)
);

INVx1_ASAP7_75t_L g12434 ( 
.A(n_10678),
.Y(n_12434)
);

INVx1_ASAP7_75t_L g12435 ( 
.A(n_10682),
.Y(n_12435)
);

BUFx2_ASAP7_75t_L g12436 ( 
.A(n_10823),
.Y(n_12436)
);

AOI221xp5_ASAP7_75t_L g12437 ( 
.A1(n_11364),
.A2(n_9123),
.B1(n_9122),
.B2(n_9096),
.C(n_9979),
.Y(n_12437)
);

INVx1_ASAP7_75t_SL g12438 ( 
.A(n_11432),
.Y(n_12438)
);

OAI22xp5_ASAP7_75t_SL g12439 ( 
.A1(n_11145),
.A2(n_7690),
.B1(n_7684),
.B2(n_7472),
.Y(n_12439)
);

AOI22xp33_ASAP7_75t_SL g12440 ( 
.A1(n_11436),
.A2(n_8918),
.B1(n_8979),
.B2(n_8873),
.Y(n_12440)
);

AOI22xp33_ASAP7_75t_SL g12441 ( 
.A1(n_11436),
.A2(n_8979),
.B1(n_8961),
.B2(n_8923),
.Y(n_12441)
);

OAI211xp5_ASAP7_75t_SL g12442 ( 
.A1(n_10844),
.A2(n_10057),
.B(n_10062),
.C(n_10051),
.Y(n_12442)
);

AOI22x1_ASAP7_75t_SL g12443 ( 
.A1(n_10844),
.A2(n_7476),
.B1(n_7469),
.B2(n_7439),
.Y(n_12443)
);

AOI22xp33_ASAP7_75t_L g12444 ( 
.A1(n_11214),
.A2(n_7992),
.B1(n_8415),
.B2(n_11232),
.Y(n_12444)
);

AOI22xp33_ASAP7_75t_L g12445 ( 
.A1(n_11214),
.A2(n_7992),
.B1(n_8415),
.B2(n_7964),
.Y(n_12445)
);

AOI21xp5_ASAP7_75t_L g12446 ( 
.A1(n_10589),
.A2(n_8961),
.B(n_9426),
.Y(n_12446)
);

NAND3xp33_ASAP7_75t_L g12447 ( 
.A(n_10764),
.B(n_7741),
.C(n_9681),
.Y(n_12447)
);

AOI22xp33_ASAP7_75t_L g12448 ( 
.A1(n_11232),
.A2(n_7992),
.B1(n_8415),
.B2(n_7964),
.Y(n_12448)
);

INVx1_ASAP7_75t_L g12449 ( 
.A(n_10684),
.Y(n_12449)
);

CKINVDCx11_ASAP7_75t_R g12450 ( 
.A(n_10407),
.Y(n_12450)
);

AND2x2_ASAP7_75t_L g12451 ( 
.A(n_11461),
.B(n_9394),
.Y(n_12451)
);

AOI21xp33_ASAP7_75t_L g12452 ( 
.A1(n_11145),
.A2(n_9730),
.B(n_9708),
.Y(n_12452)
);

BUFx3_ASAP7_75t_L g12453 ( 
.A(n_10844),
.Y(n_12453)
);

INVx1_ASAP7_75t_L g12454 ( 
.A(n_10686),
.Y(n_12454)
);

AOI22xp33_ASAP7_75t_L g12455 ( 
.A1(n_11461),
.A2(n_7992),
.B1(n_8415),
.B2(n_11463),
.Y(n_12455)
);

AOI22xp33_ASAP7_75t_L g12456 ( 
.A1(n_11463),
.A2(n_7992),
.B1(n_8415),
.B2(n_7964),
.Y(n_12456)
);

NAND3xp33_ASAP7_75t_L g12457 ( 
.A(n_10764),
.B(n_7741),
.C(n_9708),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_10693),
.Y(n_12458)
);

OR2x2_ASAP7_75t_L g12459 ( 
.A(n_10633),
.B(n_8872),
.Y(n_12459)
);

NAND2x1p5_ASAP7_75t_L g12460 ( 
.A(n_10901),
.B(n_8953),
.Y(n_12460)
);

HB1xp67_ASAP7_75t_L g12461 ( 
.A(n_10494),
.Y(n_12461)
);

INVx1_ASAP7_75t_L g12462 ( 
.A(n_10695),
.Y(n_12462)
);

AOI22xp33_ASAP7_75t_L g12463 ( 
.A1(n_10679),
.A2(n_7992),
.B1(n_8415),
.B2(n_7964),
.Y(n_12463)
);

INVx4_ASAP7_75t_SL g12464 ( 
.A(n_10494),
.Y(n_12464)
);

AOI22xp33_ASAP7_75t_SL g12465 ( 
.A1(n_11249),
.A2(n_8961),
.B1(n_8952),
.B2(n_8923),
.Y(n_12465)
);

OAI22xp5_ASAP7_75t_L g12466 ( 
.A1(n_10901),
.A2(n_7465),
.B1(n_7489),
.B2(n_7464),
.Y(n_12466)
);

OAI211xp5_ASAP7_75t_L g12467 ( 
.A1(n_10901),
.A2(n_9517),
.B(n_9373),
.C(n_9351),
.Y(n_12467)
);

OAI221xp5_ASAP7_75t_L g12468 ( 
.A1(n_11175),
.A2(n_10057),
.B1(n_10072),
.B2(n_10062),
.C(n_10051),
.Y(n_12468)
);

OAI221xp5_ASAP7_75t_L g12469 ( 
.A1(n_11175),
.A2(n_10062),
.B1(n_10087),
.B2(n_10072),
.C(n_10057),
.Y(n_12469)
);

CKINVDCx11_ASAP7_75t_R g12470 ( 
.A(n_10412),
.Y(n_12470)
);

NAND4xp25_ASAP7_75t_SL g12471 ( 
.A(n_11269),
.B(n_9921),
.C(n_9394),
.D(n_9464),
.Y(n_12471)
);

BUFx6f_ASAP7_75t_L g12472 ( 
.A(n_10945),
.Y(n_12472)
);

AOI222xp33_ASAP7_75t_L g12473 ( 
.A1(n_11269),
.A2(n_8518),
.B1(n_8701),
.B2(n_7417),
.C1(n_7410),
.C2(n_9036),
.Y(n_12473)
);

INVx1_ASAP7_75t_L g12474 ( 
.A(n_10698),
.Y(n_12474)
);

AOI22xp33_ASAP7_75t_L g12475 ( 
.A1(n_10679),
.A2(n_7992),
.B1(n_8415),
.B2(n_7964),
.Y(n_12475)
);

AOI21xp33_ASAP7_75t_L g12476 ( 
.A1(n_10945),
.A2(n_9730),
.B(n_9708),
.Y(n_12476)
);

OAI221xp5_ASAP7_75t_L g12477 ( 
.A1(n_11175),
.A2(n_10072),
.B1(n_10090),
.B2(n_10087),
.C(n_10062),
.Y(n_12477)
);

AOI22xp33_ASAP7_75t_SL g12478 ( 
.A1(n_11273),
.A2(n_8961),
.B1(n_8952),
.B2(n_8923),
.Y(n_12478)
);

AOI221xp5_ASAP7_75t_L g12479 ( 
.A1(n_11273),
.A2(n_9123),
.B1(n_9122),
.B2(n_10098),
.C(n_9979),
.Y(n_12479)
);

NAND2xp5_ASAP7_75t_L g12480 ( 
.A(n_10633),
.B(n_10286),
.Y(n_12480)
);

AOI22xp33_ASAP7_75t_L g12481 ( 
.A1(n_10700),
.A2(n_8415),
.B1(n_8841),
.B2(n_7964),
.Y(n_12481)
);

AND2x4_ASAP7_75t_L g12482 ( 
.A(n_10945),
.B(n_9400),
.Y(n_12482)
);

OAI221xp5_ASAP7_75t_L g12483 ( 
.A1(n_11184),
.A2(n_10090),
.B1(n_10110),
.B2(n_10087),
.C(n_10072),
.Y(n_12483)
);

INVx1_ASAP7_75t_L g12484 ( 
.A(n_10706),
.Y(n_12484)
);

INVx2_ASAP7_75t_L g12485 ( 
.A(n_10995),
.Y(n_12485)
);

OR2x2_ASAP7_75t_L g12486 ( 
.A(n_10802),
.B(n_8872),
.Y(n_12486)
);

AOI22xp33_ASAP7_75t_L g12487 ( 
.A1(n_10700),
.A2(n_8841),
.B1(n_8870),
.B2(n_7964),
.Y(n_12487)
);

OR2x6_ASAP7_75t_L g12488 ( 
.A(n_10995),
.B(n_9708),
.Y(n_12488)
);

OAI22xp5_ASAP7_75t_L g12489 ( 
.A1(n_10995),
.A2(n_7465),
.B1(n_7489),
.B2(n_7464),
.Y(n_12489)
);

OR2x2_ASAP7_75t_L g12490 ( 
.A(n_10802),
.B(n_8872),
.Y(n_12490)
);

INVxp67_ASAP7_75t_L g12491 ( 
.A(n_10707),
.Y(n_12491)
);

CKINVDCx5p33_ASAP7_75t_R g12492 ( 
.A(n_11062),
.Y(n_12492)
);

AO31x2_ASAP7_75t_L g12493 ( 
.A1(n_10712),
.A2(n_9515),
.A3(n_9511),
.B(n_9189),
.Y(n_12493)
);

AOI221xp5_ASAP7_75t_L g12494 ( 
.A1(n_11520),
.A2(n_9123),
.B1(n_10098),
.B2(n_10227),
.C(n_9979),
.Y(n_12494)
);

INVx1_ASAP7_75t_L g12495 ( 
.A(n_10714),
.Y(n_12495)
);

HB1xp67_ASAP7_75t_L g12496 ( 
.A(n_10494),
.Y(n_12496)
);

AND2x2_ASAP7_75t_L g12497 ( 
.A(n_10722),
.B(n_9400),
.Y(n_12497)
);

OAI22xp5_ASAP7_75t_L g12498 ( 
.A1(n_11006),
.A2(n_7465),
.B1(n_7489),
.B2(n_7464),
.Y(n_12498)
);

INVx1_ASAP7_75t_L g12499 ( 
.A(n_10721),
.Y(n_12499)
);

BUFx6f_ASAP7_75t_L g12500 ( 
.A(n_11006),
.Y(n_12500)
);

INVx1_ASAP7_75t_L g12501 ( 
.A(n_10724),
.Y(n_12501)
);

AOI222xp33_ASAP7_75t_L g12502 ( 
.A1(n_10722),
.A2(n_7417),
.B1(n_9047),
.B2(n_9068),
.C1(n_9044),
.C2(n_6661),
.Y(n_12502)
);

INVx1_ASAP7_75t_L g12503 ( 
.A(n_10726),
.Y(n_12503)
);

NAND3xp33_ASAP7_75t_L g12504 ( 
.A(n_11061),
.B(n_9752),
.C(n_9730),
.Y(n_12504)
);

OAI22xp33_ASAP7_75t_SL g12505 ( 
.A1(n_11061),
.A2(n_10090),
.B1(n_10110),
.B2(n_10087),
.Y(n_12505)
);

OA21x2_ASAP7_75t_L g12506 ( 
.A1(n_10595),
.A2(n_9515),
.B(n_9195),
.Y(n_12506)
);

AO21x2_ASAP7_75t_L g12507 ( 
.A1(n_10507),
.A2(n_9515),
.B(n_9195),
.Y(n_12507)
);

AOI22xp33_ASAP7_75t_L g12508 ( 
.A1(n_10728),
.A2(n_8870),
.B1(n_8975),
.B2(n_8841),
.Y(n_12508)
);

OAI221xp5_ASAP7_75t_L g12509 ( 
.A1(n_11184),
.A2(n_10154),
.B1(n_10216),
.B2(n_10110),
.C(n_10090),
.Y(n_12509)
);

AOI22xp33_ASAP7_75t_L g12510 ( 
.A1(n_10728),
.A2(n_8870),
.B1(n_8975),
.B2(n_8841),
.Y(n_12510)
);

INVxp67_ASAP7_75t_L g12511 ( 
.A(n_10729),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_10736),
.Y(n_12512)
);

OAI22xp5_ASAP7_75t_L g12513 ( 
.A1(n_11061),
.A2(n_7504),
.B1(n_7505),
.B2(n_7489),
.Y(n_12513)
);

AOI22xp33_ASAP7_75t_L g12514 ( 
.A1(n_10741),
.A2(n_8870),
.B1(n_8975),
.B2(n_8841),
.Y(n_12514)
);

AND2x2_ASAP7_75t_L g12515 ( 
.A(n_10741),
.B(n_9464),
.Y(n_12515)
);

INVx1_ASAP7_75t_L g12516 ( 
.A(n_10737),
.Y(n_12516)
);

AOI221xp5_ASAP7_75t_L g12517 ( 
.A1(n_10738),
.A2(n_10227),
.B1(n_10228),
.B2(n_10098),
.C(n_9979),
.Y(n_12517)
);

AND2x4_ASAP7_75t_L g12518 ( 
.A(n_11062),
.B(n_10286),
.Y(n_12518)
);

OAI22xp33_ASAP7_75t_L g12519 ( 
.A1(n_11062),
.A2(n_8954),
.B1(n_8896),
.B2(n_8952),
.Y(n_12519)
);

OR2x2_ASAP7_75t_L g12520 ( 
.A(n_10887),
.B(n_8872),
.Y(n_12520)
);

OAI221xp5_ASAP7_75t_L g12521 ( 
.A1(n_11184),
.A2(n_10216),
.B1(n_10255),
.B2(n_10154),
.C(n_10110),
.Y(n_12521)
);

AOI22xp33_ASAP7_75t_L g12522 ( 
.A1(n_10749),
.A2(n_8870),
.B1(n_8975),
.B2(n_8841),
.Y(n_12522)
);

INVx1_ASAP7_75t_L g12523 ( 
.A(n_11542),
.Y(n_12523)
);

AND2x2_ASAP7_75t_L g12524 ( 
.A(n_11552),
.B(n_9678),
.Y(n_12524)
);

INVx1_ASAP7_75t_SL g12525 ( 
.A(n_12128),
.Y(n_12525)
);

OR2x2_ASAP7_75t_L g12526 ( 
.A(n_12093),
.B(n_12206),
.Y(n_12526)
);

INVx2_ASAP7_75t_L g12527 ( 
.A(n_11678),
.Y(n_12527)
);

BUFx2_ASAP7_75t_L g12528 ( 
.A(n_11700),
.Y(n_12528)
);

INVx2_ASAP7_75t_L g12529 ( 
.A(n_11896),
.Y(n_12529)
);

NAND2xp5_ASAP7_75t_L g12530 ( 
.A(n_11780),
.B(n_10494),
.Y(n_12530)
);

HB1xp67_ASAP7_75t_L g12531 ( 
.A(n_11707),
.Y(n_12531)
);

NAND2xp5_ASAP7_75t_L g12532 ( 
.A(n_11610),
.B(n_11739),
.Y(n_12532)
);

AOI22xp33_ASAP7_75t_L g12533 ( 
.A1(n_11558),
.A2(n_11258),
.B1(n_11272),
.B2(n_11197),
.Y(n_12533)
);

AND2x4_ASAP7_75t_L g12534 ( 
.A(n_11739),
.B(n_11068),
.Y(n_12534)
);

INVx1_ASAP7_75t_L g12535 ( 
.A(n_11725),
.Y(n_12535)
);

AND2x2_ASAP7_75t_L g12536 ( 
.A(n_11559),
.B(n_9487),
.Y(n_12536)
);

OR2x2_ASAP7_75t_L g12537 ( 
.A(n_12243),
.B(n_12064),
.Y(n_12537)
);

AND2x2_ASAP7_75t_L g12538 ( 
.A(n_11602),
.B(n_9487),
.Y(n_12538)
);

OR2x2_ASAP7_75t_L g12539 ( 
.A(n_12080),
.B(n_10887),
.Y(n_12539)
);

AND2x2_ASAP7_75t_L g12540 ( 
.A(n_11887),
.B(n_9627),
.Y(n_12540)
);

AND2x2_ASAP7_75t_SL g12541 ( 
.A(n_11879),
.B(n_11068),
.Y(n_12541)
);

HB1xp67_ASAP7_75t_L g12542 ( 
.A(n_12316),
.Y(n_12542)
);

INVx1_ASAP7_75t_L g12543 ( 
.A(n_11802),
.Y(n_12543)
);

BUFx3_ASAP7_75t_L g12544 ( 
.A(n_11669),
.Y(n_12544)
);

AND2x2_ASAP7_75t_L g12545 ( 
.A(n_11963),
.B(n_9627),
.Y(n_12545)
);

HB1xp67_ASAP7_75t_L g12546 ( 
.A(n_12366),
.Y(n_12546)
);

NAND2xp5_ASAP7_75t_L g12547 ( 
.A(n_11741),
.B(n_10740),
.Y(n_12547)
);

NAND2xp5_ASAP7_75t_L g12548 ( 
.A(n_11637),
.B(n_11768),
.Y(n_12548)
);

INVx1_ASAP7_75t_L g12549 ( 
.A(n_11907),
.Y(n_12549)
);

INVx1_ASAP7_75t_L g12550 ( 
.A(n_11918),
.Y(n_12550)
);

INVx2_ASAP7_75t_SL g12551 ( 
.A(n_11569),
.Y(n_12551)
);

INVx1_ASAP7_75t_L g12552 ( 
.A(n_11943),
.Y(n_12552)
);

INVx1_ASAP7_75t_L g12553 ( 
.A(n_12085),
.Y(n_12553)
);

AND2x4_ASAP7_75t_L g12554 ( 
.A(n_11974),
.B(n_11990),
.Y(n_12554)
);

INVx2_ASAP7_75t_L g12555 ( 
.A(n_11804),
.Y(n_12555)
);

INVx1_ASAP7_75t_L g12556 ( 
.A(n_12124),
.Y(n_12556)
);

BUFx2_ASAP7_75t_L g12557 ( 
.A(n_11700),
.Y(n_12557)
);

AND2x4_ASAP7_75t_SL g12558 ( 
.A(n_11581),
.B(n_11068),
.Y(n_12558)
);

AND2x2_ASAP7_75t_L g12559 ( 
.A(n_11973),
.B(n_10749),
.Y(n_12559)
);

AND2x2_ASAP7_75t_L g12560 ( 
.A(n_11996),
.B(n_10787),
.Y(n_12560)
);

INVx1_ASAP7_75t_L g12561 ( 
.A(n_12392),
.Y(n_12561)
);

BUFx2_ASAP7_75t_L g12562 ( 
.A(n_12226),
.Y(n_12562)
);

OR2x2_ASAP7_75t_L g12563 ( 
.A(n_12144),
.B(n_10740),
.Y(n_12563)
);

AND2x2_ASAP7_75t_L g12564 ( 
.A(n_12057),
.B(n_10787),
.Y(n_12564)
);

AND2x2_ASAP7_75t_L g12565 ( 
.A(n_11579),
.B(n_12078),
.Y(n_12565)
);

INVx2_ASAP7_75t_L g12566 ( 
.A(n_11804),
.Y(n_12566)
);

HB1xp67_ASAP7_75t_L g12567 ( 
.A(n_12429),
.Y(n_12567)
);

OR2x2_ASAP7_75t_L g12568 ( 
.A(n_12438),
.B(n_11567),
.Y(n_12568)
);

AND2x2_ASAP7_75t_L g12569 ( 
.A(n_12096),
.B(n_10794),
.Y(n_12569)
);

AND2x2_ASAP7_75t_L g12570 ( 
.A(n_11690),
.B(n_10794),
.Y(n_12570)
);

OR2x2_ASAP7_75t_L g12571 ( 
.A(n_11607),
.B(n_10740),
.Y(n_12571)
);

AND2x2_ASAP7_75t_L g12572 ( 
.A(n_11603),
.B(n_10816),
.Y(n_12572)
);

INVx1_ASAP7_75t_SL g12573 ( 
.A(n_11751),
.Y(n_12573)
);

INVx1_ASAP7_75t_L g12574 ( 
.A(n_11668),
.Y(n_12574)
);

AND2x2_ASAP7_75t_L g12575 ( 
.A(n_11734),
.B(n_10816),
.Y(n_12575)
);

INVx3_ASAP7_75t_SL g12576 ( 
.A(n_11937),
.Y(n_12576)
);

INVx1_ASAP7_75t_L g12577 ( 
.A(n_11683),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_11711),
.Y(n_12578)
);

INVx2_ASAP7_75t_L g12579 ( 
.A(n_11874),
.Y(n_12579)
);

AND2x2_ASAP7_75t_L g12580 ( 
.A(n_12154),
.B(n_10832),
.Y(n_12580)
);

INVx2_ASAP7_75t_L g12581 ( 
.A(n_11874),
.Y(n_12581)
);

INVx2_ASAP7_75t_L g12582 ( 
.A(n_12024),
.Y(n_12582)
);

HB1xp67_ASAP7_75t_L g12583 ( 
.A(n_12436),
.Y(n_12583)
);

AND2x2_ASAP7_75t_L g12584 ( 
.A(n_12175),
.B(n_10832),
.Y(n_12584)
);

INVx4_ASAP7_75t_L g12585 ( 
.A(n_11554),
.Y(n_12585)
);

INVx1_ASAP7_75t_L g12586 ( 
.A(n_11718),
.Y(n_12586)
);

INVx2_ASAP7_75t_L g12587 ( 
.A(n_12024),
.Y(n_12587)
);

AOI22xp33_ASAP7_75t_L g12588 ( 
.A1(n_11606),
.A2(n_11258),
.B1(n_11272),
.B2(n_11197),
.Y(n_12588)
);

INVx3_ASAP7_75t_L g12589 ( 
.A(n_11554),
.Y(n_12589)
);

AND2x4_ASAP7_75t_L g12590 ( 
.A(n_12116),
.B(n_11157),
.Y(n_12590)
);

BUFx2_ASAP7_75t_L g12591 ( 
.A(n_12226),
.Y(n_12591)
);

INVx1_ASAP7_75t_L g12592 ( 
.A(n_11723),
.Y(n_12592)
);

INVx2_ASAP7_75t_L g12593 ( 
.A(n_12072),
.Y(n_12593)
);

INVx1_ASAP7_75t_L g12594 ( 
.A(n_11744),
.Y(n_12594)
);

AND2x2_ASAP7_75t_L g12595 ( 
.A(n_12156),
.B(n_10834),
.Y(n_12595)
);

BUFx2_ASAP7_75t_L g12596 ( 
.A(n_11554),
.Y(n_12596)
);

AND2x2_ASAP7_75t_L g12597 ( 
.A(n_12156),
.B(n_10834),
.Y(n_12597)
);

INVx2_ASAP7_75t_L g12598 ( 
.A(n_12072),
.Y(n_12598)
);

INVx1_ASAP7_75t_L g12599 ( 
.A(n_11747),
.Y(n_12599)
);

INVxp67_ASAP7_75t_L g12600 ( 
.A(n_11546),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_11752),
.Y(n_12601)
);

BUFx3_ASAP7_75t_L g12602 ( 
.A(n_11570),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_11761),
.Y(n_12603)
);

INVx1_ASAP7_75t_L g12604 ( 
.A(n_11763),
.Y(n_12604)
);

AND2x2_ASAP7_75t_L g12605 ( 
.A(n_12130),
.B(n_10876),
.Y(n_12605)
);

INVx1_ASAP7_75t_L g12606 ( 
.A(n_11771),
.Y(n_12606)
);

BUFx6f_ASAP7_75t_L g12607 ( 
.A(n_11570),
.Y(n_12607)
);

INVx2_ASAP7_75t_L g12608 ( 
.A(n_12301),
.Y(n_12608)
);

AND2x2_ASAP7_75t_L g12609 ( 
.A(n_12143),
.B(n_10876),
.Y(n_12609)
);

INVx2_ASAP7_75t_SL g12610 ( 
.A(n_11569),
.Y(n_12610)
);

INVx1_ASAP7_75t_L g12611 ( 
.A(n_11778),
.Y(n_12611)
);

AND2x2_ASAP7_75t_L g12612 ( 
.A(n_12147),
.B(n_10877),
.Y(n_12612)
);

INVxp67_ASAP7_75t_L g12613 ( 
.A(n_11570),
.Y(n_12613)
);

AND2x2_ASAP7_75t_L g12614 ( 
.A(n_12151),
.B(n_10877),
.Y(n_12614)
);

AND2x2_ASAP7_75t_L g12615 ( 
.A(n_12285),
.B(n_9475),
.Y(n_12615)
);

INVx1_ASAP7_75t_L g12616 ( 
.A(n_11788),
.Y(n_12616)
);

INVx3_ASAP7_75t_SL g12617 ( 
.A(n_11945),
.Y(n_12617)
);

OR2x2_ASAP7_75t_L g12618 ( 
.A(n_11712),
.B(n_10740),
.Y(n_12618)
);

INVx2_ASAP7_75t_L g12619 ( 
.A(n_12301),
.Y(n_12619)
);

INVx2_ASAP7_75t_L g12620 ( 
.A(n_12301),
.Y(n_12620)
);

INVx1_ASAP7_75t_L g12621 ( 
.A(n_11792),
.Y(n_12621)
);

AND2x2_ASAP7_75t_L g12622 ( 
.A(n_12285),
.B(n_9475),
.Y(n_12622)
);

INVx3_ASAP7_75t_L g12623 ( 
.A(n_12254),
.Y(n_12623)
);

AND2x2_ASAP7_75t_L g12624 ( 
.A(n_11677),
.B(n_9494),
.Y(n_12624)
);

INVx2_ASAP7_75t_SL g12625 ( 
.A(n_11569),
.Y(n_12625)
);

INVx2_ASAP7_75t_L g12626 ( 
.A(n_12019),
.Y(n_12626)
);

HB1xp67_ASAP7_75t_L g12627 ( 
.A(n_12464),
.Y(n_12627)
);

OAI222xp33_ASAP7_75t_L g12628 ( 
.A1(n_11622),
.A2(n_11157),
.B1(n_11272),
.B2(n_11276),
.C1(n_11258),
.C2(n_11197),
.Y(n_12628)
);

NAND2xp5_ASAP7_75t_L g12629 ( 
.A(n_11595),
.B(n_10739),
.Y(n_12629)
);

AND2x4_ASAP7_75t_L g12630 ( 
.A(n_12116),
.B(n_11625),
.Y(n_12630)
);

AND2x2_ASAP7_75t_L g12631 ( 
.A(n_11677),
.B(n_9494),
.Y(n_12631)
);

INVx4_ASAP7_75t_L g12632 ( 
.A(n_11581),
.Y(n_12632)
);

AND2x2_ASAP7_75t_L g12633 ( 
.A(n_11708),
.B(n_9495),
.Y(n_12633)
);

HB1xp67_ASAP7_75t_L g12634 ( 
.A(n_12464),
.Y(n_12634)
);

INVx1_ASAP7_75t_L g12635 ( 
.A(n_11801),
.Y(n_12635)
);

INVx2_ASAP7_75t_L g12636 ( 
.A(n_12240),
.Y(n_12636)
);

AND2x2_ASAP7_75t_L g12637 ( 
.A(n_11708),
.B(n_9495),
.Y(n_12637)
);

INVx2_ASAP7_75t_SL g12638 ( 
.A(n_11766),
.Y(n_12638)
);

NAND2x1_ASAP7_75t_L g12639 ( 
.A(n_11625),
.B(n_11157),
.Y(n_12639)
);

AND2x2_ASAP7_75t_L g12640 ( 
.A(n_12173),
.B(n_9927),
.Y(n_12640)
);

INVx1_ASAP7_75t_L g12641 ( 
.A(n_11811),
.Y(n_12641)
);

INVx4_ASAP7_75t_L g12642 ( 
.A(n_11581),
.Y(n_12642)
);

INVx1_ASAP7_75t_L g12643 ( 
.A(n_11819),
.Y(n_12643)
);

INVx1_ASAP7_75t_L g12644 ( 
.A(n_11821),
.Y(n_12644)
);

BUFx2_ASAP7_75t_L g12645 ( 
.A(n_11568),
.Y(n_12645)
);

INVx1_ASAP7_75t_L g12646 ( 
.A(n_11826),
.Y(n_12646)
);

AND2x2_ASAP7_75t_L g12647 ( 
.A(n_12186),
.B(n_11960),
.Y(n_12647)
);

BUFx2_ASAP7_75t_SL g12648 ( 
.A(n_11754),
.Y(n_12648)
);

NAND2xp5_ASAP7_75t_L g12649 ( 
.A(n_11545),
.B(n_10743),
.Y(n_12649)
);

INVx2_ASAP7_75t_L g12650 ( 
.A(n_12240),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_11841),
.Y(n_12651)
);

AND2x2_ASAP7_75t_L g12652 ( 
.A(n_11713),
.B(n_9927),
.Y(n_12652)
);

INVx3_ASAP7_75t_L g12653 ( 
.A(n_12254),
.Y(n_12653)
);

OR2x2_ASAP7_75t_L g12654 ( 
.A(n_12338),
.B(n_8737),
.Y(n_12654)
);

BUFx2_ASAP7_75t_L g12655 ( 
.A(n_11954),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_11687),
.B(n_10058),
.Y(n_12656)
);

NAND2xp5_ASAP7_75t_L g12657 ( 
.A(n_11565),
.B(n_10746),
.Y(n_12657)
);

INVx3_ASAP7_75t_L g12658 ( 
.A(n_11681),
.Y(n_12658)
);

INVx2_ASAP7_75t_L g12659 ( 
.A(n_12240),
.Y(n_12659)
);

NAND2xp5_ASAP7_75t_L g12660 ( 
.A(n_11621),
.B(n_10748),
.Y(n_12660)
);

INVx1_ASAP7_75t_L g12661 ( 
.A(n_11844),
.Y(n_12661)
);

INVx1_ASAP7_75t_L g12662 ( 
.A(n_11854),
.Y(n_12662)
);

INVxp67_ASAP7_75t_SL g12663 ( 
.A(n_11576),
.Y(n_12663)
);

INVx2_ASAP7_75t_L g12664 ( 
.A(n_12268),
.Y(n_12664)
);

INVx1_ASAP7_75t_L g12665 ( 
.A(n_11863),
.Y(n_12665)
);

INVx2_ASAP7_75t_L g12666 ( 
.A(n_12268),
.Y(n_12666)
);

AND2x2_ASAP7_75t_L g12667 ( 
.A(n_11650),
.B(n_10058),
.Y(n_12667)
);

INVx1_ASAP7_75t_L g12668 ( 
.A(n_11866),
.Y(n_12668)
);

BUFx3_ASAP7_75t_L g12669 ( 
.A(n_11875),
.Y(n_12669)
);

INVx1_ASAP7_75t_L g12670 ( 
.A(n_11898),
.Y(n_12670)
);

NOR2x1_ASAP7_75t_L g12671 ( 
.A(n_11643),
.B(n_11276),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_11901),
.Y(n_12672)
);

BUFx3_ASAP7_75t_L g12673 ( 
.A(n_12120),
.Y(n_12673)
);

OAI22xp5_ASAP7_75t_L g12674 ( 
.A1(n_11543),
.A2(n_11276),
.B1(n_11347),
.B2(n_11291),
.Y(n_12674)
);

INVx2_ASAP7_75t_L g12675 ( 
.A(n_12268),
.Y(n_12675)
);

INVx1_ASAP7_75t_L g12676 ( 
.A(n_11902),
.Y(n_12676)
);

AND2x2_ASAP7_75t_L g12677 ( 
.A(n_11652),
.B(n_10061),
.Y(n_12677)
);

AND2x2_ASAP7_75t_L g12678 ( 
.A(n_11658),
.B(n_10061),
.Y(n_12678)
);

HB1xp67_ASAP7_75t_L g12679 ( 
.A(n_12342),
.Y(n_12679)
);

INVx1_ASAP7_75t_L g12680 ( 
.A(n_11920),
.Y(n_12680)
);

AND2x2_ASAP7_75t_L g12681 ( 
.A(n_11580),
.B(n_10066),
.Y(n_12681)
);

AND2x2_ASAP7_75t_L g12682 ( 
.A(n_12012),
.B(n_10066),
.Y(n_12682)
);

INVx2_ASAP7_75t_L g12683 ( 
.A(n_12426),
.Y(n_12683)
);

AND2x2_ASAP7_75t_L g12684 ( 
.A(n_12065),
.B(n_10100),
.Y(n_12684)
);

AND2x2_ASAP7_75t_L g12685 ( 
.A(n_11705),
.B(n_11706),
.Y(n_12685)
);

INVx1_ASAP7_75t_L g12686 ( 
.A(n_11936),
.Y(n_12686)
);

INVx2_ASAP7_75t_L g12687 ( 
.A(n_12426),
.Y(n_12687)
);

AND2x2_ASAP7_75t_L g12688 ( 
.A(n_11716),
.B(n_10100),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_11952),
.Y(n_12689)
);

OR2x2_ASAP7_75t_L g12690 ( 
.A(n_11544),
.B(n_8737),
.Y(n_12690)
);

INVx1_ASAP7_75t_L g12691 ( 
.A(n_11961),
.Y(n_12691)
);

INVx1_ASAP7_75t_L g12692 ( 
.A(n_11981),
.Y(n_12692)
);

AND2x2_ASAP7_75t_L g12693 ( 
.A(n_11726),
.B(n_10103),
.Y(n_12693)
);

INVx1_ASAP7_75t_L g12694 ( 
.A(n_11992),
.Y(n_12694)
);

AND2x4_ASAP7_75t_L g12695 ( 
.A(n_12244),
.B(n_11291),
.Y(n_12695)
);

AND2x2_ASAP7_75t_L g12696 ( 
.A(n_11799),
.B(n_10103),
.Y(n_12696)
);

OAI22xp5_ASAP7_75t_L g12697 ( 
.A1(n_11550),
.A2(n_11291),
.B1(n_11349),
.B2(n_11347),
.Y(n_12697)
);

INVx2_ASAP7_75t_L g12698 ( 
.A(n_12426),
.Y(n_12698)
);

INVx1_ASAP7_75t_L g12699 ( 
.A(n_11994),
.Y(n_12699)
);

INVx3_ASAP7_75t_L g12700 ( 
.A(n_12094),
.Y(n_12700)
);

AND2x2_ASAP7_75t_L g12701 ( 
.A(n_11809),
.B(n_10202),
.Y(n_12701)
);

INVx2_ASAP7_75t_L g12702 ( 
.A(n_12472),
.Y(n_12702)
);

BUFx2_ASAP7_75t_L g12703 ( 
.A(n_12122),
.Y(n_12703)
);

AND2x2_ASAP7_75t_L g12704 ( 
.A(n_11848),
.B(n_10202),
.Y(n_12704)
);

INVx4_ASAP7_75t_L g12705 ( 
.A(n_11663),
.Y(n_12705)
);

INVx1_ASAP7_75t_L g12706 ( 
.A(n_12000),
.Y(n_12706)
);

OR2x2_ASAP7_75t_L g12707 ( 
.A(n_11549),
.B(n_8737),
.Y(n_12707)
);

INVx2_ASAP7_75t_L g12708 ( 
.A(n_12472),
.Y(n_12708)
);

INVx2_ASAP7_75t_L g12709 ( 
.A(n_12472),
.Y(n_12709)
);

INVx2_ASAP7_75t_L g12710 ( 
.A(n_12500),
.Y(n_12710)
);

AND2x2_ASAP7_75t_L g12711 ( 
.A(n_11861),
.B(n_10213),
.Y(n_12711)
);

HB1xp67_ASAP7_75t_L g12712 ( 
.A(n_11624),
.Y(n_12712)
);

OR2x2_ASAP7_75t_L g12713 ( 
.A(n_11553),
.B(n_8737),
.Y(n_12713)
);

INVx1_ASAP7_75t_L g12714 ( 
.A(n_12028),
.Y(n_12714)
);

AND2x2_ASAP7_75t_L g12715 ( 
.A(n_11871),
.B(n_10213),
.Y(n_12715)
);

INVx2_ASAP7_75t_L g12716 ( 
.A(n_12500),
.Y(n_12716)
);

INVx1_ASAP7_75t_L g12717 ( 
.A(n_12032),
.Y(n_12717)
);

INVx1_ASAP7_75t_L g12718 ( 
.A(n_12036),
.Y(n_12718)
);

INVx2_ASAP7_75t_L g12719 ( 
.A(n_12500),
.Y(n_12719)
);

AND2x2_ASAP7_75t_L g12720 ( 
.A(n_11878),
.B(n_10243),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_11631),
.B(n_10752),
.Y(n_12721)
);

AND2x2_ASAP7_75t_L g12722 ( 
.A(n_11888),
.B(n_10243),
.Y(n_12722)
);

INVx1_ASAP7_75t_L g12723 ( 
.A(n_12042),
.Y(n_12723)
);

INVx2_ASAP7_75t_L g12724 ( 
.A(n_11796),
.Y(n_12724)
);

AOI22xp33_ASAP7_75t_L g12725 ( 
.A1(n_11583),
.A2(n_11349),
.B1(n_11357),
.B2(n_11347),
.Y(n_12725)
);

AND2x2_ASAP7_75t_L g12726 ( 
.A(n_11893),
.B(n_10251),
.Y(n_12726)
);

HB1xp67_ASAP7_75t_L g12727 ( 
.A(n_11656),
.Y(n_12727)
);

NAND2xp5_ASAP7_75t_L g12728 ( 
.A(n_11662),
.B(n_10753),
.Y(n_12728)
);

INVx1_ASAP7_75t_L g12729 ( 
.A(n_12051),
.Y(n_12729)
);

INVx1_ASAP7_75t_L g12730 ( 
.A(n_12052),
.Y(n_12730)
);

NAND2xp5_ASAP7_75t_L g12731 ( 
.A(n_11675),
.B(n_10754),
.Y(n_12731)
);

INVx2_ASAP7_75t_L g12732 ( 
.A(n_12357),
.Y(n_12732)
);

NOR2xp33_ASAP7_75t_L g12733 ( 
.A(n_11663),
.B(n_7469),
.Y(n_12733)
);

INVx1_ASAP7_75t_L g12734 ( 
.A(n_12055),
.Y(n_12734)
);

INVx1_ASAP7_75t_L g12735 ( 
.A(n_12095),
.Y(n_12735)
);

HB1xp67_ASAP7_75t_L g12736 ( 
.A(n_11686),
.Y(n_12736)
);

AND2x2_ASAP7_75t_L g12737 ( 
.A(n_11906),
.B(n_10251),
.Y(n_12737)
);

INVx1_ASAP7_75t_L g12738 ( 
.A(n_12117),
.Y(n_12738)
);

HB1xp67_ASAP7_75t_L g12739 ( 
.A(n_11695),
.Y(n_12739)
);

AND2x2_ASAP7_75t_L g12740 ( 
.A(n_12308),
.B(n_10269),
.Y(n_12740)
);

INVx1_ASAP7_75t_L g12741 ( 
.A(n_12133),
.Y(n_12741)
);

INVx2_ASAP7_75t_L g12742 ( 
.A(n_12357),
.Y(n_12742)
);

INVx4_ASAP7_75t_L g12743 ( 
.A(n_11663),
.Y(n_12743)
);

INVx2_ASAP7_75t_L g12744 ( 
.A(n_12518),
.Y(n_12744)
);

OR2x2_ASAP7_75t_L g12745 ( 
.A(n_11572),
.B(n_8737),
.Y(n_12745)
);

INVxp67_ASAP7_75t_SL g12746 ( 
.A(n_11803),
.Y(n_12746)
);

AND2x2_ASAP7_75t_L g12747 ( 
.A(n_12094),
.B(n_12139),
.Y(n_12747)
);

AND2x4_ASAP7_75t_L g12748 ( 
.A(n_11958),
.B(n_11349),
.Y(n_12748)
);

INVx2_ASAP7_75t_L g12749 ( 
.A(n_12518),
.Y(n_12749)
);

NOR2x1p5_ASAP7_75t_L g12750 ( 
.A(n_11551),
.B(n_7476),
.Y(n_12750)
);

NAND2xp5_ASAP7_75t_SL g12751 ( 
.A(n_11548),
.B(n_9303),
.Y(n_12751)
);

BUFx2_ASAP7_75t_L g12752 ( 
.A(n_12122),
.Y(n_12752)
);

HB1xp67_ASAP7_75t_L g12753 ( 
.A(n_11709),
.Y(n_12753)
);

NAND2xp5_ASAP7_75t_SL g12754 ( 
.A(n_11555),
.B(n_9303),
.Y(n_12754)
);

INVx2_ASAP7_75t_L g12755 ( 
.A(n_12330),
.Y(n_12755)
);

INVx1_ASAP7_75t_L g12756 ( 
.A(n_12155),
.Y(n_12756)
);

NAND2x1p5_ASAP7_75t_L g12757 ( 
.A(n_12098),
.B(n_8953),
.Y(n_12757)
);

OR2x2_ASAP7_75t_L g12758 ( 
.A(n_11573),
.B(n_8737),
.Y(n_12758)
);

CKINVDCx5p33_ASAP7_75t_R g12759 ( 
.A(n_11742),
.Y(n_12759)
);

OR2x2_ASAP7_75t_L g12760 ( 
.A(n_11598),
.B(n_8737),
.Y(n_12760)
);

BUFx3_ASAP7_75t_L g12761 ( 
.A(n_11660),
.Y(n_12761)
);

INVx1_ASAP7_75t_L g12762 ( 
.A(n_12159),
.Y(n_12762)
);

INVx1_ASAP7_75t_L g12763 ( 
.A(n_12160),
.Y(n_12763)
);

INVx2_ASAP7_75t_L g12764 ( 
.A(n_12330),
.Y(n_12764)
);

AND2x2_ASAP7_75t_L g12765 ( 
.A(n_12139),
.B(n_10269),
.Y(n_12765)
);

OR2x2_ASAP7_75t_L g12766 ( 
.A(n_11616),
.B(n_8737),
.Y(n_12766)
);

BUFx2_ASAP7_75t_L g12767 ( 
.A(n_12122),
.Y(n_12767)
);

INVx1_ASAP7_75t_L g12768 ( 
.A(n_12165),
.Y(n_12768)
);

NOR2xp33_ASAP7_75t_L g12769 ( 
.A(n_11660),
.B(n_7439),
.Y(n_12769)
);

INVx1_ASAP7_75t_L g12770 ( 
.A(n_12182),
.Y(n_12770)
);

AND2x2_ASAP7_75t_L g12771 ( 
.A(n_12174),
.B(n_10308),
.Y(n_12771)
);

BUFx3_ASAP7_75t_L g12772 ( 
.A(n_11676),
.Y(n_12772)
);

HB1xp67_ASAP7_75t_L g12773 ( 
.A(n_11748),
.Y(n_12773)
);

INVx1_ASAP7_75t_L g12774 ( 
.A(n_12187),
.Y(n_12774)
);

INVx1_ASAP7_75t_L g12775 ( 
.A(n_12189),
.Y(n_12775)
);

INVx1_ASAP7_75t_L g12776 ( 
.A(n_12192),
.Y(n_12776)
);

AND2x2_ASAP7_75t_L g12777 ( 
.A(n_12174),
.B(n_10308),
.Y(n_12777)
);

AND2x2_ASAP7_75t_L g12778 ( 
.A(n_11946),
.B(n_9921),
.Y(n_12778)
);

INVx1_ASAP7_75t_L g12779 ( 
.A(n_12195),
.Y(n_12779)
);

AND2x4_ASAP7_75t_L g12780 ( 
.A(n_11958),
.B(n_11357),
.Y(n_12780)
);

HB1xp67_ASAP7_75t_L g12781 ( 
.A(n_11770),
.Y(n_12781)
);

INVx2_ASAP7_75t_L g12782 ( 
.A(n_12348),
.Y(n_12782)
);

INVx1_ASAP7_75t_L g12783 ( 
.A(n_12199),
.Y(n_12783)
);

AND2x2_ASAP7_75t_L g12784 ( 
.A(n_11950),
.B(n_11357),
.Y(n_12784)
);

HB1xp67_ASAP7_75t_L g12785 ( 
.A(n_11629),
.Y(n_12785)
);

INVx2_ASAP7_75t_L g12786 ( 
.A(n_12348),
.Y(n_12786)
);

INVx2_ASAP7_75t_L g12787 ( 
.A(n_12351),
.Y(n_12787)
);

HB1xp67_ASAP7_75t_L g12788 ( 
.A(n_11633),
.Y(n_12788)
);

NAND2xp5_ASAP7_75t_L g12789 ( 
.A(n_11597),
.B(n_10758),
.Y(n_12789)
);

OR2x2_ASAP7_75t_L g12790 ( 
.A(n_11641),
.B(n_10759),
.Y(n_12790)
);

INVx1_ASAP7_75t_L g12791 ( 
.A(n_12208),
.Y(n_12791)
);

AND2x4_ASAP7_75t_L g12792 ( 
.A(n_12191),
.B(n_11423),
.Y(n_12792)
);

INVx2_ASAP7_75t_L g12793 ( 
.A(n_12351),
.Y(n_12793)
);

INVx2_ASAP7_75t_SL g12794 ( 
.A(n_11766),
.Y(n_12794)
);

INVx2_ASAP7_75t_L g12795 ( 
.A(n_12371),
.Y(n_12795)
);

INVx2_ASAP7_75t_L g12796 ( 
.A(n_12377),
.Y(n_12796)
);

BUFx3_ASAP7_75t_L g12797 ( 
.A(n_11676),
.Y(n_12797)
);

INVx1_ASAP7_75t_L g12798 ( 
.A(n_12210),
.Y(n_12798)
);

INVx1_ASAP7_75t_L g12799 ( 
.A(n_12211),
.Y(n_12799)
);

AND2x4_ASAP7_75t_L g12800 ( 
.A(n_11941),
.B(n_11423),
.Y(n_12800)
);

BUFx2_ASAP7_75t_L g12801 ( 
.A(n_12122),
.Y(n_12801)
);

INVx2_ASAP7_75t_L g12802 ( 
.A(n_12453),
.Y(n_12802)
);

AND2x4_ASAP7_75t_L g12803 ( 
.A(n_11941),
.B(n_11423),
.Y(n_12803)
);

OR2x2_ASAP7_75t_L g12804 ( 
.A(n_11665),
.B(n_10763),
.Y(n_12804)
);

OR2x2_ASAP7_75t_L g12805 ( 
.A(n_11626),
.B(n_10773),
.Y(n_12805)
);

BUFx2_ASAP7_75t_L g12806 ( 
.A(n_12386),
.Y(n_12806)
);

NOR2xp33_ASAP7_75t_SL g12807 ( 
.A(n_12061),
.B(n_7383),
.Y(n_12807)
);

INVx3_ASAP7_75t_L g12808 ( 
.A(n_12218),
.Y(n_12808)
);

NAND2xp5_ASAP7_75t_L g12809 ( 
.A(n_11645),
.B(n_10774),
.Y(n_12809)
);

INVx2_ASAP7_75t_L g12810 ( 
.A(n_12482),
.Y(n_12810)
);

INVx1_ASAP7_75t_L g12811 ( 
.A(n_12213),
.Y(n_12811)
);

HB1xp67_ASAP7_75t_L g12812 ( 
.A(n_12461),
.Y(n_12812)
);

BUFx2_ASAP7_75t_L g12813 ( 
.A(n_12198),
.Y(n_12813)
);

HB1xp67_ASAP7_75t_L g12814 ( 
.A(n_12496),
.Y(n_12814)
);

INVx2_ASAP7_75t_L g12815 ( 
.A(n_12482),
.Y(n_12815)
);

AND2x2_ASAP7_75t_L g12816 ( 
.A(n_11651),
.B(n_11460),
.Y(n_12816)
);

INVx1_ASAP7_75t_L g12817 ( 
.A(n_12214),
.Y(n_12817)
);

OR2x2_ASAP7_75t_L g12818 ( 
.A(n_11601),
.B(n_10776),
.Y(n_12818)
);

OR2x2_ASAP7_75t_L g12819 ( 
.A(n_11661),
.B(n_10778),
.Y(n_12819)
);

HB1xp67_ASAP7_75t_L g12820 ( 
.A(n_11944),
.Y(n_12820)
);

INVx1_ASAP7_75t_L g12821 ( 
.A(n_12222),
.Y(n_12821)
);

AND2x2_ASAP7_75t_L g12822 ( 
.A(n_12108),
.B(n_11460),
.Y(n_12822)
);

AOI22xp33_ASAP7_75t_SL g12823 ( 
.A1(n_11594),
.A2(n_8015),
.B1(n_11464),
.B2(n_11460),
.Y(n_12823)
);

AOI22xp33_ASAP7_75t_L g12824 ( 
.A1(n_11578),
.A2(n_11538),
.B1(n_11464),
.B2(n_9752),
.Y(n_12824)
);

AND2x2_ASAP7_75t_L g12825 ( 
.A(n_11955),
.B(n_11464),
.Y(n_12825)
);

INVx1_ASAP7_75t_L g12826 ( 
.A(n_12248),
.Y(n_12826)
);

INVx5_ASAP7_75t_L g12827 ( 
.A(n_11618),
.Y(n_12827)
);

OR2x2_ASAP7_75t_L g12828 ( 
.A(n_11968),
.B(n_10782),
.Y(n_12828)
);

INVx1_ASAP7_75t_L g12829 ( 
.A(n_12278),
.Y(n_12829)
);

AND2x2_ASAP7_75t_L g12830 ( 
.A(n_11988),
.B(n_11762),
.Y(n_12830)
);

INVx1_ASAP7_75t_L g12831 ( 
.A(n_12320),
.Y(n_12831)
);

AOI21xp33_ASAP7_75t_L g12832 ( 
.A1(n_11635),
.A2(n_9752),
.B(n_9730),
.Y(n_12832)
);

INVx2_ASAP7_75t_SL g12833 ( 
.A(n_12236),
.Y(n_12833)
);

AND2x2_ASAP7_75t_L g12834 ( 
.A(n_11825),
.B(n_11538),
.Y(n_12834)
);

AND2x2_ASAP7_75t_L g12835 ( 
.A(n_11730),
.B(n_11538),
.Y(n_12835)
);

INVx2_ASAP7_75t_L g12836 ( 
.A(n_11998),
.Y(n_12836)
);

AOI22xp33_ASAP7_75t_L g12837 ( 
.A1(n_11563),
.A2(n_9752),
.B1(n_9754),
.B2(n_9730),
.Y(n_12837)
);

HB1xp67_ASAP7_75t_L g12838 ( 
.A(n_11758),
.Y(n_12838)
);

INVx2_ASAP7_75t_L g12839 ( 
.A(n_12066),
.Y(n_12839)
);

NAND2xp5_ASAP7_75t_L g12840 ( 
.A(n_11596),
.B(n_10783),
.Y(n_12840)
);

INVx2_ASAP7_75t_SL g12841 ( 
.A(n_11773),
.Y(n_12841)
);

AND2x2_ASAP7_75t_L g12842 ( 
.A(n_11817),
.B(n_10154),
.Y(n_12842)
);

INVx2_ASAP7_75t_L g12843 ( 
.A(n_11758),
.Y(n_12843)
);

INVxp67_ASAP7_75t_SL g12844 ( 
.A(n_12018),
.Y(n_12844)
);

AND2x4_ASAP7_75t_L g12845 ( 
.A(n_12164),
.B(n_10711),
.Y(n_12845)
);

INVx1_ASAP7_75t_L g12846 ( 
.A(n_12326),
.Y(n_12846)
);

INVx2_ASAP7_75t_L g12847 ( 
.A(n_11758),
.Y(n_12847)
);

INVx2_ASAP7_75t_SL g12848 ( 
.A(n_12097),
.Y(n_12848)
);

BUFx2_ASAP7_75t_L g12849 ( 
.A(n_12217),
.Y(n_12849)
);

INVx1_ASAP7_75t_L g12850 ( 
.A(n_12339),
.Y(n_12850)
);

NAND2xp5_ASAP7_75t_L g12851 ( 
.A(n_11591),
.B(n_10788),
.Y(n_12851)
);

OR2x2_ASAP7_75t_L g12852 ( 
.A(n_12420),
.B(n_10789),
.Y(n_12852)
);

BUFx2_ASAP7_75t_L g12853 ( 
.A(n_12181),
.Y(n_12853)
);

AND2x2_ASAP7_75t_L g12854 ( 
.A(n_12075),
.B(n_10154),
.Y(n_12854)
);

HB1xp67_ASAP7_75t_L g12855 ( 
.A(n_11856),
.Y(n_12855)
);

AND2x2_ASAP7_75t_L g12856 ( 
.A(n_12075),
.B(n_10216),
.Y(n_12856)
);

NOR2xp33_ASAP7_75t_L g12857 ( 
.A(n_11649),
.B(n_7452),
.Y(n_12857)
);

AND2x2_ASAP7_75t_L g12858 ( 
.A(n_12400),
.B(n_10216),
.Y(n_12858)
);

AND2x2_ASAP7_75t_L g12859 ( 
.A(n_12419),
.B(n_10255),
.Y(n_12859)
);

NAND2xp5_ASAP7_75t_L g12860 ( 
.A(n_11592),
.B(n_10800),
.Y(n_12860)
);

INVx1_ASAP7_75t_L g12861 ( 
.A(n_12350),
.Y(n_12861)
);

INVxp67_ASAP7_75t_SL g12862 ( 
.A(n_12291),
.Y(n_12862)
);

INVx2_ASAP7_75t_L g12863 ( 
.A(n_11856),
.Y(n_12863)
);

AND2x4_ASAP7_75t_SL g12864 ( 
.A(n_11872),
.B(n_7732),
.Y(n_12864)
);

INVx1_ASAP7_75t_L g12865 ( 
.A(n_12353),
.Y(n_12865)
);

NAND2xp5_ASAP7_75t_L g12866 ( 
.A(n_11599),
.B(n_10801),
.Y(n_12866)
);

INVx2_ASAP7_75t_L g12867 ( 
.A(n_11856),
.Y(n_12867)
);

INVx1_ASAP7_75t_SL g12868 ( 
.A(n_12234),
.Y(n_12868)
);

INVx3_ASAP7_75t_L g12869 ( 
.A(n_12488),
.Y(n_12869)
);

AND2x2_ASAP7_75t_L g12870 ( 
.A(n_12451),
.B(n_10255),
.Y(n_12870)
);

INVx1_ASAP7_75t_L g12871 ( 
.A(n_12356),
.Y(n_12871)
);

AND2x2_ASAP7_75t_L g12872 ( 
.A(n_11999),
.B(n_10255),
.Y(n_12872)
);

INVx1_ASAP7_75t_L g12873 ( 
.A(n_12359),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_12363),
.Y(n_12874)
);

NAND2xp5_ASAP7_75t_L g12875 ( 
.A(n_11584),
.B(n_10804),
.Y(n_12875)
);

INVx1_ASAP7_75t_L g12876 ( 
.A(n_12375),
.Y(n_12876)
);

OR2x2_ASAP7_75t_L g12877 ( 
.A(n_12480),
.B(n_10807),
.Y(n_12877)
);

NAND2xp5_ASAP7_75t_L g12878 ( 
.A(n_11775),
.B(n_10810),
.Y(n_12878)
);

AND2x2_ASAP7_75t_L g12879 ( 
.A(n_12003),
.B(n_10303),
.Y(n_12879)
);

INVx1_ASAP7_75t_L g12880 ( 
.A(n_12384),
.Y(n_12880)
);

INVx1_ASAP7_75t_L g12881 ( 
.A(n_12390),
.Y(n_12881)
);

INVx1_ASAP7_75t_L g12882 ( 
.A(n_12391),
.Y(n_12882)
);

NAND2xp5_ASAP7_75t_L g12883 ( 
.A(n_11783),
.B(n_10812),
.Y(n_12883)
);

INVx2_ASAP7_75t_SL g12884 ( 
.A(n_12097),
.Y(n_12884)
);

INVx2_ASAP7_75t_L g12885 ( 
.A(n_12004),
.Y(n_12885)
);

AND2x2_ASAP7_75t_L g12886 ( 
.A(n_12258),
.B(n_10303),
.Y(n_12886)
);

OR2x2_ASAP7_75t_L g12887 ( 
.A(n_11769),
.B(n_10814),
.Y(n_12887)
);

AND2x2_ASAP7_75t_L g12888 ( 
.A(n_12276),
.B(n_10303),
.Y(n_12888)
);

AND2x2_ASAP7_75t_L g12889 ( 
.A(n_12300),
.B(n_10303),
.Y(n_12889)
);

INVx1_ASAP7_75t_L g12890 ( 
.A(n_12407),
.Y(n_12890)
);

INVxp67_ASAP7_75t_L g12891 ( 
.A(n_12349),
.Y(n_12891)
);

AND2x2_ASAP7_75t_L g12892 ( 
.A(n_12315),
.B(n_10313),
.Y(n_12892)
);

INVx1_ASAP7_75t_L g12893 ( 
.A(n_12408),
.Y(n_12893)
);

AND2x2_ASAP7_75t_L g12894 ( 
.A(n_12166),
.B(n_10313),
.Y(n_12894)
);

AND2x4_ASAP7_75t_L g12895 ( 
.A(n_11779),
.B(n_10711),
.Y(n_12895)
);

INVx2_ASAP7_75t_L g12896 ( 
.A(n_12004),
.Y(n_12896)
);

AND2x2_ASAP7_75t_L g12897 ( 
.A(n_12341),
.B(n_12381),
.Y(n_12897)
);

NAND2xp5_ASAP7_75t_L g12898 ( 
.A(n_11586),
.B(n_11588),
.Y(n_12898)
);

INVxp67_ASAP7_75t_L g12899 ( 
.A(n_12404),
.Y(n_12899)
);

INVx2_ASAP7_75t_L g12900 ( 
.A(n_12004),
.Y(n_12900)
);

AND2x2_ASAP7_75t_L g12901 ( 
.A(n_11642),
.B(n_10313),
.Y(n_12901)
);

INVx2_ASAP7_75t_L g12902 ( 
.A(n_12053),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_12412),
.Y(n_12903)
);

AND2x2_ASAP7_75t_L g12904 ( 
.A(n_12054),
.B(n_10313),
.Y(n_12904)
);

AND2x2_ASAP7_75t_L g12905 ( 
.A(n_12101),
.B(n_10333),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_12414),
.Y(n_12906)
);

OR2x2_ASAP7_75t_L g12907 ( 
.A(n_12360),
.B(n_10818),
.Y(n_12907)
);

INVx1_ASAP7_75t_L g12908 ( 
.A(n_12434),
.Y(n_12908)
);

OR2x2_ASAP7_75t_L g12909 ( 
.A(n_11688),
.B(n_10819),
.Y(n_12909)
);

BUFx3_ASAP7_75t_L g12910 ( 
.A(n_11831),
.Y(n_12910)
);

INVx3_ASAP7_75t_L g12911 ( 
.A(n_12488),
.Y(n_12911)
);

INVxp67_ASAP7_75t_L g12912 ( 
.A(n_12053),
.Y(n_12912)
);

HB1xp67_ASAP7_75t_L g12913 ( 
.A(n_12053),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_12435),
.Y(n_12914)
);

HB1xp67_ASAP7_75t_L g12915 ( 
.A(n_12197),
.Y(n_12915)
);

AND2x2_ASAP7_75t_L g12916 ( 
.A(n_12074),
.B(n_10333),
.Y(n_12916)
);

AND2x4_ASAP7_75t_L g12917 ( 
.A(n_11779),
.B(n_10333),
.Y(n_12917)
);

INVx2_ASAP7_75t_L g12918 ( 
.A(n_12207),
.Y(n_12918)
);

OR2x2_ASAP7_75t_L g12919 ( 
.A(n_11702),
.B(n_10820),
.Y(n_12919)
);

HB1xp67_ASAP7_75t_L g12920 ( 
.A(n_12373),
.Y(n_12920)
);

AND2x2_ASAP7_75t_L g12921 ( 
.A(n_12237),
.B(n_10333),
.Y(n_12921)
);

AND2x2_ASAP7_75t_L g12922 ( 
.A(n_11753),
.B(n_8375),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12449),
.Y(n_12923)
);

BUFx2_ASAP7_75t_L g12924 ( 
.A(n_11872),
.Y(n_12924)
);

AND2x2_ASAP7_75t_L g12925 ( 
.A(n_11757),
.B(n_8377),
.Y(n_12925)
);

INVx2_ASAP7_75t_L g12926 ( 
.A(n_12132),
.Y(n_12926)
);

INVx2_ASAP7_75t_L g12927 ( 
.A(n_12430),
.Y(n_12927)
);

INVx2_ASAP7_75t_L g12928 ( 
.A(n_12460),
.Y(n_12928)
);

AND2x2_ASAP7_75t_L g12929 ( 
.A(n_12109),
.B(n_8377),
.Y(n_12929)
);

AND2x2_ASAP7_75t_L g12930 ( 
.A(n_12148),
.B(n_8391),
.Y(n_12930)
);

AOI22xp33_ASAP7_75t_L g12931 ( 
.A1(n_11560),
.A2(n_9752),
.B1(n_9754),
.B2(n_9730),
.Y(n_12931)
);

BUFx6f_ASAP7_75t_L g12932 ( 
.A(n_12113),
.Y(n_12932)
);

AND2x2_ASAP7_75t_L g12933 ( 
.A(n_12152),
.B(n_8391),
.Y(n_12933)
);

BUFx2_ASAP7_75t_L g12934 ( 
.A(n_12327),
.Y(n_12934)
);

AND2x2_ASAP7_75t_L g12935 ( 
.A(n_11760),
.B(n_8391),
.Y(n_12935)
);

INVxp67_ASAP7_75t_L g12936 ( 
.A(n_12157),
.Y(n_12936)
);

INVx2_ASAP7_75t_L g12937 ( 
.A(n_11980),
.Y(n_12937)
);

INVx1_ASAP7_75t_L g12938 ( 
.A(n_12454),
.Y(n_12938)
);

NAND2xp5_ASAP7_75t_L g12939 ( 
.A(n_11564),
.B(n_10821),
.Y(n_12939)
);

AND2x2_ASAP7_75t_L g12940 ( 
.A(n_12171),
.B(n_8393),
.Y(n_12940)
);

INVx3_ASAP7_75t_SL g12941 ( 
.A(n_12115),
.Y(n_12941)
);

INVx1_ASAP7_75t_L g12942 ( 
.A(n_12458),
.Y(n_12942)
);

INVx2_ASAP7_75t_L g12943 ( 
.A(n_11980),
.Y(n_12943)
);

NAND2xp5_ASAP7_75t_L g12944 ( 
.A(n_11605),
.B(n_10822),
.Y(n_12944)
);

OR2x2_ASAP7_75t_L g12945 ( 
.A(n_11786),
.B(n_10842),
.Y(n_12945)
);

INVx1_ASAP7_75t_SL g12946 ( 
.A(n_12443),
.Y(n_12946)
);

BUFx3_ASAP7_75t_L g12947 ( 
.A(n_11664),
.Y(n_12947)
);

NAND2xp5_ASAP7_75t_L g12948 ( 
.A(n_11585),
.B(n_10850),
.Y(n_12948)
);

INVx3_ASAP7_75t_L g12949 ( 
.A(n_11834),
.Y(n_12949)
);

INVx2_ASAP7_75t_L g12950 ( 
.A(n_12013),
.Y(n_12950)
);

INVx2_ASAP7_75t_L g12951 ( 
.A(n_12013),
.Y(n_12951)
);

INVx1_ASAP7_75t_L g12952 ( 
.A(n_12462),
.Y(n_12952)
);

INVx2_ASAP7_75t_L g12953 ( 
.A(n_12025),
.Y(n_12953)
);

HB1xp67_ASAP7_75t_L g12954 ( 
.A(n_12425),
.Y(n_12954)
);

AND2x2_ASAP7_75t_L g12955 ( 
.A(n_12176),
.B(n_8393),
.Y(n_12955)
);

INVx2_ASAP7_75t_L g12956 ( 
.A(n_12025),
.Y(n_12956)
);

OR2x2_ASAP7_75t_L g12957 ( 
.A(n_11800),
.B(n_10866),
.Y(n_12957)
);

BUFx2_ASAP7_75t_L g12958 ( 
.A(n_12331),
.Y(n_12958)
);

INVx3_ASAP7_75t_L g12959 ( 
.A(n_11834),
.Y(n_12959)
);

INVx2_ASAP7_75t_L g12960 ( 
.A(n_12089),
.Y(n_12960)
);

AND2x2_ASAP7_75t_L g12961 ( 
.A(n_12178),
.B(n_8393),
.Y(n_12961)
);

INVx2_ASAP7_75t_L g12962 ( 
.A(n_12089),
.Y(n_12962)
);

AND2x2_ASAP7_75t_L g12963 ( 
.A(n_12179),
.B(n_8395),
.Y(n_12963)
);

AND2x2_ASAP7_75t_L g12964 ( 
.A(n_12183),
.B(n_8395),
.Y(n_12964)
);

AND2x2_ASAP7_75t_L g12965 ( 
.A(n_12184),
.B(n_8395),
.Y(n_12965)
);

INVx1_ASAP7_75t_L g12966 ( 
.A(n_12474),
.Y(n_12966)
);

INVx1_ASAP7_75t_L g12967 ( 
.A(n_12484),
.Y(n_12967)
);

BUFx3_ASAP7_75t_L g12968 ( 
.A(n_11679),
.Y(n_12968)
);

HB1xp67_ASAP7_75t_L g12969 ( 
.A(n_11620),
.Y(n_12969)
);

INVx2_ASAP7_75t_L g12970 ( 
.A(n_12105),
.Y(n_12970)
);

INVx1_ASAP7_75t_L g12971 ( 
.A(n_12495),
.Y(n_12971)
);

INVx1_ASAP7_75t_L g12972 ( 
.A(n_12499),
.Y(n_12972)
);

AND2x2_ASAP7_75t_L g12973 ( 
.A(n_12188),
.B(n_11806),
.Y(n_12973)
);

INVx1_ASAP7_75t_L g12974 ( 
.A(n_12501),
.Y(n_12974)
);

INVx2_ASAP7_75t_L g12975 ( 
.A(n_12105),
.Y(n_12975)
);

NOR2x1_ASAP7_75t_L g12976 ( 
.A(n_11671),
.B(n_10867),
.Y(n_12976)
);

NAND2xp5_ASAP7_75t_L g12977 ( 
.A(n_11755),
.B(n_10868),
.Y(n_12977)
);

AND2x2_ASAP7_75t_L g12978 ( 
.A(n_12497),
.B(n_8451),
.Y(n_12978)
);

INVx1_ASAP7_75t_L g12979 ( 
.A(n_12503),
.Y(n_12979)
);

AND2x2_ASAP7_75t_L g12980 ( 
.A(n_12515),
.B(n_8451),
.Y(n_12980)
);

INVx2_ASAP7_75t_L g12981 ( 
.A(n_11823),
.Y(n_12981)
);

INVx2_ASAP7_75t_L g12982 ( 
.A(n_11858),
.Y(n_12982)
);

AND2x4_ASAP7_75t_L g12983 ( 
.A(n_11977),
.B(n_10871),
.Y(n_12983)
);

INVx1_ASAP7_75t_L g12984 ( 
.A(n_12512),
.Y(n_12984)
);

AND2x2_ASAP7_75t_L g12985 ( 
.A(n_11795),
.B(n_8451),
.Y(n_12985)
);

INVx2_ASAP7_75t_L g12986 ( 
.A(n_11860),
.Y(n_12986)
);

HB1xp67_ASAP7_75t_L g12987 ( 
.A(n_11620),
.Y(n_12987)
);

AND2x2_ASAP7_75t_L g12988 ( 
.A(n_11805),
.B(n_12141),
.Y(n_12988)
);

BUFx2_ASAP7_75t_SL g12989 ( 
.A(n_11977),
.Y(n_12989)
);

AND2x2_ASAP7_75t_L g12990 ( 
.A(n_12146),
.B(n_8477),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_12516),
.Y(n_12991)
);

OR2x2_ASAP7_75t_L g12992 ( 
.A(n_11881),
.B(n_10873),
.Y(n_12992)
);

INVx1_ASAP7_75t_L g12993 ( 
.A(n_12511),
.Y(n_12993)
);

AND2x2_ASAP7_75t_L g12994 ( 
.A(n_11781),
.B(n_8477),
.Y(n_12994)
);

INVx2_ASAP7_75t_L g12995 ( 
.A(n_11909),
.Y(n_12995)
);

INVx2_ASAP7_75t_L g12996 ( 
.A(n_11921),
.Y(n_12996)
);

NAND2xp5_ASAP7_75t_L g12997 ( 
.A(n_11600),
.B(n_10875),
.Y(n_12997)
);

INVx4_ASAP7_75t_L g12998 ( 
.A(n_12098),
.Y(n_12998)
);

INVx2_ASAP7_75t_L g12999 ( 
.A(n_11932),
.Y(n_12999)
);

AND2x2_ASAP7_75t_L g13000 ( 
.A(n_11736),
.B(n_8477),
.Y(n_13000)
);

INVx2_ASAP7_75t_SL g13001 ( 
.A(n_11947),
.Y(n_13001)
);

NAND2xp5_ASAP7_75t_L g13002 ( 
.A(n_11556),
.B(n_10884),
.Y(n_13002)
);

AND2x2_ASAP7_75t_L g13003 ( 
.A(n_11740),
.B(n_8486),
.Y(n_13003)
);

INVx3_ASAP7_75t_L g13004 ( 
.A(n_11807),
.Y(n_13004)
);

AND2x4_ASAP7_75t_L g13005 ( 
.A(n_11764),
.B(n_10890),
.Y(n_13005)
);

INVx2_ASAP7_75t_L g13006 ( 
.A(n_11959),
.Y(n_13006)
);

INVx2_ASAP7_75t_L g13007 ( 
.A(n_12048),
.Y(n_13007)
);

INVx1_ASAP7_75t_L g13008 ( 
.A(n_12491),
.Y(n_13008)
);

HB1xp67_ASAP7_75t_L g13009 ( 
.A(n_12068),
.Y(n_13009)
);

INVx2_ASAP7_75t_L g13010 ( 
.A(n_12083),
.Y(n_13010)
);

INVx1_ASAP7_75t_L g13011 ( 
.A(n_12493),
.Y(n_13011)
);

INVx1_ASAP7_75t_L g13012 ( 
.A(n_12493),
.Y(n_13012)
);

OR2x2_ASAP7_75t_L g13013 ( 
.A(n_11659),
.B(n_10894),
.Y(n_13013)
);

AND2x2_ASAP7_75t_L g13014 ( 
.A(n_12150),
.B(n_8486),
.Y(n_13014)
);

BUFx3_ASAP7_75t_L g13015 ( 
.A(n_11692),
.Y(n_13015)
);

INVx2_ASAP7_75t_L g13016 ( 
.A(n_12084),
.Y(n_13016)
);

AND2x2_ASAP7_75t_L g13017 ( 
.A(n_12242),
.B(n_8486),
.Y(n_13017)
);

AND2x2_ASAP7_75t_L g13018 ( 
.A(n_12167),
.B(n_8503),
.Y(n_13018)
);

AND2x2_ASAP7_75t_L g13019 ( 
.A(n_11827),
.B(n_8503),
.Y(n_13019)
);

INVx2_ASAP7_75t_L g13020 ( 
.A(n_12125),
.Y(n_13020)
);

AOI222xp33_ASAP7_75t_L g13021 ( 
.A1(n_11674),
.A2(n_11547),
.B1(n_11608),
.B2(n_11562),
.C1(n_11647),
.C2(n_11571),
.Y(n_13021)
);

AND2x4_ASAP7_75t_L g13022 ( 
.A(n_11764),
.B(n_10895),
.Y(n_13022)
);

HB1xp67_ASAP7_75t_L g13023 ( 
.A(n_12129),
.Y(n_13023)
);

AND2x4_ASAP7_75t_L g13024 ( 
.A(n_11764),
.B(n_10897),
.Y(n_13024)
);

INVx1_ASAP7_75t_L g13025 ( 
.A(n_12493),
.Y(n_13025)
);

OR2x2_ASAP7_75t_L g13026 ( 
.A(n_11746),
.B(n_10907),
.Y(n_13026)
);

INVx1_ASAP7_75t_L g13027 ( 
.A(n_12138),
.Y(n_13027)
);

INVx2_ASAP7_75t_L g13028 ( 
.A(n_12228),
.Y(n_13028)
);

OR2x2_ASAP7_75t_L g13029 ( 
.A(n_11911),
.B(n_12050),
.Y(n_13029)
);

BUFx2_ASAP7_75t_L g13030 ( 
.A(n_12492),
.Y(n_13030)
);

CKINVDCx20_ASAP7_75t_R g13031 ( 
.A(n_12318),
.Y(n_13031)
);

INVxp67_ASAP7_75t_L g13032 ( 
.A(n_11617),
.Y(n_13032)
);

AND2x2_ASAP7_75t_L g13033 ( 
.A(n_11830),
.B(n_8503),
.Y(n_13033)
);

INVx1_ASAP7_75t_L g13034 ( 
.A(n_12251),
.Y(n_13034)
);

HB1xp67_ASAP7_75t_L g13035 ( 
.A(n_12274),
.Y(n_13035)
);

AND2x4_ASAP7_75t_L g13036 ( 
.A(n_12047),
.B(n_10908),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12284),
.Y(n_13037)
);

AND2x2_ASAP7_75t_L g13038 ( 
.A(n_11776),
.B(n_8509),
.Y(n_13038)
);

AND2x2_ASAP7_75t_L g13039 ( 
.A(n_11733),
.B(n_11880),
.Y(n_13039)
);

AND2x2_ASAP7_75t_L g13040 ( 
.A(n_12221),
.B(n_8509),
.Y(n_13040)
);

INVx3_ASAP7_75t_L g13041 ( 
.A(n_11899),
.Y(n_13041)
);

BUFx2_ASAP7_75t_L g13042 ( 
.A(n_11947),
.Y(n_13042)
);

AND2x2_ASAP7_75t_L g13043 ( 
.A(n_12252),
.B(n_11991),
.Y(n_13043)
);

INVx1_ASAP7_75t_L g13044 ( 
.A(n_12324),
.Y(n_13044)
);

INVx2_ASAP7_75t_L g13045 ( 
.A(n_12334),
.Y(n_13045)
);

INVx1_ASAP7_75t_L g13046 ( 
.A(n_12369),
.Y(n_13046)
);

AND2x2_ASAP7_75t_L g13047 ( 
.A(n_11993),
.B(n_8509),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_12376),
.Y(n_13048)
);

BUFx12f_ASAP7_75t_L g13049 ( 
.A(n_12450),
.Y(n_13049)
);

BUFx2_ASAP7_75t_L g13050 ( 
.A(n_11947),
.Y(n_13050)
);

INVx2_ASAP7_75t_L g13051 ( 
.A(n_12382),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12402),
.Y(n_13052)
);

INVx3_ASAP7_75t_L g13053 ( 
.A(n_11899),
.Y(n_13053)
);

INVx1_ASAP7_75t_L g13054 ( 
.A(n_12421),
.Y(n_13054)
);

AND2x2_ASAP7_75t_L g13055 ( 
.A(n_12006),
.B(n_8547),
.Y(n_13055)
);

NAND2xp5_ASAP7_75t_L g13056 ( 
.A(n_11577),
.B(n_10911),
.Y(n_13056)
);

INVx1_ASAP7_75t_L g13057 ( 
.A(n_12422),
.Y(n_13057)
);

CKINVDCx5p33_ASAP7_75t_R g13058 ( 
.A(n_11966),
.Y(n_13058)
);

INVx1_ASAP7_75t_L g13059 ( 
.A(n_12216),
.Y(n_13059)
);

AND2x2_ASAP7_75t_L g13060 ( 
.A(n_11870),
.B(n_8547),
.Y(n_13060)
);

INVx2_ASAP7_75t_L g13061 ( 
.A(n_12423),
.Y(n_13061)
);

AND2x2_ASAP7_75t_L g13062 ( 
.A(n_11914),
.B(n_8547),
.Y(n_13062)
);

INVx1_ASAP7_75t_L g13063 ( 
.A(n_12216),
.Y(n_13063)
);

BUFx3_ASAP7_75t_L g13064 ( 
.A(n_12149),
.Y(n_13064)
);

AND2x2_ASAP7_75t_L g13065 ( 
.A(n_11917),
.B(n_8626),
.Y(n_13065)
);

BUFx6f_ASAP7_75t_L g13066 ( 
.A(n_12470),
.Y(n_13066)
);

INVx2_ASAP7_75t_L g13067 ( 
.A(n_12431),
.Y(n_13067)
);

HB1xp67_ASAP7_75t_L g13068 ( 
.A(n_12485),
.Y(n_13068)
);

INVx2_ASAP7_75t_L g13069 ( 
.A(n_11684),
.Y(n_13069)
);

INVx3_ASAP7_75t_L g13070 ( 
.A(n_11684),
.Y(n_13070)
);

INVx1_ASAP7_75t_L g13071 ( 
.A(n_12216),
.Y(n_13071)
);

INVxp67_ASAP7_75t_L g13072 ( 
.A(n_11623),
.Y(n_13072)
);

AND2x4_ASAP7_75t_L g13073 ( 
.A(n_12020),
.B(n_10912),
.Y(n_13073)
);

NOR2x1_ASAP7_75t_L g13074 ( 
.A(n_11737),
.B(n_10916),
.Y(n_13074)
);

INVx1_ASAP7_75t_L g13075 ( 
.A(n_12255),
.Y(n_13075)
);

INVx4_ASAP7_75t_L g13076 ( 
.A(n_11759),
.Y(n_13076)
);

AND2x4_ASAP7_75t_SL g13077 ( 
.A(n_11785),
.B(n_7732),
.Y(n_13077)
);

AND2x2_ASAP7_75t_L g13078 ( 
.A(n_11922),
.B(n_8626),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12255),
.Y(n_13079)
);

AND2x2_ASAP7_75t_L g13080 ( 
.A(n_11923),
.B(n_8626),
.Y(n_13080)
);

AND2x2_ASAP7_75t_L g13081 ( 
.A(n_11926),
.B(n_8715),
.Y(n_13081)
);

INVx2_ASAP7_75t_L g13082 ( 
.A(n_11759),
.Y(n_13082)
);

AND2x2_ASAP7_75t_L g13083 ( 
.A(n_11928),
.B(n_11929),
.Y(n_13083)
);

INVx2_ASAP7_75t_L g13084 ( 
.A(n_11840),
.Y(n_13084)
);

BUFx8_ASAP7_75t_SL g13085 ( 
.A(n_11840),
.Y(n_13085)
);

BUFx6f_ASAP7_75t_L g13086 ( 
.A(n_11850),
.Y(n_13086)
);

AND2x4_ASAP7_75t_L g13087 ( 
.A(n_11672),
.B(n_10918),
.Y(n_13087)
);

AOI22xp5_ASAP7_75t_SL g13088 ( 
.A1(n_11615),
.A2(n_7452),
.B1(n_7555),
.B2(n_7551),
.Y(n_13088)
);

OR2x2_ASAP7_75t_L g13089 ( 
.A(n_11849),
.B(n_10922),
.Y(n_13089)
);

BUFx2_ASAP7_75t_L g13090 ( 
.A(n_12439),
.Y(n_13090)
);

AND2x2_ASAP7_75t_L g13091 ( 
.A(n_11938),
.B(n_8715),
.Y(n_13091)
);

INVx1_ASAP7_75t_L g13092 ( 
.A(n_12264),
.Y(n_13092)
);

INVx2_ASAP7_75t_L g13093 ( 
.A(n_11850),
.Y(n_13093)
);

OR2x2_ASAP7_75t_L g13094 ( 
.A(n_11868),
.B(n_10923),
.Y(n_13094)
);

NAND2xp5_ASAP7_75t_L g13095 ( 
.A(n_11590),
.B(n_10928),
.Y(n_13095)
);

INVx5_ASAP7_75t_L g13096 ( 
.A(n_11890),
.Y(n_13096)
);

AND2x2_ASAP7_75t_L g13097 ( 
.A(n_11940),
.B(n_8715),
.Y(n_13097)
);

NAND2xp5_ASAP7_75t_L g13098 ( 
.A(n_11589),
.B(n_10929),
.Y(n_13098)
);

INVx2_ASAP7_75t_L g13099 ( 
.A(n_11890),
.Y(n_13099)
);

INVx2_ASAP7_75t_SL g13100 ( 
.A(n_11722),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_12264),
.Y(n_13101)
);

OR2x2_ASAP7_75t_L g13102 ( 
.A(n_11908),
.B(n_10933),
.Y(n_13102)
);

INVxp67_ASAP7_75t_SL g13103 ( 
.A(n_11612),
.Y(n_13103)
);

INVx1_ASAP7_75t_L g13104 ( 
.A(n_12092),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12092),
.Y(n_13105)
);

INVx1_ASAP7_75t_L g13106 ( 
.A(n_12246),
.Y(n_13106)
);

NAND2xp5_ASAP7_75t_L g13107 ( 
.A(n_11883),
.B(n_10936),
.Y(n_13107)
);

INVx2_ASAP7_75t_L g13108 ( 
.A(n_11722),
.Y(n_13108)
);

INVx1_ASAP7_75t_L g13109 ( 
.A(n_12246),
.Y(n_13109)
);

NAND2x1p5_ASAP7_75t_L g13110 ( 
.A(n_11685),
.B(n_8953),
.Y(n_13110)
);

AND2x2_ASAP7_75t_L g13111 ( 
.A(n_11942),
.B(n_8720),
.Y(n_13111)
);

AND2x4_ASAP7_75t_L g13112 ( 
.A(n_11962),
.B(n_10937),
.Y(n_13112)
);

AND2x2_ASAP7_75t_L g13113 ( 
.A(n_11953),
.B(n_8720),
.Y(n_13113)
);

INVx1_ASAP7_75t_L g13114 ( 
.A(n_12266),
.Y(n_13114)
);

INVx2_ASAP7_75t_L g13115 ( 
.A(n_11822),
.Y(n_13115)
);

BUFx3_ASAP7_75t_L g13116 ( 
.A(n_11956),
.Y(n_13116)
);

INVx2_ASAP7_75t_L g13117 ( 
.A(n_11822),
.Y(n_13117)
);

INVx1_ASAP7_75t_L g13118 ( 
.A(n_12266),
.Y(n_13118)
);

AND2x2_ASAP7_75t_L g13119 ( 
.A(n_11985),
.B(n_8720),
.Y(n_13119)
);

AND2x2_ASAP7_75t_L g13120 ( 
.A(n_11986),
.B(n_8725),
.Y(n_13120)
);

INVx1_ASAP7_75t_L g13121 ( 
.A(n_12267),
.Y(n_13121)
);

INVx2_ASAP7_75t_L g13122 ( 
.A(n_12239),
.Y(n_13122)
);

AND2x2_ASAP7_75t_L g13123 ( 
.A(n_11987),
.B(n_8725),
.Y(n_13123)
);

INVx2_ASAP7_75t_L g13124 ( 
.A(n_12281),
.Y(n_13124)
);

NAND2xp5_ASAP7_75t_L g13125 ( 
.A(n_11835),
.B(n_11639),
.Y(n_13125)
);

AND2x2_ASAP7_75t_L g13126 ( 
.A(n_11989),
.B(n_8725),
.Y(n_13126)
);

OR2x2_ASAP7_75t_L g13127 ( 
.A(n_12005),
.B(n_10949),
.Y(n_13127)
);

NAND2xp5_ASAP7_75t_L g13128 ( 
.A(n_11566),
.B(n_10957),
.Y(n_13128)
);

AND2x2_ASAP7_75t_L g13129 ( 
.A(n_12282),
.B(n_8748),
.Y(n_13129)
);

INVx2_ASAP7_75t_L g13130 ( 
.A(n_11915),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_12267),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12411),
.Y(n_13132)
);

HB1xp67_ASAP7_75t_L g13133 ( 
.A(n_11750),
.Y(n_13133)
);

INVx2_ASAP7_75t_L g13134 ( 
.A(n_11724),
.Y(n_13134)
);

AND2x4_ASAP7_75t_L g13135 ( 
.A(n_11916),
.B(n_10959),
.Y(n_13135)
);

INVx2_ASAP7_75t_L g13136 ( 
.A(n_11756),
.Y(n_13136)
);

INVx2_ASAP7_75t_L g13137 ( 
.A(n_11828),
.Y(n_13137)
);

AOI22xp33_ASAP7_75t_L g13138 ( 
.A1(n_11561),
.A2(n_9754),
.B1(n_9768),
.B2(n_9752),
.Y(n_13138)
);

OR2x2_ASAP7_75t_L g13139 ( 
.A(n_12007),
.B(n_10962),
.Y(n_13139)
);

INVx1_ASAP7_75t_L g13140 ( 
.A(n_12411),
.Y(n_13140)
);

OR2x2_ASAP7_75t_L g13141 ( 
.A(n_12015),
.B(n_10967),
.Y(n_13141)
);

NAND2x1_ASAP7_75t_L g13142 ( 
.A(n_11897),
.B(n_10589),
.Y(n_13142)
);

AND2x2_ASAP7_75t_L g13143 ( 
.A(n_12297),
.B(n_8748),
.Y(n_13143)
);

INVx2_ASAP7_75t_L g13144 ( 
.A(n_11865),
.Y(n_13144)
);

NAND2x1_ASAP7_75t_L g13145 ( 
.A(n_12161),
.B(n_11039),
.Y(n_13145)
);

INVx1_ASAP7_75t_L g13146 ( 
.A(n_11798),
.Y(n_13146)
);

INVx2_ASAP7_75t_L g13147 ( 
.A(n_12273),
.Y(n_13147)
);

INVxp67_ASAP7_75t_L g13148 ( 
.A(n_11557),
.Y(n_13148)
);

BUFx6f_ASAP7_75t_L g13149 ( 
.A(n_12504),
.Y(n_13149)
);

OR2x2_ASAP7_75t_L g13150 ( 
.A(n_12471),
.B(n_10968),
.Y(n_13150)
);

HB1xp67_ASAP7_75t_L g13151 ( 
.A(n_11939),
.Y(n_13151)
);

CKINVDCx20_ASAP7_75t_R g13152 ( 
.A(n_11873),
.Y(n_13152)
);

AND2x2_ASAP7_75t_L g13153 ( 
.A(n_11838),
.B(n_8748),
.Y(n_13153)
);

HB1xp67_ASAP7_75t_L g13154 ( 
.A(n_11787),
.Y(n_13154)
);

AND2x2_ASAP7_75t_L g13155 ( 
.A(n_11919),
.B(n_8779),
.Y(n_13155)
);

AND2x2_ASAP7_75t_L g13156 ( 
.A(n_11701),
.B(n_8779),
.Y(n_13156)
);

OR2x2_ASAP7_75t_L g13157 ( 
.A(n_12410),
.B(n_10969),
.Y(n_13157)
);

INVx2_ASAP7_75t_L g13158 ( 
.A(n_12397),
.Y(n_13158)
);

HB1xp67_ASAP7_75t_L g13159 ( 
.A(n_11964),
.Y(n_13159)
);

AND2x2_ASAP7_75t_L g13160 ( 
.A(n_11714),
.B(n_8779),
.Y(n_13160)
);

INVx2_ASAP7_75t_L g13161 ( 
.A(n_12137),
.Y(n_13161)
);

OR2x2_ASAP7_75t_L g13162 ( 
.A(n_12459),
.B(n_10970),
.Y(n_13162)
);

INVx2_ASAP7_75t_L g13163 ( 
.A(n_12058),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_11719),
.B(n_8782),
.Y(n_13164)
);

INVxp67_ASAP7_75t_SL g13165 ( 
.A(n_12153),
.Y(n_13165)
);

INVx4_ASAP7_75t_L g13166 ( 
.A(n_11884),
.Y(n_13166)
);

HB1xp67_ASAP7_75t_L g13167 ( 
.A(n_11777),
.Y(n_13167)
);

INVxp67_ASAP7_75t_L g13168 ( 
.A(n_11710),
.Y(n_13168)
);

AO21x2_ASAP7_75t_L g13169 ( 
.A1(n_11593),
.A2(n_10976),
.B(n_10973),
.Y(n_13169)
);

NAND2xp5_ASAP7_75t_L g13170 ( 
.A(n_11604),
.B(n_10982),
.Y(n_13170)
);

INVx1_ASAP7_75t_L g13171 ( 
.A(n_11798),
.Y(n_13171)
);

NAND2xp5_ASAP7_75t_L g13172 ( 
.A(n_11582),
.B(n_10986),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_12058),
.Y(n_13173)
);

INVx1_ASAP7_75t_L g13174 ( 
.A(n_11857),
.Y(n_13174)
);

AND2x2_ASAP7_75t_L g13175 ( 
.A(n_12162),
.B(n_8782),
.Y(n_13175)
);

AND2x4_ASAP7_75t_SL g13176 ( 
.A(n_11885),
.B(n_11900),
.Y(n_13176)
);

INVx1_ASAP7_75t_L g13177 ( 
.A(n_11857),
.Y(n_13177)
);

AND2x2_ASAP7_75t_L g13178 ( 
.A(n_11836),
.B(n_8782),
.Y(n_13178)
);

OR2x2_ASAP7_75t_L g13179 ( 
.A(n_12486),
.B(n_10990),
.Y(n_13179)
);

INVxp67_ASAP7_75t_SL g13180 ( 
.A(n_12102),
.Y(n_13180)
);

INVx2_ASAP7_75t_L g13181 ( 
.A(n_12058),
.Y(n_13181)
);

OR2x2_ASAP7_75t_L g13182 ( 
.A(n_12490),
.B(n_10994),
.Y(n_13182)
);

AND2x2_ASAP7_75t_L g13183 ( 
.A(n_11912),
.B(n_8829),
.Y(n_13183)
);

AND2x2_ASAP7_75t_L g13184 ( 
.A(n_11913),
.B(n_8829),
.Y(n_13184)
);

INVx1_ASAP7_75t_L g13185 ( 
.A(n_12099),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_11654),
.B(n_8829),
.Y(n_13186)
);

INVx3_ASAP7_75t_SL g13187 ( 
.A(n_12317),
.Y(n_13187)
);

BUFx2_ASAP7_75t_L g13188 ( 
.A(n_11933),
.Y(n_13188)
);

INVx1_ASAP7_75t_L g13189 ( 
.A(n_12099),
.Y(n_13189)
);

HB1xp67_ASAP7_75t_L g13190 ( 
.A(n_11777),
.Y(n_13190)
);

HB1xp67_ASAP7_75t_L g13191 ( 
.A(n_11851),
.Y(n_13191)
);

INVx1_ASAP7_75t_L g13192 ( 
.A(n_12223),
.Y(n_13192)
);

NAND2xp5_ASAP7_75t_L g13193 ( 
.A(n_11816),
.B(n_10997),
.Y(n_13193)
);

AND2x2_ASAP7_75t_L g13194 ( 
.A(n_11666),
.B(n_8849),
.Y(n_13194)
);

INVx1_ASAP7_75t_L g13195 ( 
.A(n_12223),
.Y(n_13195)
);

AND2x2_ASAP7_75t_L g13196 ( 
.A(n_11680),
.B(n_11698),
.Y(n_13196)
);

AND2x2_ASAP7_75t_L g13197 ( 
.A(n_12039),
.B(n_12041),
.Y(n_13197)
);

INVx1_ASAP7_75t_L g13198 ( 
.A(n_12507),
.Y(n_13198)
);

INVxp67_ASAP7_75t_L g13199 ( 
.A(n_12292),
.Y(n_13199)
);

NOR2x1_ASAP7_75t_L g13200 ( 
.A(n_11982),
.B(n_10998),
.Y(n_13200)
);

NAND2xp5_ASAP7_75t_L g13201 ( 
.A(n_11613),
.B(n_11000),
.Y(n_13201)
);

AND2x2_ASAP7_75t_L g13202 ( 
.A(n_12059),
.B(n_8849),
.Y(n_13202)
);

AND2x2_ASAP7_75t_L g13203 ( 
.A(n_12063),
.B(n_8849),
.Y(n_13203)
);

HB1xp67_ASAP7_75t_L g13204 ( 
.A(n_12081),
.Y(n_13204)
);

AOI22xp33_ASAP7_75t_L g13205 ( 
.A1(n_11673),
.A2(n_9768),
.B1(n_9874),
.B2(n_9754),
.Y(n_13205)
);

INVx2_ASAP7_75t_L g13206 ( 
.A(n_12100),
.Y(n_13206)
);

OR2x2_ASAP7_75t_L g13207 ( 
.A(n_12520),
.B(n_11007),
.Y(n_13207)
);

AND2x2_ASAP7_75t_L g13208 ( 
.A(n_12110),
.B(n_12333),
.Y(n_13208)
);

AO21x2_ASAP7_75t_L g13209 ( 
.A1(n_12298),
.A2(n_11012),
.B(n_11009),
.Y(n_13209)
);

HB1xp67_ASAP7_75t_L g13210 ( 
.A(n_12038),
.Y(n_13210)
);

AND2x2_ASAP7_75t_L g13211 ( 
.A(n_11951),
.B(n_8850),
.Y(n_13211)
);

INVx1_ASAP7_75t_L g13212 ( 
.A(n_12507),
.Y(n_13212)
);

INVxp67_ASAP7_75t_L g13213 ( 
.A(n_11882),
.Y(n_13213)
);

INVx2_ASAP7_75t_L g13214 ( 
.A(n_11889),
.Y(n_13214)
);

BUFx3_ASAP7_75t_L g13215 ( 
.A(n_11924),
.Y(n_13215)
);

NAND2x1p5_ASAP7_75t_L g13216 ( 
.A(n_11813),
.B(n_8953),
.Y(n_13216)
);

INVx2_ASAP7_75t_L g13217 ( 
.A(n_11891),
.Y(n_13217)
);

AND2x2_ASAP7_75t_L g13218 ( 
.A(n_11644),
.B(n_8850),
.Y(n_13218)
);

INVx1_ASAP7_75t_L g13219 ( 
.A(n_12029),
.Y(n_13219)
);

INVx1_ASAP7_75t_L g13220 ( 
.A(n_11824),
.Y(n_13220)
);

NOR2xp33_ASAP7_75t_L g13221 ( 
.A(n_11886),
.B(n_7551),
.Y(n_13221)
);

AND2x2_ASAP7_75t_L g13222 ( 
.A(n_12070),
.B(n_8850),
.Y(n_13222)
);

AND2x2_ASAP7_75t_L g13223 ( 
.A(n_12190),
.B(n_8856),
.Y(n_13223)
);

HB1xp67_ASAP7_75t_L g13224 ( 
.A(n_12233),
.Y(n_13224)
);

AND2x2_ASAP7_75t_L g13225 ( 
.A(n_12196),
.B(n_8856),
.Y(n_13225)
);

INVx1_ASAP7_75t_L g13226 ( 
.A(n_12289),
.Y(n_13226)
);

AND2x2_ASAP7_75t_L g13227 ( 
.A(n_11640),
.B(n_8856),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_11648),
.B(n_8874),
.Y(n_13228)
);

INVx1_ASAP7_75t_L g13229 ( 
.A(n_12296),
.Y(n_13229)
);

INVx2_ASAP7_75t_L g13230 ( 
.A(n_11927),
.Y(n_13230)
);

OR2x2_ASAP7_75t_L g13231 ( 
.A(n_11949),
.B(n_11657),
.Y(n_13231)
);

AND2x2_ASAP7_75t_L g13232 ( 
.A(n_11965),
.B(n_8874),
.Y(n_13232)
);

OR2x2_ASAP7_75t_L g13233 ( 
.A(n_11691),
.B(n_11018),
.Y(n_13233)
);

AND2x2_ASAP7_75t_L g13234 ( 
.A(n_12008),
.B(n_8874),
.Y(n_13234)
);

INVx2_ASAP7_75t_L g13235 ( 
.A(n_12259),
.Y(n_13235)
);

OR2x2_ASAP7_75t_L g13236 ( 
.A(n_11869),
.B(n_11019),
.Y(n_13236)
);

HB1xp67_ASAP7_75t_L g13237 ( 
.A(n_12082),
.Y(n_13237)
);

INVxp67_ASAP7_75t_L g13238 ( 
.A(n_12002),
.Y(n_13238)
);

INVx1_ASAP7_75t_SL g13239 ( 
.A(n_11774),
.Y(n_13239)
);

BUFx4f_ASAP7_75t_SL g13240 ( 
.A(n_11976),
.Y(n_13240)
);

INVx2_ASAP7_75t_L g13241 ( 
.A(n_12224),
.Y(n_13241)
);

INVxp67_ASAP7_75t_L g13242 ( 
.A(n_11735),
.Y(n_13242)
);

OR2x2_ASAP7_75t_L g13243 ( 
.A(n_11653),
.B(n_11026),
.Y(n_13243)
);

INVx2_ASAP7_75t_L g13244 ( 
.A(n_12224),
.Y(n_13244)
);

OR2x2_ASAP7_75t_L g13245 ( 
.A(n_12077),
.B(n_11033),
.Y(n_13245)
);

INVx1_ASAP7_75t_L g13246 ( 
.A(n_12062),
.Y(n_13246)
);

INVx1_ASAP7_75t_L g13247 ( 
.A(n_12294),
.Y(n_13247)
);

AND2x2_ASAP7_75t_L g13248 ( 
.A(n_12017),
.B(n_8915),
.Y(n_13248)
);

NOR2x1_ASAP7_75t_L g13249 ( 
.A(n_11704),
.B(n_11048),
.Y(n_13249)
);

INVx2_ASAP7_75t_L g13250 ( 
.A(n_12293),
.Y(n_13250)
);

AND2x2_ASAP7_75t_L g13251 ( 
.A(n_11791),
.B(n_8915),
.Y(n_13251)
);

INVx2_ASAP7_75t_L g13252 ( 
.A(n_12305),
.Y(n_13252)
);

AND2x2_ASAP7_75t_L g13253 ( 
.A(n_11720),
.B(n_11721),
.Y(n_13253)
);

OR2x2_ASAP7_75t_L g13254 ( 
.A(n_11765),
.B(n_11051),
.Y(n_13254)
);

INVx1_ASAP7_75t_L g13255 ( 
.A(n_12215),
.Y(n_13255)
);

INVx1_ASAP7_75t_L g13256 ( 
.A(n_11628),
.Y(n_13256)
);

INVxp67_ASAP7_75t_L g13257 ( 
.A(n_11575),
.Y(n_13257)
);

INVx2_ASAP7_75t_L g13258 ( 
.A(n_12313),
.Y(n_13258)
);

INVx1_ASAP7_75t_L g13259 ( 
.A(n_11818),
.Y(n_13259)
);

BUFx3_ASAP7_75t_L g13260 ( 
.A(n_11983),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_12329),
.Y(n_13261)
);

INVx2_ASAP7_75t_L g13262 ( 
.A(n_12346),
.Y(n_13262)
);

INVx1_ASAP7_75t_L g13263 ( 
.A(n_12394),
.Y(n_13263)
);

HB1xp67_ASAP7_75t_L g13264 ( 
.A(n_11749),
.Y(n_13264)
);

INVx2_ASAP7_75t_L g13265 ( 
.A(n_11728),
.Y(n_13265)
);

INVx1_ASAP7_75t_L g13266 ( 
.A(n_11699),
.Y(n_13266)
);

OR2x2_ASAP7_75t_L g13267 ( 
.A(n_11703),
.B(n_11053),
.Y(n_13267)
);

INVx2_ASAP7_75t_L g13268 ( 
.A(n_11728),
.Y(n_13268)
);

NAND2xp5_ASAP7_75t_L g13269 ( 
.A(n_11634),
.B(n_11054),
.Y(n_13269)
);

AND2x2_ASAP7_75t_L g13270 ( 
.A(n_12361),
.B(n_8915),
.Y(n_13270)
);

HB1xp67_ASAP7_75t_L g13271 ( 
.A(n_11984),
.Y(n_13271)
);

AND2x4_ASAP7_75t_SL g13272 ( 
.A(n_12114),
.B(n_7732),
.Y(n_13272)
);

INVx1_ASAP7_75t_L g13273 ( 
.A(n_11699),
.Y(n_13273)
);

AND2x2_ASAP7_75t_L g13274 ( 
.A(n_12362),
.B(n_8916),
.Y(n_13274)
);

INVx1_ASAP7_75t_L g13275 ( 
.A(n_12229),
.Y(n_13275)
);

INVx2_ASAP7_75t_L g13276 ( 
.A(n_11972),
.Y(n_13276)
);

INVx1_ASAP7_75t_L g13277 ( 
.A(n_11967),
.Y(n_13277)
);

OA21x2_ASAP7_75t_L g13278 ( 
.A1(n_11646),
.A2(n_10453),
.B(n_10445),
.Y(n_13278)
);

HB1xp67_ASAP7_75t_L g13279 ( 
.A(n_12415),
.Y(n_13279)
);

INVx1_ASAP7_75t_L g13280 ( 
.A(n_12505),
.Y(n_13280)
);

INVx2_ASAP7_75t_L g13281 ( 
.A(n_12279),
.Y(n_13281)
);

AND2x2_ASAP7_75t_L g13282 ( 
.A(n_12364),
.B(n_8916),
.Y(n_13282)
);

AND2x2_ASAP7_75t_L g13283 ( 
.A(n_11767),
.B(n_8916),
.Y(n_13283)
);

AND2x2_ASAP7_75t_L g13284 ( 
.A(n_12067),
.B(n_12127),
.Y(n_13284)
);

INVx2_ASAP7_75t_L g13285 ( 
.A(n_12468),
.Y(n_13285)
);

NAND2xp5_ASAP7_75t_L g13286 ( 
.A(n_11797),
.B(n_11057),
.Y(n_13286)
);

INVx1_ASAP7_75t_L g13287 ( 
.A(n_12506),
.Y(n_13287)
);

INVx2_ASAP7_75t_L g13288 ( 
.A(n_12469),
.Y(n_13288)
);

AND2x2_ASAP7_75t_L g13289 ( 
.A(n_11632),
.B(n_8955),
.Y(n_13289)
);

OR2x2_ASAP7_75t_L g13290 ( 
.A(n_12014),
.B(n_11060),
.Y(n_13290)
);

INVx2_ASAP7_75t_L g13291 ( 
.A(n_12477),
.Y(n_13291)
);

AND2x4_ASAP7_75t_L g13292 ( 
.A(n_12344),
.B(n_11063),
.Y(n_13292)
);

AND2x2_ASAP7_75t_L g13293 ( 
.A(n_12202),
.B(n_8955),
.Y(n_13293)
);

INVx1_ASAP7_75t_L g13294 ( 
.A(n_12506),
.Y(n_13294)
);

HB1xp67_ASAP7_75t_L g13295 ( 
.A(n_11743),
.Y(n_13295)
);

OR2x2_ASAP7_75t_L g13296 ( 
.A(n_11627),
.B(n_11065),
.Y(n_13296)
);

AND2x2_ASAP7_75t_L g13297 ( 
.A(n_12204),
.B(n_8955),
.Y(n_13297)
);

AND2x2_ASAP7_75t_L g13298 ( 
.A(n_12205),
.B(n_8970),
.Y(n_13298)
);

NAND2xp5_ASAP7_75t_L g13299 ( 
.A(n_12011),
.B(n_11066),
.Y(n_13299)
);

INVx2_ASAP7_75t_L g13300 ( 
.A(n_12483),
.Y(n_13300)
);

INVx3_ASAP7_75t_L g13301 ( 
.A(n_12335),
.Y(n_13301)
);

NAND2xp5_ASAP7_75t_L g13302 ( 
.A(n_11978),
.B(n_11078),
.Y(n_13302)
);

AND2x2_ASAP7_75t_L g13303 ( 
.A(n_12209),
.B(n_8970),
.Y(n_13303)
);

INVx1_ASAP7_75t_L g13304 ( 
.A(n_11694),
.Y(n_13304)
);

HB1xp67_ASAP7_75t_L g13305 ( 
.A(n_11772),
.Y(n_13305)
);

BUFx3_ASAP7_75t_L g13306 ( 
.A(n_12241),
.Y(n_13306)
);

INVx2_ASAP7_75t_L g13307 ( 
.A(n_12509),
.Y(n_13307)
);

INVx1_ASAP7_75t_L g13308 ( 
.A(n_11715),
.Y(n_13308)
);

INVx2_ASAP7_75t_SL g13309 ( 
.A(n_12136),
.Y(n_13309)
);

INVx4_ASAP7_75t_SL g13310 ( 
.A(n_11727),
.Y(n_13310)
);

BUFx3_ASAP7_75t_L g13311 ( 
.A(n_12261),
.Y(n_13311)
);

INVx1_ASAP7_75t_SL g13312 ( 
.A(n_11689),
.Y(n_13312)
);

AND2x2_ASAP7_75t_L g13313 ( 
.A(n_12245),
.B(n_8970),
.Y(n_13313)
);

INVx2_ASAP7_75t_L g13314 ( 
.A(n_12521),
.Y(n_13314)
);

AND2x4_ASAP7_75t_L g13315 ( 
.A(n_12172),
.B(n_11975),
.Y(n_13315)
);

INVx1_ASAP7_75t_L g13316 ( 
.A(n_11630),
.Y(n_13316)
);

INVx1_ASAP7_75t_L g13317 ( 
.A(n_11829),
.Y(n_13317)
);

AND2x2_ASAP7_75t_L g13318 ( 
.A(n_12247),
.B(n_9007),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_12304),
.Y(n_13319)
);

INVx1_ASAP7_75t_L g13320 ( 
.A(n_12355),
.Y(n_13320)
);

AOI22xp33_ASAP7_75t_L g13321 ( 
.A1(n_11574),
.A2(n_9768),
.B1(n_9874),
.B2(n_9754),
.Y(n_13321)
);

NAND2xp5_ASAP7_75t_L g13322 ( 
.A(n_11969),
.B(n_11085),
.Y(n_13322)
);

AND2x4_ASAP7_75t_L g13323 ( 
.A(n_12031),
.B(n_11086),
.Y(n_13323)
);

OR2x2_ASAP7_75t_L g13324 ( 
.A(n_11609),
.B(n_11089),
.Y(n_13324)
);

AND2x2_ASAP7_75t_L g13325 ( 
.A(n_12253),
.B(n_9007),
.Y(n_13325)
);

OR2x2_ASAP7_75t_L g13326 ( 
.A(n_12022),
.B(n_11099),
.Y(n_13326)
);

INVx1_ASAP7_75t_L g13327 ( 
.A(n_12368),
.Y(n_13327)
);

INVxp67_ASAP7_75t_SL g13328 ( 
.A(n_11638),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_12227),
.Y(n_13329)
);

NAND2xp5_ASAP7_75t_L g13330 ( 
.A(n_11979),
.B(n_11102),
.Y(n_13330)
);

AND2x4_ASAP7_75t_L g13331 ( 
.A(n_12302),
.B(n_11105),
.Y(n_13331)
);

AND2x2_ASAP7_75t_L g13332 ( 
.A(n_12365),
.B(n_9007),
.Y(n_13332)
);

INVx1_ASAP7_75t_L g13333 ( 
.A(n_11732),
.Y(n_13333)
);

INVx2_ASAP7_75t_L g13334 ( 
.A(n_12270),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_11670),
.Y(n_13335)
);

INVx1_ASAP7_75t_L g13336 ( 
.A(n_12433),
.Y(n_13336)
);

AND2x2_ASAP7_75t_L g13337 ( 
.A(n_12310),
.B(n_9754),
.Y(n_13337)
);

AND2x2_ASAP7_75t_L g13338 ( 
.A(n_12312),
.B(n_9768),
.Y(n_13338)
);

OR2x2_ASAP7_75t_L g13339 ( 
.A(n_11682),
.B(n_11117),
.Y(n_13339)
);

NAND2xp5_ASAP7_75t_L g13340 ( 
.A(n_11784),
.B(n_11118),
.Y(n_13340)
);

INVx1_ASAP7_75t_L g13341 ( 
.A(n_12163),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_12314),
.B(n_9768),
.Y(n_13342)
);

AND2x2_ASAP7_75t_L g13343 ( 
.A(n_12319),
.B(n_9768),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_12322),
.B(n_9874),
.Y(n_13344)
);

INVx1_ASAP7_75t_L g13345 ( 
.A(n_12389),
.Y(n_13345)
);

HB1xp67_ASAP7_75t_L g13346 ( 
.A(n_11910),
.Y(n_13346)
);

AND2x2_ASAP7_75t_L g13347 ( 
.A(n_12079),
.B(n_9874),
.Y(n_13347)
);

INVx2_ASAP7_75t_L g13348 ( 
.A(n_12056),
.Y(n_13348)
);

INVx2_ASAP7_75t_L g13349 ( 
.A(n_12194),
.Y(n_13349)
);

AND2x2_ASAP7_75t_L g13350 ( 
.A(n_12086),
.B(n_9874),
.Y(n_13350)
);

NAND2xp5_ASAP7_75t_L g13351 ( 
.A(n_11655),
.B(n_11121),
.Y(n_13351)
);

INVx2_ASAP7_75t_L g13352 ( 
.A(n_12201),
.Y(n_13352)
);

INVx3_ASAP7_75t_L g13353 ( 
.A(n_12134),
.Y(n_13353)
);

INVx2_ASAP7_75t_L g13354 ( 
.A(n_12272),
.Y(n_13354)
);

AND2x2_ASAP7_75t_L g13355 ( 
.A(n_12087),
.B(n_9874),
.Y(n_13355)
);

INVx1_ASAP7_75t_L g13356 ( 
.A(n_11905),
.Y(n_13356)
);

INVxp67_ASAP7_75t_L g13357 ( 
.A(n_11745),
.Y(n_13357)
);

INVx3_ASAP7_75t_SL g13358 ( 
.A(n_11837),
.Y(n_13358)
);

OR2x2_ASAP7_75t_L g13359 ( 
.A(n_11611),
.B(n_11123),
.Y(n_13359)
);

BUFx3_ASAP7_75t_L g13360 ( 
.A(n_12090),
.Y(n_13360)
);

INVx1_ASAP7_75t_L g13361 ( 
.A(n_11935),
.Y(n_13361)
);

INVx2_ASAP7_75t_L g13362 ( 
.A(n_12232),
.Y(n_13362)
);

INVxp67_ASAP7_75t_L g13363 ( 
.A(n_11862),
.Y(n_13363)
);

INVx1_ASAP7_75t_L g13364 ( 
.A(n_12168),
.Y(n_13364)
);

CKINVDCx20_ASAP7_75t_R g13365 ( 
.A(n_11782),
.Y(n_13365)
);

HB1xp67_ASAP7_75t_L g13366 ( 
.A(n_12112),
.Y(n_13366)
);

INVx2_ASAP7_75t_L g13367 ( 
.A(n_12260),
.Y(n_13367)
);

INVx2_ASAP7_75t_L g13368 ( 
.A(n_12271),
.Y(n_13368)
);

INVx2_ASAP7_75t_L g13369 ( 
.A(n_12193),
.Y(n_13369)
);

AND2x2_ASAP7_75t_L g13370 ( 
.A(n_12088),
.B(n_9963),
.Y(n_13370)
);

AND2x2_ASAP7_75t_L g13371 ( 
.A(n_12091),
.B(n_9963),
.Y(n_13371)
);

INVx1_ASAP7_75t_L g13372 ( 
.A(n_12517),
.Y(n_13372)
);

INVxp67_ASAP7_75t_L g13373 ( 
.A(n_11587),
.Y(n_13373)
);

INVx2_ASAP7_75t_L g13374 ( 
.A(n_12393),
.Y(n_13374)
);

OR2x2_ASAP7_75t_L g13375 ( 
.A(n_11693),
.B(n_11125),
.Y(n_13375)
);

INVx2_ASAP7_75t_L g13376 ( 
.A(n_12403),
.Y(n_13376)
);

INVx2_ASAP7_75t_L g13377 ( 
.A(n_12466),
.Y(n_13377)
);

INVx1_ASAP7_75t_L g13378 ( 
.A(n_11614),
.Y(n_13378)
);

AND2x2_ASAP7_75t_L g13379 ( 
.A(n_12332),
.B(n_9963),
.Y(n_13379)
);

INVx1_ASAP7_75t_L g13380 ( 
.A(n_12519),
.Y(n_13380)
);

AND2x2_ASAP7_75t_L g13381 ( 
.A(n_12347),
.B(n_9963),
.Y(n_13381)
);

HB1xp67_ASAP7_75t_L g13382 ( 
.A(n_12131),
.Y(n_13382)
);

AND2x2_ASAP7_75t_L g13383 ( 
.A(n_12126),
.B(n_9963),
.Y(n_13383)
);

AND2x2_ASAP7_75t_L g13384 ( 
.A(n_12262),
.B(n_9963),
.Y(n_13384)
);

INVx1_ASAP7_75t_L g13385 ( 
.A(n_11845),
.Y(n_13385)
);

INVx1_ASAP7_75t_L g13386 ( 
.A(n_12398),
.Y(n_13386)
);

AND2x4_ASAP7_75t_L g13387 ( 
.A(n_12283),
.B(n_11126),
.Y(n_13387)
);

OR2x2_ASAP7_75t_L g13388 ( 
.A(n_11930),
.B(n_11129),
.Y(n_13388)
);

NAND2xp5_ASAP7_75t_L g13389 ( 
.A(n_11696),
.B(n_11134),
.Y(n_13389)
);

INVx2_ASAP7_75t_L g13390 ( 
.A(n_12489),
.Y(n_13390)
);

INVx2_ASAP7_75t_L g13391 ( 
.A(n_12498),
.Y(n_13391)
);

INVx2_ASAP7_75t_L g13392 ( 
.A(n_12513),
.Y(n_13392)
);

INVx1_ASAP7_75t_L g13393 ( 
.A(n_12409),
.Y(n_13393)
);

INVx2_ASAP7_75t_L g13394 ( 
.A(n_12009),
.Y(n_13394)
);

NAND2xp5_ASAP7_75t_L g13395 ( 
.A(n_11619),
.B(n_11139),
.Y(n_13395)
);

AND2x2_ASAP7_75t_L g13396 ( 
.A(n_12263),
.B(n_9983),
.Y(n_13396)
);

INVx2_ASAP7_75t_L g13397 ( 
.A(n_12417),
.Y(n_13397)
);

INVx1_ASAP7_75t_L g13398 ( 
.A(n_12427),
.Y(n_13398)
);

AND2x2_ASAP7_75t_L g13399 ( 
.A(n_12256),
.B(n_9983),
.Y(n_13399)
);

INVx1_ASAP7_75t_L g13400 ( 
.A(n_12494),
.Y(n_13400)
);

AND2x2_ASAP7_75t_L g13401 ( 
.A(n_12107),
.B(n_9983),
.Y(n_13401)
);

INVxp67_ASAP7_75t_L g13402 ( 
.A(n_11852),
.Y(n_13402)
);

INVx3_ASAP7_75t_L g13403 ( 
.A(n_12203),
.Y(n_13403)
);

AND2x2_ASAP7_75t_L g13404 ( 
.A(n_12444),
.B(n_9983),
.Y(n_13404)
);

HB1xp67_ASAP7_75t_L g13405 ( 
.A(n_11892),
.Y(n_13405)
);

BUFx6f_ASAP7_75t_L g13406 ( 
.A(n_12311),
.Y(n_13406)
);

INVx1_ASAP7_75t_L g13407 ( 
.A(n_12388),
.Y(n_13407)
);

INVx1_ASAP7_75t_L g13408 ( 
.A(n_12401),
.Y(n_13408)
);

AND2x2_ASAP7_75t_L g13409 ( 
.A(n_12111),
.B(n_9983),
.Y(n_13409)
);

BUFx3_ASAP7_75t_L g13410 ( 
.A(n_11789),
.Y(n_13410)
);

HB1xp67_ASAP7_75t_L g13411 ( 
.A(n_11904),
.Y(n_13411)
);

INVx4_ASAP7_75t_R g13412 ( 
.A(n_11636),
.Y(n_13412)
);

HB1xp67_ASAP7_75t_L g13413 ( 
.A(n_12060),
.Y(n_13413)
);

BUFx3_ASAP7_75t_L g13414 ( 
.A(n_11842),
.Y(n_13414)
);

BUFx3_ASAP7_75t_L g13415 ( 
.A(n_12212),
.Y(n_13415)
);

INVxp67_ASAP7_75t_SL g13416 ( 
.A(n_11877),
.Y(n_13416)
);

INVx2_ASAP7_75t_L g13417 ( 
.A(n_12219),
.Y(n_13417)
);

AND2x2_ASAP7_75t_L g13418 ( 
.A(n_12288),
.B(n_9983),
.Y(n_13418)
);

INVx2_ASAP7_75t_L g13419 ( 
.A(n_12225),
.Y(n_13419)
);

OR2x2_ASAP7_75t_L g13420 ( 
.A(n_11793),
.B(n_11141),
.Y(n_13420)
);

BUFx2_ASAP7_75t_L g13421 ( 
.A(n_12010),
.Y(n_13421)
);

OR2x6_ASAP7_75t_L g13422 ( 
.A(n_11895),
.B(n_9990),
.Y(n_13422)
);

HB1xp67_ASAP7_75t_L g13423 ( 
.A(n_12336),
.Y(n_13423)
);

INVx2_ASAP7_75t_L g13424 ( 
.A(n_12230),
.Y(n_13424)
);

INVx1_ASAP7_75t_L g13425 ( 
.A(n_12405),
.Y(n_13425)
);

INVx1_ASAP7_75t_L g13426 ( 
.A(n_12447),
.Y(n_13426)
);

INVx4_ASAP7_75t_R g13427 ( 
.A(n_11843),
.Y(n_13427)
);

HB1xp67_ASAP7_75t_L g13428 ( 
.A(n_12343),
.Y(n_13428)
);

AND2x2_ASAP7_75t_L g13429 ( 
.A(n_12295),
.B(n_9990),
.Y(n_13429)
);

INVx2_ASAP7_75t_L g13430 ( 
.A(n_12023),
.Y(n_13430)
);

INVx2_ASAP7_75t_L g13431 ( 
.A(n_12307),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_12306),
.B(n_9990),
.Y(n_13432)
);

INVx2_ASAP7_75t_SL g13433 ( 
.A(n_12340),
.Y(n_13433)
);

INVx2_ASAP7_75t_L g13434 ( 
.A(n_12049),
.Y(n_13434)
);

INVx1_ASAP7_75t_L g13435 ( 
.A(n_12457),
.Y(n_13435)
);

NAND2xp5_ASAP7_75t_L g13436 ( 
.A(n_12123),
.B(n_11142),
.Y(n_13436)
);

INVx2_ASAP7_75t_L g13437 ( 
.A(n_12043),
.Y(n_13437)
);

BUFx12f_ASAP7_75t_L g13438 ( 
.A(n_11790),
.Y(n_13438)
);

INVx1_ASAP7_75t_L g13439 ( 
.A(n_12069),
.Y(n_13439)
);

INVx1_ASAP7_75t_L g13440 ( 
.A(n_12467),
.Y(n_13440)
);

NAND2xp5_ASAP7_75t_L g13441 ( 
.A(n_11855),
.B(n_11155),
.Y(n_13441)
);

AND2x2_ASAP7_75t_L g13442 ( 
.A(n_12525),
.B(n_11833),
.Y(n_13442)
);

INVx1_ASAP7_75t_L g13443 ( 
.A(n_12542),
.Y(n_13443)
);

INVx1_ASAP7_75t_L g13444 ( 
.A(n_12546),
.Y(n_13444)
);

INVxp67_ASAP7_75t_SL g13445 ( 
.A(n_12607),
.Y(n_13445)
);

AND2x2_ASAP7_75t_L g13446 ( 
.A(n_12573),
.B(n_11995),
.Y(n_13446)
);

INVx1_ASAP7_75t_L g13447 ( 
.A(n_12567),
.Y(n_13447)
);

NAND2xp5_ASAP7_75t_L g13448 ( 
.A(n_12663),
.B(n_12527),
.Y(n_13448)
);

AND2x2_ASAP7_75t_L g13449 ( 
.A(n_12626),
.B(n_11731),
.Y(n_13449)
);

OR2x2_ASAP7_75t_L g13450 ( 
.A(n_12568),
.B(n_11717),
.Y(n_13450)
);

AND2x4_ASAP7_75t_L g13451 ( 
.A(n_12700),
.B(n_9990),
.Y(n_13451)
);

OR2x2_ASAP7_75t_L g13452 ( 
.A(n_13170),
.B(n_11808),
.Y(n_13452)
);

AOI22xp5_ASAP7_75t_L g13453 ( 
.A1(n_13328),
.A2(n_11667),
.B1(n_12119),
.B2(n_12257),
.Y(n_13453)
);

INVx2_ASAP7_75t_SL g13454 ( 
.A(n_12607),
.Y(n_13454)
);

NOR2x1p5_ASAP7_75t_L g13455 ( 
.A(n_13049),
.B(n_7555),
.Y(n_13455)
);

HB1xp67_ASAP7_75t_L g13456 ( 
.A(n_12583),
.Y(n_13456)
);

INVx1_ASAP7_75t_L g13457 ( 
.A(n_12531),
.Y(n_13457)
);

OR2x2_ASAP7_75t_L g13458 ( 
.A(n_12537),
.B(n_12185),
.Y(n_13458)
);

AND2x2_ASAP7_75t_L g13459 ( 
.A(n_12524),
.B(n_11738),
.Y(n_13459)
);

AND2x4_ASAP7_75t_L g13460 ( 
.A(n_12700),
.B(n_9990),
.Y(n_13460)
);

NOR2x1_ASAP7_75t_L g13461 ( 
.A(n_13074),
.B(n_12016),
.Y(n_13461)
);

INVx1_ASAP7_75t_SL g13462 ( 
.A(n_12596),
.Y(n_13462)
);

INVx2_ASAP7_75t_L g13463 ( 
.A(n_12602),
.Y(n_13463)
);

INVx1_ASAP7_75t_L g13464 ( 
.A(n_12561),
.Y(n_13464)
);

NAND2xp5_ASAP7_75t_L g13465 ( 
.A(n_13239),
.B(n_12030),
.Y(n_13465)
);

INVx1_ASAP7_75t_L g13466 ( 
.A(n_12561),
.Y(n_13466)
);

AND2x2_ASAP7_75t_L g13467 ( 
.A(n_12655),
.B(n_12455),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_12785),
.Y(n_13468)
);

OR2x2_ASAP7_75t_L g13469 ( 
.A(n_13002),
.B(n_11820),
.Y(n_13469)
);

INVxp67_ASAP7_75t_L g13470 ( 
.A(n_12607),
.Y(n_13470)
);

AND2x2_ASAP7_75t_L g13471 ( 
.A(n_12868),
.B(n_13066),
.Y(n_13471)
);

INVx1_ASAP7_75t_SL g13472 ( 
.A(n_12648),
.Y(n_13472)
);

INVx1_ASAP7_75t_L g13473 ( 
.A(n_12788),
.Y(n_13473)
);

AND2x2_ASAP7_75t_L g13474 ( 
.A(n_13066),
.B(n_12286),
.Y(n_13474)
);

INVxp33_ASAP7_75t_SL g13475 ( 
.A(n_12733),
.Y(n_13475)
);

INVx1_ASAP7_75t_L g13476 ( 
.A(n_12523),
.Y(n_13476)
);

INVx1_ASAP7_75t_L g13477 ( 
.A(n_12523),
.Y(n_13477)
);

BUFx2_ASAP7_75t_L g13478 ( 
.A(n_13066),
.Y(n_13478)
);

AND2x2_ASAP7_75t_L g13479 ( 
.A(n_12747),
.B(n_12536),
.Y(n_13479)
);

INVx1_ASAP7_75t_L g13480 ( 
.A(n_12535),
.Y(n_13480)
);

INVx1_ASAP7_75t_L g13481 ( 
.A(n_12535),
.Y(n_13481)
);

INVx1_ASAP7_75t_L g13482 ( 
.A(n_12543),
.Y(n_13482)
);

INVx3_ASAP7_75t_L g13483 ( 
.A(n_12585),
.Y(n_13483)
);

NAND2xp5_ASAP7_75t_L g13484 ( 
.A(n_13246),
.B(n_11859),
.Y(n_13484)
);

INVx1_ASAP7_75t_L g13485 ( 
.A(n_12543),
.Y(n_13485)
);

INVx1_ASAP7_75t_L g13486 ( 
.A(n_12549),
.Y(n_13486)
);

OA21x2_ASAP7_75t_L g13487 ( 
.A1(n_13266),
.A2(n_12479),
.B(n_11957),
.Y(n_13487)
);

NAND2xp5_ASAP7_75t_L g13488 ( 
.A(n_13246),
.B(n_11812),
.Y(n_13488)
);

BUFx2_ASAP7_75t_L g13489 ( 
.A(n_13085),
.Y(n_13489)
);

INVx1_ASAP7_75t_L g13490 ( 
.A(n_12549),
.Y(n_13490)
);

INVx2_ASAP7_75t_L g13491 ( 
.A(n_12589),
.Y(n_13491)
);

INVx1_ASAP7_75t_L g13492 ( 
.A(n_12550),
.Y(n_13492)
);

NAND2xp5_ASAP7_75t_L g13493 ( 
.A(n_13255),
.B(n_11814),
.Y(n_13493)
);

NAND2xp5_ASAP7_75t_L g13494 ( 
.A(n_13255),
.B(n_11847),
.Y(n_13494)
);

AOI22xp33_ASAP7_75t_L g13495 ( 
.A1(n_13295),
.A2(n_11697),
.B1(n_12145),
.B2(n_12044),
.Y(n_13495)
);

CKINVDCx5p33_ASAP7_75t_R g13496 ( 
.A(n_12544),
.Y(n_13496)
);

INVx2_ASAP7_75t_SL g13497 ( 
.A(n_12827),
.Y(n_13497)
);

AND2x2_ASAP7_75t_L g13498 ( 
.A(n_12538),
.B(n_12440),
.Y(n_13498)
);

AND2x2_ASAP7_75t_L g13499 ( 
.A(n_12562),
.B(n_12073),
.Y(n_13499)
);

INVx1_ASAP7_75t_L g13500 ( 
.A(n_12550),
.Y(n_13500)
);

INVx2_ASAP7_75t_L g13501 ( 
.A(n_12589),
.Y(n_13501)
);

INVx3_ASAP7_75t_L g13502 ( 
.A(n_12585),
.Y(n_13502)
);

NOR2xp33_ASAP7_75t_L g13503 ( 
.A(n_12613),
.B(n_7557),
.Y(n_13503)
);

AND2x2_ASAP7_75t_L g13504 ( 
.A(n_12591),
.B(n_12104),
.Y(n_13504)
);

AND2x2_ASAP7_75t_L g13505 ( 
.A(n_12853),
.B(n_12238),
.Y(n_13505)
);

NAND2xp5_ASAP7_75t_L g13506 ( 
.A(n_13416),
.B(n_12473),
.Y(n_13506)
);

AOI22xp33_ASAP7_75t_L g13507 ( 
.A1(n_13305),
.A2(n_11794),
.B1(n_12033),
.B2(n_12158),
.Y(n_13507)
);

AND2x2_ASAP7_75t_L g13508 ( 
.A(n_12565),
.B(n_12445),
.Y(n_13508)
);

INVx1_ASAP7_75t_L g13509 ( 
.A(n_12552),
.Y(n_13509)
);

NAND2xp5_ASAP7_75t_L g13510 ( 
.A(n_13242),
.B(n_12502),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_12552),
.Y(n_13511)
);

HB1xp67_ASAP7_75t_L g13512 ( 
.A(n_13100),
.Y(n_13512)
);

BUFx2_ASAP7_75t_L g13513 ( 
.A(n_12630),
.Y(n_13513)
);

INVx2_ASAP7_75t_L g13514 ( 
.A(n_12761),
.Y(n_13514)
);

INVx1_ASAP7_75t_L g13515 ( 
.A(n_12553),
.Y(n_13515)
);

AOI22xp33_ASAP7_75t_L g13516 ( 
.A1(n_13438),
.A2(n_12249),
.B1(n_12250),
.B2(n_11832),
.Y(n_13516)
);

AND2x2_ASAP7_75t_L g13517 ( 
.A(n_12724),
.B(n_12448),
.Y(n_13517)
);

AND2x4_ASAP7_75t_L g13518 ( 
.A(n_12630),
.B(n_9990),
.Y(n_13518)
);

INVx1_ASAP7_75t_L g13519 ( 
.A(n_12553),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_12556),
.Y(n_13520)
);

NAND2xp5_ASAP7_75t_L g13521 ( 
.A(n_13151),
.B(n_12235),
.Y(n_13521)
);

INVx1_ASAP7_75t_L g13522 ( 
.A(n_12556),
.Y(n_13522)
);

OAI22xp5_ASAP7_75t_L g13523 ( 
.A1(n_12931),
.A2(n_12478),
.B1(n_12465),
.B2(n_12441),
.Y(n_13523)
);

INVx1_ASAP7_75t_L g13524 ( 
.A(n_12812),
.Y(n_13524)
);

OR2x2_ASAP7_75t_L g13525 ( 
.A(n_13095),
.B(n_11971),
.Y(n_13525)
);

INVx2_ASAP7_75t_L g13526 ( 
.A(n_12590),
.Y(n_13526)
);

HB1xp67_ASAP7_75t_L g13527 ( 
.A(n_13154),
.Y(n_13527)
);

INVx1_ASAP7_75t_L g13528 ( 
.A(n_12814),
.Y(n_13528)
);

INVx1_ASAP7_75t_L g13529 ( 
.A(n_12574),
.Y(n_13529)
);

OAI22xp33_ASAP7_75t_L g13530 ( 
.A1(n_12547),
.A2(n_12118),
.B1(n_12395),
.B2(n_12345),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_12574),
.Y(n_13531)
);

INVxp67_ASAP7_75t_L g13532 ( 
.A(n_12989),
.Y(n_13532)
);

INVx2_ASAP7_75t_L g13533 ( 
.A(n_12590),
.Y(n_13533)
);

NAND2xp5_ASAP7_75t_L g13534 ( 
.A(n_12836),
.B(n_12321),
.Y(n_13534)
);

INVx2_ASAP7_75t_L g13535 ( 
.A(n_12669),
.Y(n_13535)
);

NAND2xp5_ASAP7_75t_SL g13536 ( 
.A(n_12541),
.B(n_11853),
.Y(n_13536)
);

AND2x2_ASAP7_75t_L g13537 ( 
.A(n_12647),
.B(n_12554),
.Y(n_13537)
);

INVx2_ASAP7_75t_SL g13538 ( 
.A(n_12827),
.Y(n_13538)
);

INVx2_ASAP7_75t_L g13539 ( 
.A(n_12554),
.Y(n_13539)
);

INVx1_ASAP7_75t_L g13540 ( 
.A(n_12577),
.Y(n_13540)
);

INVx1_ASAP7_75t_L g13541 ( 
.A(n_12577),
.Y(n_13541)
);

HB1xp67_ASAP7_75t_L g13542 ( 
.A(n_13159),
.Y(n_13542)
);

INVx2_ASAP7_75t_L g13543 ( 
.A(n_12534),
.Y(n_13543)
);

AND2x4_ASAP7_75t_L g13544 ( 
.A(n_12827),
.B(n_10011),
.Y(n_13544)
);

INVx2_ASAP7_75t_SL g13545 ( 
.A(n_13096),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_12578),
.Y(n_13546)
);

OAI222xp33_ASAP7_75t_L g13547 ( 
.A1(n_12823),
.A2(n_11864),
.B1(n_12299),
.B2(n_12328),
.C1(n_12354),
.C2(n_12352),
.Y(n_13547)
);

AND2x2_ASAP7_75t_L g13548 ( 
.A(n_12540),
.B(n_12487),
.Y(n_13548)
);

AND2x2_ASAP7_75t_L g13549 ( 
.A(n_12545),
.B(n_12508),
.Y(n_13549)
);

INVx1_ASAP7_75t_SL g13550 ( 
.A(n_12576),
.Y(n_13550)
);

AOI22xp33_ASAP7_75t_L g13551 ( 
.A1(n_13403),
.A2(n_11839),
.B1(n_11876),
.B2(n_11903),
.Y(n_13551)
);

INVx1_ASAP7_75t_L g13552 ( 
.A(n_12578),
.Y(n_13552)
);

BUFx2_ASAP7_75t_SL g13553 ( 
.A(n_12705),
.Y(n_13553)
);

HB1xp67_ASAP7_75t_L g13554 ( 
.A(n_12915),
.Y(n_13554)
);

AND2x2_ASAP7_75t_L g13555 ( 
.A(n_12806),
.B(n_12510),
.Y(n_13555)
);

NAND2xp5_ASAP7_75t_L g13556 ( 
.A(n_12839),
.B(n_12280),
.Y(n_13556)
);

AOI22xp33_ASAP7_75t_L g13557 ( 
.A1(n_13403),
.A2(n_11925),
.B1(n_12177),
.B2(n_12046),
.Y(n_13557)
);

HB1xp67_ASAP7_75t_L g13558 ( 
.A(n_13108),
.Y(n_13558)
);

NAND2xp5_ASAP7_75t_L g13559 ( 
.A(n_13210),
.B(n_12287),
.Y(n_13559)
);

INVx2_ASAP7_75t_L g13560 ( 
.A(n_12534),
.Y(n_13560)
);

INVx2_ASAP7_75t_L g13561 ( 
.A(n_12673),
.Y(n_13561)
);

BUFx2_ASAP7_75t_L g13562 ( 
.A(n_13169),
.Y(n_13562)
);

NOR2xp33_ASAP7_75t_L g13563 ( 
.A(n_12705),
.B(n_7557),
.Y(n_13563)
);

NAND2xp5_ASAP7_75t_L g13564 ( 
.A(n_13220),
.B(n_13237),
.Y(n_13564)
);

INVx1_ASAP7_75t_L g13565 ( 
.A(n_12586),
.Y(n_13565)
);

NAND2xp5_ASAP7_75t_L g13566 ( 
.A(n_13220),
.B(n_12303),
.Y(n_13566)
);

INVx1_ASAP7_75t_SL g13567 ( 
.A(n_12617),
.Y(n_13567)
);

AND2x2_ASAP7_75t_L g13568 ( 
.A(n_12559),
.B(n_12560),
.Y(n_13568)
);

INVx2_ASAP7_75t_L g13569 ( 
.A(n_12623),
.Y(n_13569)
);

AND2x2_ASAP7_75t_L g13570 ( 
.A(n_12564),
.B(n_12514),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_12586),
.Y(n_13571)
);

INVx1_ASAP7_75t_L g13572 ( 
.A(n_12592),
.Y(n_13572)
);

INVx1_ASAP7_75t_L g13573 ( 
.A(n_12592),
.Y(n_13573)
);

OAI221xp5_ASAP7_75t_L g13574 ( 
.A1(n_12533),
.A2(n_12035),
.B1(n_12037),
.B2(n_12027),
.C(n_12370),
.Y(n_13574)
);

OR2x2_ASAP7_75t_L g13575 ( 
.A(n_12526),
.B(n_11159),
.Y(n_13575)
);

HB1xp67_ASAP7_75t_L g13576 ( 
.A(n_12679),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_12594),
.Y(n_13577)
);

AND2x2_ASAP7_75t_L g13578 ( 
.A(n_12682),
.B(n_12522),
.Y(n_13578)
);

AND2x2_ASAP7_75t_L g13579 ( 
.A(n_12813),
.B(n_12849),
.Y(n_13579)
);

NAND2xp5_ASAP7_75t_L g13580 ( 
.A(n_13213),
.B(n_12275),
.Y(n_13580)
);

INVx2_ASAP7_75t_L g13581 ( 
.A(n_12623),
.Y(n_13581)
);

INVx2_ASAP7_75t_SL g13582 ( 
.A(n_13096),
.Y(n_13582)
);

AND2x2_ASAP7_75t_L g13583 ( 
.A(n_12638),
.B(n_12481),
.Y(n_13583)
);

AND2x4_ASAP7_75t_L g13584 ( 
.A(n_12653),
.B(n_10011),
.Y(n_13584)
);

INVx1_ASAP7_75t_L g13585 ( 
.A(n_12594),
.Y(n_13585)
);

AOI22xp33_ASAP7_75t_L g13586 ( 
.A1(n_13021),
.A2(n_12277),
.B1(n_12220),
.B2(n_12026),
.Y(n_13586)
);

INVx2_ASAP7_75t_L g13587 ( 
.A(n_12653),
.Y(n_13587)
);

INVx2_ASAP7_75t_L g13588 ( 
.A(n_12658),
.Y(n_13588)
);

INVx1_ASAP7_75t_L g13589 ( 
.A(n_12599),
.Y(n_13589)
);

HB1xp67_ASAP7_75t_L g13590 ( 
.A(n_12820),
.Y(n_13590)
);

INVx1_ASAP7_75t_L g13591 ( 
.A(n_12599),
.Y(n_13591)
);

NAND2xp5_ASAP7_75t_L g13592 ( 
.A(n_12838),
.B(n_12385),
.Y(n_13592)
);

NAND2xp5_ASAP7_75t_L g13593 ( 
.A(n_12855),
.B(n_12378),
.Y(n_13593)
);

INVx1_ASAP7_75t_L g13594 ( 
.A(n_12601),
.Y(n_13594)
);

INVx1_ASAP7_75t_L g13595 ( 
.A(n_12601),
.Y(n_13595)
);

INVx2_ASAP7_75t_L g13596 ( 
.A(n_12658),
.Y(n_13596)
);

AND2x2_ASAP7_75t_L g13597 ( 
.A(n_12794),
.B(n_12456),
.Y(n_13597)
);

INVx1_ASAP7_75t_L g13598 ( 
.A(n_12603),
.Y(n_13598)
);

INVx2_ASAP7_75t_L g13599 ( 
.A(n_12932),
.Y(n_13599)
);

AND2x2_ASAP7_75t_L g13600 ( 
.A(n_12645),
.B(n_12685),
.Y(n_13600)
);

INVx2_ASAP7_75t_L g13601 ( 
.A(n_12932),
.Y(n_13601)
);

INVx3_ASAP7_75t_L g13602 ( 
.A(n_12743),
.Y(n_13602)
);

AND2x2_ASAP7_75t_L g13603 ( 
.A(n_12615),
.B(n_12367),
.Y(n_13603)
);

INVx3_ASAP7_75t_L g13604 ( 
.A(n_12743),
.Y(n_13604)
);

NAND2xp5_ASAP7_75t_L g13605 ( 
.A(n_12913),
.B(n_12372),
.Y(n_13605)
);

INVx1_ASAP7_75t_L g13606 ( 
.A(n_12603),
.Y(n_13606)
);

AND2x2_ASAP7_75t_L g13607 ( 
.A(n_12622),
.B(n_12463),
.Y(n_13607)
);

INVx2_ASAP7_75t_L g13608 ( 
.A(n_12932),
.Y(n_13608)
);

INVx3_ASAP7_75t_L g13609 ( 
.A(n_12632),
.Y(n_13609)
);

OAI22xp5_ASAP7_75t_SL g13610 ( 
.A1(n_13031),
.A2(n_7560),
.B1(n_7593),
.B2(n_7563),
.Y(n_13610)
);

AOI22xp33_ASAP7_75t_L g13611 ( 
.A1(n_13414),
.A2(n_13256),
.B1(n_13378),
.B2(n_13410),
.Y(n_13611)
);

INVx1_ASAP7_75t_L g13612 ( 
.A(n_12604),
.Y(n_13612)
);

AND2x2_ASAP7_75t_L g13613 ( 
.A(n_12941),
.B(n_12475),
.Y(n_13613)
);

AND2x2_ASAP7_75t_L g13614 ( 
.A(n_12624),
.B(n_12413),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_12604),
.Y(n_13615)
);

INVx1_ASAP7_75t_L g13616 ( 
.A(n_12606),
.Y(n_13616)
);

INVx2_ASAP7_75t_L g13617 ( 
.A(n_12639),
.Y(n_13617)
);

INVx1_ASAP7_75t_L g13618 ( 
.A(n_12606),
.Y(n_13618)
);

INVx1_ASAP7_75t_L g13619 ( 
.A(n_12611),
.Y(n_13619)
);

INVx1_ASAP7_75t_L g13620 ( 
.A(n_12611),
.Y(n_13620)
);

INVx1_ASAP7_75t_L g13621 ( 
.A(n_12616),
.Y(n_13621)
);

INVxp67_ASAP7_75t_L g13622 ( 
.A(n_12532),
.Y(n_13622)
);

AND2x4_ASAP7_75t_L g13623 ( 
.A(n_12551),
.B(n_10011),
.Y(n_13623)
);

HB1xp67_ASAP7_75t_L g13624 ( 
.A(n_12920),
.Y(n_13624)
);

NAND2xp5_ASAP7_75t_L g13625 ( 
.A(n_13148),
.B(n_12374),
.Y(n_13625)
);

INVx1_ASAP7_75t_L g13626 ( 
.A(n_12616),
.Y(n_13626)
);

OR2x2_ASAP7_75t_L g13627 ( 
.A(n_12977),
.B(n_11170),
.Y(n_13627)
);

OAI21xp33_ASAP7_75t_L g13628 ( 
.A1(n_13316),
.A2(n_12383),
.B(n_12379),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_12949),
.Y(n_13629)
);

INVxp67_ASAP7_75t_SL g13630 ( 
.A(n_12976),
.Y(n_13630)
);

NAND2xp5_ASAP7_75t_L g13631 ( 
.A(n_12712),
.B(n_11172),
.Y(n_13631)
);

AND2x2_ASAP7_75t_L g13632 ( 
.A(n_12631),
.B(n_12416),
.Y(n_13632)
);

OR2x2_ASAP7_75t_L g13633 ( 
.A(n_13326),
.B(n_11173),
.Y(n_13633)
);

AND2x2_ASAP7_75t_L g13634 ( 
.A(n_12633),
.B(n_12637),
.Y(n_13634)
);

INVx1_ASAP7_75t_L g13635 ( 
.A(n_12621),
.Y(n_13635)
);

BUFx2_ASAP7_75t_L g13636 ( 
.A(n_13310),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_12621),
.Y(n_13637)
);

AND2x2_ASAP7_75t_L g13638 ( 
.A(n_13166),
.B(n_12323),
.Y(n_13638)
);

OR2x2_ASAP7_75t_L g13639 ( 
.A(n_12539),
.B(n_11177),
.Y(n_13639)
);

BUFx2_ASAP7_75t_L g13640 ( 
.A(n_13310),
.Y(n_13640)
);

AOI22xp33_ASAP7_75t_SL g13641 ( 
.A1(n_13165),
.A2(n_12021),
.B1(n_11815),
.B2(n_11810),
.Y(n_13641)
);

INVx1_ASAP7_75t_L g13642 ( 
.A(n_12723),
.Y(n_13642)
);

AND2x2_ASAP7_75t_L g13643 ( 
.A(n_13166),
.B(n_12432),
.Y(n_13643)
);

AOI22xp33_ASAP7_75t_L g13644 ( 
.A1(n_13256),
.A2(n_12265),
.B1(n_12231),
.B2(n_11934),
.Y(n_13644)
);

HB1xp67_ASAP7_75t_L g13645 ( 
.A(n_12954),
.Y(n_13645)
);

NOR3xp33_ASAP7_75t_L g13646 ( 
.A(n_12998),
.B(n_11729),
.C(n_12034),
.Y(n_13646)
);

AND2x2_ASAP7_75t_L g13647 ( 
.A(n_12808),
.B(n_12452),
.Y(n_13647)
);

AND2x2_ASAP7_75t_L g13648 ( 
.A(n_12808),
.B(n_12396),
.Y(n_13648)
);

INVx1_ASAP7_75t_L g13649 ( 
.A(n_12723),
.Y(n_13649)
);

INVx2_ASAP7_75t_L g13650 ( 
.A(n_12949),
.Y(n_13650)
);

OR2x2_ASAP7_75t_L g13651 ( 
.A(n_13263),
.B(n_11185),
.Y(n_13651)
);

INVx1_ASAP7_75t_L g13652 ( 
.A(n_12729),
.Y(n_13652)
);

INVx2_ASAP7_75t_L g13653 ( 
.A(n_12959),
.Y(n_13653)
);

INVx1_ASAP7_75t_L g13654 ( 
.A(n_12729),
.Y(n_13654)
);

INVx2_ASAP7_75t_SL g13655 ( 
.A(n_13096),
.Y(n_13655)
);

INVx2_ASAP7_75t_L g13656 ( 
.A(n_12959),
.Y(n_13656)
);

OR2x2_ASAP7_75t_L g13657 ( 
.A(n_13263),
.B(n_11186),
.Y(n_13657)
);

OR2x2_ASAP7_75t_L g13658 ( 
.A(n_12629),
.B(n_11187),
.Y(n_13658)
);

AND2x2_ASAP7_75t_L g13659 ( 
.A(n_12580),
.B(n_12399),
.Y(n_13659)
);

AND2x2_ASAP7_75t_L g13660 ( 
.A(n_12584),
.B(n_12569),
.Y(n_13660)
);

OR2x2_ASAP7_75t_L g13661 ( 
.A(n_12939),
.B(n_11191),
.Y(n_13661)
);

NAND2xp5_ASAP7_75t_SL g13662 ( 
.A(n_13088),
.B(n_11846),
.Y(n_13662)
);

AND2x4_ASAP7_75t_L g13663 ( 
.A(n_12610),
.B(n_10011),
.Y(n_13663)
);

NOR2xp33_ASAP7_75t_L g13664 ( 
.A(n_12772),
.B(n_7560),
.Y(n_13664)
);

NAND2xp5_ASAP7_75t_L g13665 ( 
.A(n_12727),
.B(n_11194),
.Y(n_13665)
);

NAND2xp5_ASAP7_75t_L g13666 ( 
.A(n_12736),
.B(n_11200),
.Y(n_13666)
);

INVx2_ASAP7_75t_SL g13667 ( 
.A(n_12558),
.Y(n_13667)
);

AND2x2_ASAP7_75t_SL g13668 ( 
.A(n_13090),
.B(n_11948),
.Y(n_13668)
);

INVx2_ASAP7_75t_L g13669 ( 
.A(n_12632),
.Y(n_13669)
);

OR2x2_ASAP7_75t_L g13670 ( 
.A(n_12789),
.B(n_11201),
.Y(n_13670)
);

OR2x2_ASAP7_75t_L g13671 ( 
.A(n_13098),
.B(n_11205),
.Y(n_13671)
);

AOI22xp33_ASAP7_75t_L g13672 ( 
.A1(n_13378),
.A2(n_12337),
.B1(n_12001),
.B2(n_12358),
.Y(n_13672)
);

INVx1_ASAP7_75t_L g13673 ( 
.A(n_12730),
.Y(n_13673)
);

AND2x2_ASAP7_75t_L g13674 ( 
.A(n_12830),
.B(n_12476),
.Y(n_13674)
);

AND2x2_ASAP7_75t_L g13675 ( 
.A(n_12575),
.B(n_11207),
.Y(n_13675)
);

AND2x4_ASAP7_75t_L g13676 ( 
.A(n_12625),
.B(n_12755),
.Y(n_13676)
);

INVxp67_ASAP7_75t_SL g13677 ( 
.A(n_13301),
.Y(n_13677)
);

INVx2_ASAP7_75t_L g13678 ( 
.A(n_12642),
.Y(n_13678)
);

INVx1_ASAP7_75t_L g13679 ( 
.A(n_12730),
.Y(n_13679)
);

AND2x2_ASAP7_75t_L g13680 ( 
.A(n_12910),
.B(n_12529),
.Y(n_13680)
);

AOI22xp33_ASAP7_75t_L g13681 ( 
.A1(n_13353),
.A2(n_12269),
.B1(n_12200),
.B2(n_12180),
.Y(n_13681)
);

AND2x2_ASAP7_75t_L g13682 ( 
.A(n_12595),
.B(n_11209),
.Y(n_13682)
);

AND2x2_ASAP7_75t_L g13683 ( 
.A(n_12597),
.B(n_11212),
.Y(n_13683)
);

AND2x2_ASAP7_75t_L g13684 ( 
.A(n_12897),
.B(n_12572),
.Y(n_13684)
);

INVx1_ASAP7_75t_L g13685 ( 
.A(n_12734),
.Y(n_13685)
);

AND2x2_ASAP7_75t_L g13686 ( 
.A(n_13038),
.B(n_11215),
.Y(n_13686)
);

OR2x2_ASAP7_75t_L g13687 ( 
.A(n_13269),
.B(n_11217),
.Y(n_13687)
);

NAND2xp5_ASAP7_75t_L g13688 ( 
.A(n_12739),
.B(n_11220),
.Y(n_13688)
);

NOR2xp33_ASAP7_75t_L g13689 ( 
.A(n_12797),
.B(n_7563),
.Y(n_13689)
);

AND2x4_ASAP7_75t_SL g13690 ( 
.A(n_12642),
.B(n_6760),
.Y(n_13690)
);

CKINVDCx20_ASAP7_75t_R g13691 ( 
.A(n_13152),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_12734),
.Y(n_13692)
);

BUFx6f_ASAP7_75t_L g13693 ( 
.A(n_12759),
.Y(n_13693)
);

INVx2_ASAP7_75t_L g13694 ( 
.A(n_12748),
.Y(n_13694)
);

BUFx2_ASAP7_75t_L g13695 ( 
.A(n_12746),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_12735),
.Y(n_13696)
);

INVx1_ASAP7_75t_L g13697 ( 
.A(n_12735),
.Y(n_13697)
);

INVx2_ASAP7_75t_L g13698 ( 
.A(n_12748),
.Y(n_13698)
);

AND2x2_ASAP7_75t_L g13699 ( 
.A(n_12528),
.B(n_11223),
.Y(n_13699)
);

OAI22xp33_ASAP7_75t_L g13700 ( 
.A1(n_13187),
.A2(n_12418),
.B1(n_12446),
.B2(n_10011),
.Y(n_13700)
);

INVx2_ASAP7_75t_L g13701 ( 
.A(n_12780),
.Y(n_13701)
);

INVx1_ASAP7_75t_L g13702 ( 
.A(n_12738),
.Y(n_13702)
);

INVx1_ASAP7_75t_L g13703 ( 
.A(n_12738),
.Y(n_13703)
);

NAND2xp5_ASAP7_75t_L g13704 ( 
.A(n_12753),
.B(n_11229),
.Y(n_13704)
);

INVx1_ASAP7_75t_L g13705 ( 
.A(n_12741),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_12741),
.Y(n_13706)
);

INVx3_ASAP7_75t_L g13707 ( 
.A(n_12780),
.Y(n_13707)
);

NOR2x1_ASAP7_75t_L g13708 ( 
.A(n_13249),
.B(n_12380),
.Y(n_13708)
);

INVx2_ASAP7_75t_L g13709 ( 
.A(n_12765),
.Y(n_13709)
);

AND2x2_ASAP7_75t_L g13710 ( 
.A(n_12557),
.B(n_12934),
.Y(n_13710)
);

AND2x2_ASAP7_75t_L g13711 ( 
.A(n_12958),
.B(n_11231),
.Y(n_13711)
);

INVx1_ASAP7_75t_L g13712 ( 
.A(n_12756),
.Y(n_13712)
);

INVx2_ASAP7_75t_L g13713 ( 
.A(n_12771),
.Y(n_13713)
);

INVx2_ASAP7_75t_L g13714 ( 
.A(n_12777),
.Y(n_13714)
);

NAND2xp5_ASAP7_75t_L g13715 ( 
.A(n_12773),
.B(n_11234),
.Y(n_13715)
);

OR2x2_ASAP7_75t_L g13716 ( 
.A(n_13233),
.B(n_11235),
.Y(n_13716)
);

AND2x2_ASAP7_75t_L g13717 ( 
.A(n_13030),
.B(n_11236),
.Y(n_13717)
);

AND2x2_ASAP7_75t_L g13718 ( 
.A(n_12833),
.B(n_11238),
.Y(n_13718)
);

INVx2_ASAP7_75t_L g13719 ( 
.A(n_12869),
.Y(n_13719)
);

AND2x4_ASAP7_75t_L g13720 ( 
.A(n_12764),
.B(n_10011),
.Y(n_13720)
);

AND2x4_ASAP7_75t_L g13721 ( 
.A(n_12782),
.B(n_10037),
.Y(n_13721)
);

INVx1_ASAP7_75t_L g13722 ( 
.A(n_12756),
.Y(n_13722)
);

NAND2xp5_ASAP7_75t_L g13723 ( 
.A(n_12781),
.B(n_11240),
.Y(n_13723)
);

OR2x2_ASAP7_75t_L g13724 ( 
.A(n_12600),
.B(n_11251),
.Y(n_13724)
);

AND2x2_ASAP7_75t_L g13725 ( 
.A(n_12656),
.B(n_11256),
.Y(n_13725)
);

AND2x2_ASAP7_75t_L g13726 ( 
.A(n_12834),
.B(n_12927),
.Y(n_13726)
);

AND2x2_ASAP7_75t_L g13727 ( 
.A(n_12684),
.B(n_11264),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_12762),
.Y(n_13728)
);

INVx2_ASAP7_75t_L g13729 ( 
.A(n_12869),
.Y(n_13729)
);

INVx4_ASAP7_75t_L g13730 ( 
.A(n_12998),
.Y(n_13730)
);

AOI22xp33_ASAP7_75t_SL g13731 ( 
.A1(n_13353),
.A2(n_11867),
.B1(n_11970),
.B2(n_11931),
.Y(n_13731)
);

AND2x4_ASAP7_75t_L g13732 ( 
.A(n_12786),
.B(n_10037),
.Y(n_13732)
);

INVx2_ASAP7_75t_L g13733 ( 
.A(n_12911),
.Y(n_13733)
);

NOR2xp67_ASAP7_75t_L g13734 ( 
.A(n_13301),
.B(n_11265),
.Y(n_13734)
);

AND2x2_ASAP7_75t_L g13735 ( 
.A(n_12947),
.B(n_11270),
.Y(n_13735)
);

AND2x4_ASAP7_75t_L g13736 ( 
.A(n_12787),
.B(n_10037),
.Y(n_13736)
);

INVx2_ASAP7_75t_L g13737 ( 
.A(n_12911),
.Y(n_13737)
);

INVx1_ASAP7_75t_L g13738 ( 
.A(n_12762),
.Y(n_13738)
);

NAND2xp5_ASAP7_75t_L g13739 ( 
.A(n_13032),
.B(n_11278),
.Y(n_13739)
);

INVx1_ASAP7_75t_L g13740 ( 
.A(n_12763),
.Y(n_13740)
);

NAND2xp5_ASAP7_75t_L g13741 ( 
.A(n_12843),
.B(n_11279),
.Y(n_13741)
);

NAND2xp5_ASAP7_75t_L g13742 ( 
.A(n_12847),
.B(n_11283),
.Y(n_13742)
);

INVx2_ASAP7_75t_L g13743 ( 
.A(n_12793),
.Y(n_13743)
);

AND2x2_ASAP7_75t_L g13744 ( 
.A(n_12905),
.B(n_11287),
.Y(n_13744)
);

NAND2xp5_ASAP7_75t_L g13745 ( 
.A(n_12863),
.B(n_11292),
.Y(n_13745)
);

INVx2_ASAP7_75t_SL g13746 ( 
.A(n_12864),
.Y(n_13746)
);

INVx3_ASAP7_75t_L g13747 ( 
.A(n_12800),
.Y(n_13747)
);

INVx2_ASAP7_75t_L g13748 ( 
.A(n_12695),
.Y(n_13748)
);

OR2x2_ASAP7_75t_L g13749 ( 
.A(n_13254),
.B(n_11296),
.Y(n_13749)
);

INVx2_ASAP7_75t_L g13750 ( 
.A(n_12695),
.Y(n_13750)
);

INVx1_ASAP7_75t_L g13751 ( 
.A(n_12763),
.Y(n_13751)
);

INVx1_ASAP7_75t_L g13752 ( 
.A(n_12768),
.Y(n_13752)
);

INVx2_ASAP7_75t_L g13753 ( 
.A(n_12608),
.Y(n_13753)
);

NAND2xp5_ASAP7_75t_L g13754 ( 
.A(n_12867),
.B(n_11298),
.Y(n_13754)
);

AND2x2_ASAP7_75t_L g13755 ( 
.A(n_12605),
.B(n_11299),
.Y(n_13755)
);

AND2x4_ASAP7_75t_L g13756 ( 
.A(n_12619),
.B(n_10037),
.Y(n_13756)
);

BUFx2_ASAP7_75t_L g13757 ( 
.A(n_12671),
.Y(n_13757)
);

AND2x2_ASAP7_75t_L g13758 ( 
.A(n_12609),
.B(n_11300),
.Y(n_13758)
);

NAND2xp5_ASAP7_75t_L g13759 ( 
.A(n_12885),
.B(n_11304),
.Y(n_13759)
);

AND2x2_ASAP7_75t_L g13760 ( 
.A(n_12612),
.B(n_11308),
.Y(n_13760)
);

BUFx2_ASAP7_75t_L g13761 ( 
.A(n_13266),
.Y(n_13761)
);

NAND2xp5_ASAP7_75t_L g13762 ( 
.A(n_12896),
.B(n_11311),
.Y(n_13762)
);

INVx1_ASAP7_75t_L g13763 ( 
.A(n_12768),
.Y(n_13763)
);

INVx2_ASAP7_75t_L g13764 ( 
.A(n_12620),
.Y(n_13764)
);

AND2x2_ASAP7_75t_L g13765 ( 
.A(n_12614),
.B(n_11320),
.Y(n_13765)
);

INVx1_ASAP7_75t_L g13766 ( 
.A(n_12770),
.Y(n_13766)
);

AND2x2_ASAP7_75t_L g13767 ( 
.A(n_12835),
.B(n_11325),
.Y(n_13767)
);

INVx3_ASAP7_75t_L g13768 ( 
.A(n_12800),
.Y(n_13768)
);

NAND2x1p5_ASAP7_75t_L g13769 ( 
.A(n_12703),
.B(n_10037),
.Y(n_13769)
);

INVx2_ASAP7_75t_L g13770 ( 
.A(n_13086),
.Y(n_13770)
);

AND2x2_ASAP7_75t_L g13771 ( 
.A(n_12916),
.B(n_11333),
.Y(n_13771)
);

INVx1_ASAP7_75t_L g13772 ( 
.A(n_12770),
.Y(n_13772)
);

HB1xp67_ASAP7_75t_L g13773 ( 
.A(n_12627),
.Y(n_13773)
);

INVx1_ASAP7_75t_L g13774 ( 
.A(n_12790),
.Y(n_13774)
);

OR2x2_ASAP7_75t_L g13775 ( 
.A(n_13056),
.B(n_11335),
.Y(n_13775)
);

INVx1_ASAP7_75t_L g13776 ( 
.A(n_13026),
.Y(n_13776)
);

NAND2xp5_ASAP7_75t_L g13777 ( 
.A(n_12900),
.B(n_11341),
.Y(n_13777)
);

AND2x2_ASAP7_75t_L g13778 ( 
.A(n_12841),
.B(n_13018),
.Y(n_13778)
);

NAND2xp5_ASAP7_75t_L g13779 ( 
.A(n_12902),
.B(n_11343),
.Y(n_13779)
);

NAND2xp5_ASAP7_75t_L g13780 ( 
.A(n_13247),
.B(n_11344),
.Y(n_13780)
);

AND2x2_ASAP7_75t_L g13781 ( 
.A(n_12744),
.B(n_11348),
.Y(n_13781)
);

INVx1_ASAP7_75t_L g13782 ( 
.A(n_12635),
.Y(n_13782)
);

AOI22xp33_ASAP7_75t_SL g13783 ( 
.A1(n_13315),
.A2(n_12290),
.B1(n_11039),
.B2(n_12169),
.Y(n_13783)
);

INVx1_ASAP7_75t_L g13784 ( 
.A(n_12641),
.Y(n_13784)
);

HB1xp67_ASAP7_75t_L g13785 ( 
.A(n_12634),
.Y(n_13785)
);

AND2x2_ASAP7_75t_L g13786 ( 
.A(n_12749),
.B(n_12810),
.Y(n_13786)
);

NAND2xp5_ASAP7_75t_SL g13787 ( 
.A(n_13315),
.B(n_12106),
.Y(n_13787)
);

AND2x2_ASAP7_75t_L g13788 ( 
.A(n_12815),
.B(n_11356),
.Y(n_13788)
);

AOI22xp33_ASAP7_75t_SL g13789 ( 
.A1(n_13180),
.A2(n_11039),
.B1(n_9303),
.B2(n_8015),
.Y(n_13789)
);

HB1xp67_ASAP7_75t_L g13790 ( 
.A(n_13149),
.Y(n_13790)
);

OAI221xp5_ASAP7_75t_SL g13791 ( 
.A1(n_13231),
.A2(n_12437),
.B1(n_12325),
.B2(n_12309),
.C(n_12428),
.Y(n_13791)
);

AND2x2_ASAP7_75t_L g13792 ( 
.A(n_12822),
.B(n_11362),
.Y(n_13792)
);

INVx4_ASAP7_75t_L g13793 ( 
.A(n_12968),
.Y(n_13793)
);

AND2x2_ASAP7_75t_L g13794 ( 
.A(n_12842),
.B(n_11363),
.Y(n_13794)
);

INVx2_ASAP7_75t_L g13795 ( 
.A(n_13086),
.Y(n_13795)
);

AND2x2_ASAP7_75t_L g13796 ( 
.A(n_13015),
.B(n_11367),
.Y(n_13796)
);

INVx3_ASAP7_75t_L g13797 ( 
.A(n_12803),
.Y(n_13797)
);

AND2x2_ASAP7_75t_L g13798 ( 
.A(n_13260),
.B(n_11371),
.Y(n_13798)
);

INVxp67_ASAP7_75t_L g13799 ( 
.A(n_12844),
.Y(n_13799)
);

INVxp67_ASAP7_75t_SL g13800 ( 
.A(n_13363),
.Y(n_13800)
);

OAI22xp5_ASAP7_75t_L g13801 ( 
.A1(n_12837),
.A2(n_13247),
.B1(n_13312),
.B2(n_13316),
.Y(n_13801)
);

NOR2xp67_ASAP7_75t_L g13802 ( 
.A(n_13219),
.B(n_11373),
.Y(n_13802)
);

INVx2_ASAP7_75t_L g13803 ( 
.A(n_13086),
.Y(n_13803)
);

HB1xp67_ASAP7_75t_L g13804 ( 
.A(n_13149),
.Y(n_13804)
);

INVx3_ASAP7_75t_L g13805 ( 
.A(n_12803),
.Y(n_13805)
);

INVx1_ASAP7_75t_L g13806 ( 
.A(n_12643),
.Y(n_13806)
);

NAND2xp5_ASAP7_75t_L g13807 ( 
.A(n_13279),
.B(n_11374),
.Y(n_13807)
);

INVx1_ASAP7_75t_L g13808 ( 
.A(n_12644),
.Y(n_13808)
);

INVx3_ASAP7_75t_L g13809 ( 
.A(n_12895),
.Y(n_13809)
);

INVx1_ASAP7_75t_L g13810 ( 
.A(n_12646),
.Y(n_13810)
);

AOI22xp33_ASAP7_75t_L g13811 ( 
.A1(n_13125),
.A2(n_12170),
.B1(n_11997),
.B2(n_12121),
.Y(n_13811)
);

INVx2_ASAP7_75t_SL g13812 ( 
.A(n_12792),
.Y(n_13812)
);

INVx1_ASAP7_75t_L g13813 ( 
.A(n_12651),
.Y(n_13813)
);

AND2x2_ASAP7_75t_L g13814 ( 
.A(n_12795),
.B(n_11376),
.Y(n_13814)
);

AND2x2_ASAP7_75t_L g13815 ( 
.A(n_12796),
.B(n_11380),
.Y(n_13815)
);

NAND2xp5_ASAP7_75t_L g13816 ( 
.A(n_13226),
.B(n_11384),
.Y(n_13816)
);

INVx1_ASAP7_75t_L g13817 ( 
.A(n_12661),
.Y(n_13817)
);

BUFx3_ASAP7_75t_L g13818 ( 
.A(n_12924),
.Y(n_13818)
);

INVx2_ASAP7_75t_L g13819 ( 
.A(n_12895),
.Y(n_13819)
);

NAND2xp5_ASAP7_75t_L g13820 ( 
.A(n_13226),
.B(n_13072),
.Y(n_13820)
);

HB1xp67_ASAP7_75t_L g13821 ( 
.A(n_13149),
.Y(n_13821)
);

INVx1_ASAP7_75t_L g13822 ( 
.A(n_12662),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_12802),
.B(n_11386),
.Y(n_13823)
);

INVx1_ASAP7_75t_L g13824 ( 
.A(n_12665),
.Y(n_13824)
);

NOR2x1_ASAP7_75t_SL g13825 ( 
.A(n_13422),
.B(n_10037),
.Y(n_13825)
);

INVx1_ASAP7_75t_L g13826 ( 
.A(n_12668),
.Y(n_13826)
);

NOR2xp33_ASAP7_75t_L g13827 ( 
.A(n_13064),
.B(n_7593),
.Y(n_13827)
);

INVx2_ASAP7_75t_L g13828 ( 
.A(n_13041),
.Y(n_13828)
);

BUFx3_ASAP7_75t_L g13829 ( 
.A(n_12769),
.Y(n_13829)
);

HB1xp67_ASAP7_75t_L g13830 ( 
.A(n_13009),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_12670),
.Y(n_13831)
);

AND2x2_ASAP7_75t_L g13832 ( 
.A(n_13039),
.B(n_13083),
.Y(n_13832)
);

OR2x2_ASAP7_75t_L g13833 ( 
.A(n_13267),
.B(n_11388),
.Y(n_13833)
);

INVx1_ASAP7_75t_L g13834 ( 
.A(n_12672),
.Y(n_13834)
);

INVx1_ASAP7_75t_L g13835 ( 
.A(n_12676),
.Y(n_13835)
);

OR2x2_ASAP7_75t_L g13836 ( 
.A(n_13375),
.B(n_11390),
.Y(n_13836)
);

NOR2xp33_ASAP7_75t_L g13837 ( 
.A(n_12936),
.B(n_12442),
.Y(n_13837)
);

INVx1_ASAP7_75t_L g13838 ( 
.A(n_12680),
.Y(n_13838)
);

OR2x2_ASAP7_75t_L g13839 ( 
.A(n_13029),
.B(n_11394),
.Y(n_13839)
);

OR2x2_ASAP7_75t_L g13840 ( 
.A(n_12851),
.B(n_11398),
.Y(n_13840)
);

NAND2xp5_ASAP7_75t_L g13841 ( 
.A(n_12912),
.B(n_11404),
.Y(n_13841)
);

AND2x2_ASAP7_75t_L g13842 ( 
.A(n_12918),
.B(n_11407),
.Y(n_13842)
);

AND2x2_ASAP7_75t_L g13843 ( 
.A(n_12904),
.B(n_11410),
.Y(n_13843)
);

INVx2_ASAP7_75t_L g13844 ( 
.A(n_13041),
.Y(n_13844)
);

INVx1_ASAP7_75t_L g13845 ( 
.A(n_12686),
.Y(n_13845)
);

BUFx2_ASAP7_75t_L g13846 ( 
.A(n_13273),
.Y(n_13846)
);

INVxp67_ASAP7_75t_L g13847 ( 
.A(n_13191),
.Y(n_13847)
);

INVxp67_ASAP7_75t_L g13848 ( 
.A(n_13219),
.Y(n_13848)
);

OR2x2_ASAP7_75t_L g13849 ( 
.A(n_13243),
.B(n_11413),
.Y(n_13849)
);

INVx1_ASAP7_75t_L g13850 ( 
.A(n_12689),
.Y(n_13850)
);

AND2x2_ASAP7_75t_L g13851 ( 
.A(n_13188),
.B(n_11414),
.Y(n_13851)
);

BUFx2_ASAP7_75t_L g13852 ( 
.A(n_13273),
.Y(n_13852)
);

AOI22xp33_ASAP7_75t_L g13853 ( 
.A1(n_13257),
.A2(n_11894),
.B1(n_12142),
.B2(n_12040),
.Y(n_13853)
);

AND2x2_ASAP7_75t_L g13854 ( 
.A(n_12784),
.B(n_11415),
.Y(n_13854)
);

AND2x2_ASAP7_75t_L g13855 ( 
.A(n_12816),
.B(n_12848),
.Y(n_13855)
);

NAND2xp5_ASAP7_75t_L g13856 ( 
.A(n_12548),
.B(n_11418),
.Y(n_13856)
);

AND2x2_ASAP7_75t_L g13857 ( 
.A(n_12884),
.B(n_11427),
.Y(n_13857)
);

OR2x2_ASAP7_75t_L g13858 ( 
.A(n_12860),
.B(n_11428),
.Y(n_13858)
);

INVx1_ASAP7_75t_L g13859 ( 
.A(n_12691),
.Y(n_13859)
);

BUFx3_ASAP7_75t_L g13860 ( 
.A(n_12926),
.Y(n_13860)
);

BUFx6f_ASAP7_75t_L g13861 ( 
.A(n_12555),
.Y(n_13861)
);

OR2x2_ASAP7_75t_L g13862 ( 
.A(n_13290),
.B(n_11430),
.Y(n_13862)
);

INVx2_ASAP7_75t_L g13863 ( 
.A(n_13053),
.Y(n_13863)
);

NOR2xp33_ASAP7_75t_SL g13864 ( 
.A(n_12628),
.B(n_12946),
.Y(n_13864)
);

AOI22xp33_ASAP7_75t_L g13865 ( 
.A1(n_13329),
.A2(n_12140),
.B1(n_12135),
.B2(n_12071),
.Y(n_13865)
);

INVx2_ASAP7_75t_L g13866 ( 
.A(n_13053),
.Y(n_13866)
);

INVx1_ASAP7_75t_L g13867 ( 
.A(n_12692),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_12694),
.Y(n_13868)
);

INVx1_ASAP7_75t_L g13869 ( 
.A(n_12699),
.Y(n_13869)
);

AND2x2_ASAP7_75t_L g13870 ( 
.A(n_12570),
.B(n_11431),
.Y(n_13870)
);

AND2x2_ASAP7_75t_L g13871 ( 
.A(n_12825),
.B(n_11440),
.Y(n_13871)
);

INVx1_ASAP7_75t_L g13872 ( 
.A(n_12706),
.Y(n_13872)
);

OR2x2_ASAP7_75t_L g13873 ( 
.A(n_12948),
.B(n_11449),
.Y(n_13873)
);

AND2x2_ASAP7_75t_L g13874 ( 
.A(n_13200),
.B(n_11450),
.Y(n_13874)
);

AND2x2_ASAP7_75t_L g13875 ( 
.A(n_13304),
.B(n_11452),
.Y(n_13875)
);

INVxp67_ASAP7_75t_L g13876 ( 
.A(n_13133),
.Y(n_13876)
);

BUFx2_ASAP7_75t_L g13877 ( 
.A(n_13423),
.Y(n_13877)
);

HB1xp67_ASAP7_75t_L g13878 ( 
.A(n_13023),
.Y(n_13878)
);

AND2x2_ASAP7_75t_L g13879 ( 
.A(n_13304),
.B(n_11454),
.Y(n_13879)
);

INVx2_ASAP7_75t_L g13880 ( 
.A(n_13070),
.Y(n_13880)
);

HB1xp67_ASAP7_75t_L g13881 ( 
.A(n_13035),
.Y(n_13881)
);

NAND2xp5_ASAP7_75t_L g13882 ( 
.A(n_13168),
.B(n_11455),
.Y(n_13882)
);

AND2x2_ASAP7_75t_L g13883 ( 
.A(n_13308),
.B(n_11459),
.Y(n_13883)
);

OR2x2_ASAP7_75t_L g13884 ( 
.A(n_13259),
.B(n_11462),
.Y(n_13884)
);

AND2x2_ASAP7_75t_L g13885 ( 
.A(n_13308),
.B(n_11470),
.Y(n_13885)
);

AND2x2_ASAP7_75t_L g13886 ( 
.A(n_13335),
.B(n_11481),
.Y(n_13886)
);

OR2x2_ASAP7_75t_L g13887 ( 
.A(n_13259),
.B(n_11482),
.Y(n_13887)
);

INVxp67_ASAP7_75t_SL g13888 ( 
.A(n_12750),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13335),
.B(n_11486),
.Y(n_13889)
);

INVx1_ASAP7_75t_L g13890 ( 
.A(n_12714),
.Y(n_13890)
);

INVx1_ASAP7_75t_L g13891 ( 
.A(n_12717),
.Y(n_13891)
);

OAI221xp5_ASAP7_75t_SL g13892 ( 
.A1(n_13373),
.A2(n_12424),
.B1(n_12406),
.B2(n_12387),
.C(n_12103),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_12718),
.Y(n_13893)
);

NOR2x1_ASAP7_75t_L g13894 ( 
.A(n_13115),
.B(n_12045),
.Y(n_13894)
);

AND2x2_ASAP7_75t_L g13895 ( 
.A(n_13077),
.B(n_11487),
.Y(n_13895)
);

BUFx2_ASAP7_75t_L g13896 ( 
.A(n_13428),
.Y(n_13896)
);

INVxp67_ASAP7_75t_SL g13897 ( 
.A(n_13271),
.Y(n_13897)
);

INVx1_ASAP7_75t_L g13898 ( 
.A(n_12774),
.Y(n_13898)
);

OR2x2_ASAP7_75t_L g13899 ( 
.A(n_13339),
.B(n_13150),
.Y(n_13899)
);

AND2x2_ASAP7_75t_L g13900 ( 
.A(n_13358),
.B(n_11489),
.Y(n_13900)
);

INVx1_ASAP7_75t_L g13901 ( 
.A(n_12775),
.Y(n_13901)
);

INVx2_ASAP7_75t_L g13902 ( 
.A(n_13070),
.Y(n_13902)
);

HB1xp67_ASAP7_75t_L g13903 ( 
.A(n_13068),
.Y(n_13903)
);

HB1xp67_ASAP7_75t_L g13904 ( 
.A(n_13042),
.Y(n_13904)
);

AND2x2_ASAP7_75t_L g13905 ( 
.A(n_13222),
.B(n_11491),
.Y(n_13905)
);

OR2x2_ASAP7_75t_L g13906 ( 
.A(n_13296),
.B(n_11492),
.Y(n_13906)
);

INVx1_ASAP7_75t_L g13907 ( 
.A(n_12776),
.Y(n_13907)
);

OAI21xp33_ASAP7_75t_L g13908 ( 
.A1(n_13356),
.A2(n_11496),
.B(n_11493),
.Y(n_13908)
);

AND2x2_ASAP7_75t_L g13909 ( 
.A(n_13043),
.B(n_12922),
.Y(n_13909)
);

INVx1_ASAP7_75t_SL g13910 ( 
.A(n_13240),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_12925),
.B(n_11499),
.Y(n_13911)
);

AOI22xp33_ASAP7_75t_L g13912 ( 
.A1(n_13329),
.A2(n_12076),
.B1(n_8015),
.B2(n_10277),
.Y(n_13912)
);

AND2x4_ASAP7_75t_L g13913 ( 
.A(n_12732),
.B(n_10234),
.Y(n_13913)
);

NAND2xp5_ASAP7_75t_L g13914 ( 
.A(n_13405),
.B(n_11501),
.Y(n_13914)
);

INVx1_ASAP7_75t_L g13915 ( 
.A(n_12779),
.Y(n_13915)
);

INVx1_ASAP7_75t_L g13916 ( 
.A(n_12783),
.Y(n_13916)
);

AND2x2_ASAP7_75t_L g13917 ( 
.A(n_13208),
.B(n_11502),
.Y(n_13917)
);

NAND2x1_ASAP7_75t_L g13918 ( 
.A(n_13427),
.B(n_10452),
.Y(n_13918)
);

NAND2xp5_ASAP7_75t_L g13919 ( 
.A(n_13411),
.B(n_11506),
.Y(n_13919)
);

INVx2_ASAP7_75t_L g13920 ( 
.A(n_12917),
.Y(n_13920)
);

NAND2xp5_ASAP7_75t_SL g13921 ( 
.A(n_13058),
.B(n_12807),
.Y(n_13921)
);

AND2x4_ASAP7_75t_L g13922 ( 
.A(n_12742),
.B(n_10234),
.Y(n_13922)
);

AND2x2_ASAP7_75t_L g13923 ( 
.A(n_13317),
.B(n_11512),
.Y(n_13923)
);

AND2x2_ASAP7_75t_L g13924 ( 
.A(n_13317),
.B(n_11513),
.Y(n_13924)
);

NOR2xp33_ASAP7_75t_L g13925 ( 
.A(n_13238),
.B(n_11517),
.Y(n_13925)
);

BUFx2_ASAP7_75t_L g13926 ( 
.A(n_12752),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_12791),
.Y(n_13927)
);

AND2x2_ASAP7_75t_L g13928 ( 
.A(n_13354),
.B(n_11523),
.Y(n_13928)
);

INVx1_ASAP7_75t_L g13929 ( 
.A(n_12798),
.Y(n_13929)
);

AND2x2_ASAP7_75t_L g13930 ( 
.A(n_12985),
.B(n_11525),
.Y(n_13930)
);

INVx1_ASAP7_75t_L g13931 ( 
.A(n_12799),
.Y(n_13931)
);

INVx2_ASAP7_75t_L g13932 ( 
.A(n_12917),
.Y(n_13932)
);

AND2x2_ASAP7_75t_L g13933 ( 
.A(n_13221),
.B(n_11533),
.Y(n_13933)
);

AND2x4_ASAP7_75t_L g13934 ( 
.A(n_12566),
.B(n_10234),
.Y(n_13934)
);

AND2x2_ASAP7_75t_L g13935 ( 
.A(n_12929),
.B(n_11537),
.Y(n_13935)
);

AND2x4_ASAP7_75t_L g13936 ( 
.A(n_12579),
.B(n_12581),
.Y(n_13936)
);

OR2x2_ASAP7_75t_L g13937 ( 
.A(n_13107),
.B(n_6894),
.Y(n_13937)
);

NAND2xp5_ASAP7_75t_L g13938 ( 
.A(n_13346),
.B(n_8316),
.Y(n_13938)
);

OAI22xp5_ASAP7_75t_L g13939 ( 
.A1(n_13365),
.A2(n_8953),
.B1(n_10277),
.B2(n_10234),
.Y(n_13939)
);

AND2x4_ASAP7_75t_L g13940 ( 
.A(n_12582),
.B(n_10234),
.Y(n_13940)
);

INVx2_ASAP7_75t_L g13941 ( 
.A(n_12740),
.Y(n_13941)
);

OR2x2_ASAP7_75t_L g13942 ( 
.A(n_13172),
.B(n_6927),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_12862),
.B(n_10234),
.Y(n_13943)
);

INVx2_ASAP7_75t_L g13944 ( 
.A(n_12767),
.Y(n_13944)
);

OAI22xp5_ASAP7_75t_L g13945 ( 
.A1(n_13205),
.A2(n_8953),
.B1(n_10378),
.B2(n_10277),
.Y(n_13945)
);

AND2x2_ASAP7_75t_L g13946 ( 
.A(n_13183),
.B(n_10277),
.Y(n_13946)
);

INVx1_ASAP7_75t_L g13947 ( 
.A(n_12811),
.Y(n_13947)
);

AND2x2_ASAP7_75t_L g13948 ( 
.A(n_13184),
.B(n_10277),
.Y(n_13948)
);

AND2x2_ASAP7_75t_L g13949 ( 
.A(n_12935),
.B(n_10277),
.Y(n_13949)
);

NAND2xp5_ASAP7_75t_L g13950 ( 
.A(n_13264),
.B(n_8328),
.Y(n_13950)
);

NAND2xp5_ASAP7_75t_L g13951 ( 
.A(n_13253),
.B(n_8337),
.Y(n_13951)
);

INVx2_ASAP7_75t_L g13952 ( 
.A(n_12801),
.Y(n_13952)
);

INVx1_ASAP7_75t_L g13953 ( 
.A(n_12817),
.Y(n_13953)
);

INVx2_ASAP7_75t_L g13954 ( 
.A(n_13076),
.Y(n_13954)
);

OR2x2_ASAP7_75t_L g13955 ( 
.A(n_13245),
.B(n_6927),
.Y(n_13955)
);

INVx2_ASAP7_75t_L g13956 ( 
.A(n_13076),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_12821),
.Y(n_13957)
);

INVx1_ASAP7_75t_L g13958 ( 
.A(n_12826),
.Y(n_13958)
);

INVxp67_ASAP7_75t_SL g13959 ( 
.A(n_12969),
.Y(n_13959)
);

INVx1_ASAP7_75t_L g13960 ( 
.A(n_12829),
.Y(n_13960)
);

OAI22xp5_ASAP7_75t_L g13961 ( 
.A1(n_13439),
.A2(n_10378),
.B1(n_7732),
.B2(n_7792),
.Y(n_13961)
);

INVx2_ASAP7_75t_L g13962 ( 
.A(n_12652),
.Y(n_13962)
);

OR2x2_ASAP7_75t_L g13963 ( 
.A(n_12866),
.B(n_8337),
.Y(n_13963)
);

NAND2xp5_ASAP7_75t_L g13964 ( 
.A(n_13103),
.B(n_13345),
.Y(n_13964)
);

AOI22xp33_ASAP7_75t_L g13965 ( 
.A1(n_13439),
.A2(n_8015),
.B1(n_10378),
.B2(n_9303),
.Y(n_13965)
);

INVx1_ASAP7_75t_L g13966 ( 
.A(n_12831),
.Y(n_13966)
);

AND2x4_ASAP7_75t_L g13967 ( 
.A(n_12587),
.B(n_10378),
.Y(n_13967)
);

INVxp67_ASAP7_75t_SL g13968 ( 
.A(n_12987),
.Y(n_13968)
);

AOI22xp33_ASAP7_75t_L g13969 ( 
.A1(n_13345),
.A2(n_8015),
.B1(n_10378),
.B2(n_9303),
.Y(n_13969)
);

INVx3_ASAP7_75t_L g13970 ( 
.A(n_12792),
.Y(n_13970)
);

INVxp67_ASAP7_75t_L g13971 ( 
.A(n_13421),
.Y(n_13971)
);

INVx3_ASAP7_75t_L g13972 ( 
.A(n_12983),
.Y(n_13972)
);

INVx1_ASAP7_75t_L g13973 ( 
.A(n_12846),
.Y(n_13973)
);

INVx2_ASAP7_75t_L g13974 ( 
.A(n_12667),
.Y(n_13974)
);

AND2x2_ASAP7_75t_L g13975 ( 
.A(n_12988),
.B(n_10378),
.Y(n_13975)
);

OR2x2_ASAP7_75t_L g13976 ( 
.A(n_13359),
.B(n_8413),
.Y(n_13976)
);

BUFx6f_ASAP7_75t_L g13977 ( 
.A(n_12593),
.Y(n_13977)
);

BUFx3_ASAP7_75t_L g13978 ( 
.A(n_12857),
.Y(n_13978)
);

AND2x2_ASAP7_75t_L g13979 ( 
.A(n_13309),
.B(n_7731),
.Y(n_13979)
);

AOI221xp5_ASAP7_75t_L g13980 ( 
.A1(n_13356),
.A2(n_9209),
.B1(n_9215),
.B2(n_9195),
.C(n_9189),
.Y(n_13980)
);

OAI22xp5_ASAP7_75t_L g13981 ( 
.A1(n_13336),
.A2(n_7732),
.B1(n_7792),
.B2(n_7749),
.Y(n_13981)
);

NOR2xp33_ASAP7_75t_L g13982 ( 
.A(n_12898),
.B(n_8413),
.Y(n_13982)
);

INVx1_ASAP7_75t_L g13983 ( 
.A(n_12850),
.Y(n_13983)
);

NAND2xp5_ASAP7_75t_L g13984 ( 
.A(n_13199),
.B(n_8474),
.Y(n_13984)
);

HB1xp67_ASAP7_75t_L g13985 ( 
.A(n_13050),
.Y(n_13985)
);

INVx1_ASAP7_75t_L g13986 ( 
.A(n_12861),
.Y(n_13986)
);

OR2x2_ASAP7_75t_L g13987 ( 
.A(n_12875),
.B(n_8474),
.Y(n_13987)
);

NAND2x1_ASAP7_75t_L g13988 ( 
.A(n_13412),
.B(n_10452),
.Y(n_13988)
);

INVx1_ASAP7_75t_L g13989 ( 
.A(n_12865),
.Y(n_13989)
);

AND2x4_ASAP7_75t_L g13990 ( 
.A(n_12598),
.B(n_10770),
.Y(n_13990)
);

INVx1_ASAP7_75t_SL g13991 ( 
.A(n_13388),
.Y(n_13991)
);

AND2x2_ASAP7_75t_L g13992 ( 
.A(n_12994),
.B(n_7731),
.Y(n_13992)
);

INVx2_ASAP7_75t_L g13993 ( 
.A(n_12677),
.Y(n_13993)
);

INVx2_ASAP7_75t_L g13994 ( 
.A(n_12678),
.Y(n_13994)
);

OR2x2_ASAP7_75t_L g13995 ( 
.A(n_13420),
.B(n_9351),
.Y(n_13995)
);

HB1xp67_ASAP7_75t_L g13996 ( 
.A(n_13280),
.Y(n_13996)
);

AND2x4_ASAP7_75t_L g13997 ( 
.A(n_12636),
.B(n_10543),
.Y(n_13997)
);

INVx2_ASAP7_75t_SL g13998 ( 
.A(n_12845),
.Y(n_13998)
);

NOR2xp67_ASAP7_75t_SL g13999 ( 
.A(n_13116),
.B(n_8282),
.Y(n_13999)
);

AND2x4_ASAP7_75t_L g14000 ( 
.A(n_12650),
.B(n_10689),
.Y(n_14000)
);

INVx1_ASAP7_75t_L g14001 ( 
.A(n_12871),
.Y(n_14001)
);

INVxp67_ASAP7_75t_SL g14002 ( 
.A(n_12530),
.Y(n_14002)
);

AND2x2_ASAP7_75t_L g14003 ( 
.A(n_13176),
.B(n_7731),
.Y(n_14003)
);

BUFx2_ASAP7_75t_L g14004 ( 
.A(n_13440),
.Y(n_14004)
);

INVx1_ASAP7_75t_L g14005 ( 
.A(n_12873),
.Y(n_14005)
);

INVx2_ASAP7_75t_L g14006 ( 
.A(n_12681),
.Y(n_14006)
);

AND2x4_ASAP7_75t_SL g14007 ( 
.A(n_13073),
.B(n_6760),
.Y(n_14007)
);

INVx1_ASAP7_75t_L g14008 ( 
.A(n_12874),
.Y(n_14008)
);

AND2x2_ASAP7_75t_L g14009 ( 
.A(n_12894),
.B(n_7752),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_12876),
.Y(n_14010)
);

AND2x2_ASAP7_75t_L g14011 ( 
.A(n_13060),
.B(n_7752),
.Y(n_14011)
);

OR2x2_ASAP7_75t_L g14012 ( 
.A(n_13324),
.B(n_13277),
.Y(n_14012)
);

AND2x2_ASAP7_75t_L g14013 ( 
.A(n_12640),
.B(n_7765),
.Y(n_14013)
);

OR2x2_ASAP7_75t_L g14014 ( 
.A(n_13277),
.B(n_9351),
.Y(n_14014)
);

NAND2xp5_ASAP7_75t_L g14015 ( 
.A(n_13440),
.B(n_9783),
.Y(n_14015)
);

NAND2xp5_ASAP7_75t_L g14016 ( 
.A(n_13323),
.B(n_9785),
.Y(n_14016)
);

CKINVDCx14_ASAP7_75t_R g14017 ( 
.A(n_13215),
.Y(n_14017)
);

INVx2_ASAP7_75t_L g14018 ( 
.A(n_12688),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_12973),
.B(n_7765),
.Y(n_14019)
);

AND2x2_ASAP7_75t_L g14020 ( 
.A(n_13377),
.B(n_7826),
.Y(n_14020)
);

OR2x2_ASAP7_75t_L g14021 ( 
.A(n_12852),
.B(n_9351),
.Y(n_14021)
);

AOI22xp33_ASAP7_75t_L g14022 ( 
.A1(n_13361),
.A2(n_8015),
.B1(n_9303),
.B2(n_8036),
.Y(n_14022)
);

NAND2xp5_ASAP7_75t_L g14023 ( 
.A(n_13323),
.B(n_9785),
.Y(n_14023)
);

AND2x2_ASAP7_75t_L g14024 ( 
.A(n_13390),
.B(n_7826),
.Y(n_14024)
);

AND2x2_ASAP7_75t_L g14025 ( 
.A(n_13391),
.B(n_7827),
.Y(n_14025)
);

INVx2_ASAP7_75t_L g14026 ( 
.A(n_12693),
.Y(n_14026)
);

INVx1_ASAP7_75t_L g14027 ( 
.A(n_12880),
.Y(n_14027)
);

AND2x2_ASAP7_75t_L g14028 ( 
.A(n_13392),
.B(n_7827),
.Y(n_14028)
);

AND2x2_ASAP7_75t_L g14029 ( 
.A(n_13362),
.B(n_7827),
.Y(n_14029)
);

BUFx6f_ASAP7_75t_L g14030 ( 
.A(n_12659),
.Y(n_14030)
);

HB1xp67_ASAP7_75t_L g14031 ( 
.A(n_13280),
.Y(n_14031)
);

INVx1_ASAP7_75t_L g14032 ( 
.A(n_12881),
.Y(n_14032)
);

OAI22xp5_ASAP7_75t_L g14033 ( 
.A1(n_13336),
.A2(n_7749),
.B1(n_7823),
.B2(n_7792),
.Y(n_14033)
);

AND2x2_ASAP7_75t_L g14034 ( 
.A(n_13367),
.B(n_7830),
.Y(n_14034)
);

INVx2_ASAP7_75t_L g14035 ( 
.A(n_12696),
.Y(n_14035)
);

NAND2xp5_ASAP7_75t_L g14036 ( 
.A(n_13361),
.B(n_9787),
.Y(n_14036)
);

INVx2_ASAP7_75t_L g14037 ( 
.A(n_12701),
.Y(n_14037)
);

INVx2_ASAP7_75t_L g14038 ( 
.A(n_12704),
.Y(n_14038)
);

INVx1_ASAP7_75t_L g14039 ( 
.A(n_12882),
.Y(n_14039)
);

INVx1_ASAP7_75t_L g14040 ( 
.A(n_12890),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_12893),
.Y(n_14041)
);

OAI22xp5_ASAP7_75t_L g14042 ( 
.A1(n_13333),
.A2(n_7749),
.B1(n_7823),
.B2(n_7792),
.Y(n_14042)
);

INVx3_ASAP7_75t_L g14043 ( 
.A(n_12983),
.Y(n_14043)
);

INVx1_ASAP7_75t_L g14044 ( 
.A(n_12903),
.Y(n_14044)
);

INVx2_ASAP7_75t_L g14045 ( 
.A(n_12711),
.Y(n_14045)
);

AND2x2_ASAP7_75t_L g14046 ( 
.A(n_13368),
.B(n_7830),
.Y(n_14046)
);

OR2x2_ASAP7_75t_L g14047 ( 
.A(n_13389),
.B(n_9373),
.Y(n_14047)
);

NOR2x1_ASAP7_75t_L g14048 ( 
.A(n_13117),
.B(n_10507),
.Y(n_14048)
);

INVx2_ASAP7_75t_L g14049 ( 
.A(n_12715),
.Y(n_14049)
);

INVx1_ASAP7_75t_L g14050 ( 
.A(n_12906),
.Y(n_14050)
);

AOI22xp33_ASAP7_75t_L g14051 ( 
.A1(n_13360),
.A2(n_9303),
.B1(n_8036),
.B2(n_8037),
.Y(n_14051)
);

AND2x2_ASAP7_75t_L g14052 ( 
.A(n_12921),
.B(n_7830),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13283),
.B(n_9303),
.Y(n_14053)
);

NAND2xp5_ASAP7_75t_L g14054 ( 
.A(n_12664),
.B(n_9787),
.Y(n_14054)
);

INVx1_ASAP7_75t_L g14055 ( 
.A(n_12908),
.Y(n_14055)
);

NAND2xp5_ASAP7_75t_L g14056 ( 
.A(n_12666),
.B(n_9792),
.Y(n_14056)
);

INVx2_ASAP7_75t_L g14057 ( 
.A(n_12720),
.Y(n_14057)
);

AND2x2_ASAP7_75t_L g14058 ( 
.A(n_13415),
.B(n_9303),
.Y(n_14058)
);

AND2x2_ASAP7_75t_L g14059 ( 
.A(n_12899),
.B(n_9303),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_12914),
.Y(n_14060)
);

AND2x2_ASAP7_75t_L g14061 ( 
.A(n_13197),
.B(n_8008),
.Y(n_14061)
);

INVx1_ASAP7_75t_L g14062 ( 
.A(n_12923),
.Y(n_14062)
);

AND2x2_ASAP7_75t_L g14063 ( 
.A(n_12891),
.B(n_8008),
.Y(n_14063)
);

INVx1_ASAP7_75t_L g14064 ( 
.A(n_12938),
.Y(n_14064)
);

INVx1_ASAP7_75t_L g14065 ( 
.A(n_12942),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13000),
.B(n_8008),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13003),
.B(n_8008),
.Y(n_14067)
);

AND2x2_ASAP7_75t_L g14068 ( 
.A(n_13227),
.B(n_8008),
.Y(n_14068)
);

NOR2xp67_ASAP7_75t_L g14069 ( 
.A(n_13004),
.B(n_10513),
.Y(n_14069)
);

AOI22xp33_ASAP7_75t_SL g14070 ( 
.A1(n_13413),
.A2(n_13385),
.B1(n_13333),
.B2(n_13406),
.Y(n_14070)
);

BUFx2_ASAP7_75t_L g14071 ( 
.A(n_13278),
.Y(n_14071)
);

INVx1_ASAP7_75t_SL g14072 ( 
.A(n_13236),
.Y(n_14072)
);

OR2x2_ASAP7_75t_L g14073 ( 
.A(n_12997),
.B(n_9373),
.Y(n_14073)
);

AND2x2_ASAP7_75t_L g14074 ( 
.A(n_13019),
.B(n_8048),
.Y(n_14074)
);

BUFx2_ASAP7_75t_L g14075 ( 
.A(n_13278),
.Y(n_14075)
);

INVx3_ASAP7_75t_L g14076 ( 
.A(n_12845),
.Y(n_14076)
);

INVx1_ASAP7_75t_L g14077 ( 
.A(n_12952),
.Y(n_14077)
);

HB1xp67_ASAP7_75t_L g14078 ( 
.A(n_13275),
.Y(n_14078)
);

INVx3_ASAP7_75t_L g14079 ( 
.A(n_12757),
.Y(n_14079)
);

BUFx6f_ASAP7_75t_L g14080 ( 
.A(n_12675),
.Y(n_14080)
);

BUFx3_ASAP7_75t_L g14081 ( 
.A(n_12937),
.Y(n_14081)
);

INVx1_ASAP7_75t_L g14082 ( 
.A(n_12966),
.Y(n_14082)
);

HB1xp67_ASAP7_75t_L g14083 ( 
.A(n_13275),
.Y(n_14083)
);

AND2x2_ASAP7_75t_L g14084 ( 
.A(n_13033),
.B(n_8048),
.Y(n_14084)
);

INVx1_ASAP7_75t_L g14085 ( 
.A(n_12967),
.Y(n_14085)
);

AND2x2_ASAP7_75t_L g14086 ( 
.A(n_13062),
.B(n_8048),
.Y(n_14086)
);

OR2x2_ASAP7_75t_L g14087 ( 
.A(n_13395),
.B(n_9373),
.Y(n_14087)
);

NAND2xp5_ASAP7_75t_L g14088 ( 
.A(n_12683),
.B(n_9792),
.Y(n_14088)
);

AOI22xp33_ASAP7_75t_L g14089 ( 
.A1(n_13402),
.A2(n_8036),
.B1(n_8037),
.B2(n_8005),
.Y(n_14089)
);

AND2x2_ASAP7_75t_L g14090 ( 
.A(n_13065),
.B(n_8048),
.Y(n_14090)
);

AOI22xp33_ASAP7_75t_L g14091 ( 
.A1(n_13372),
.A2(n_8036),
.B1(n_8037),
.B2(n_8005),
.Y(n_14091)
);

AND2x2_ASAP7_75t_L g14092 ( 
.A(n_13078),
.B(n_8048),
.Y(n_14092)
);

INVxp67_ASAP7_75t_L g14093 ( 
.A(n_13366),
.Y(n_14093)
);

AND2x4_ASAP7_75t_SL g14094 ( 
.A(n_13073),
.B(n_6760),
.Y(n_14094)
);

NOR2xp67_ASAP7_75t_L g14095 ( 
.A(n_13004),
.B(n_10513),
.Y(n_14095)
);

NAND2xp5_ASAP7_75t_L g14096 ( 
.A(n_12687),
.B(n_9798),
.Y(n_14096)
);

INVx2_ASAP7_75t_L g14097 ( 
.A(n_12722),
.Y(n_14097)
);

AND2x2_ASAP7_75t_L g14098 ( 
.A(n_13080),
.B(n_13081),
.Y(n_14098)
);

AND2x2_ASAP7_75t_L g14099 ( 
.A(n_13091),
.B(n_8053),
.Y(n_14099)
);

INVx1_ASAP7_75t_L g14100 ( 
.A(n_12971),
.Y(n_14100)
);

OAI21xp33_ASAP7_75t_L g14101 ( 
.A1(n_12809),
.A2(n_7858),
.B(n_7852),
.Y(n_14101)
);

BUFx3_ASAP7_75t_L g14102 ( 
.A(n_12943),
.Y(n_14102)
);

INVx1_ASAP7_75t_L g14103 ( 
.A(n_12972),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_12974),
.Y(n_14104)
);

OR2x2_ASAP7_75t_L g14105 ( 
.A(n_13380),
.B(n_12840),
.Y(n_14105)
);

NOR2xp33_ASAP7_75t_L g14106 ( 
.A(n_13357),
.B(n_8094),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_L g14107 ( 
.A(n_12698),
.B(n_9798),
.Y(n_14107)
);

NAND2xp5_ASAP7_75t_L g14108 ( 
.A(n_12702),
.B(n_9799),
.Y(n_14108)
);

OR2x2_ASAP7_75t_L g14109 ( 
.A(n_13380),
.B(n_8094),
.Y(n_14109)
);

AND2x2_ASAP7_75t_L g14110 ( 
.A(n_13097),
.B(n_8053),
.Y(n_14110)
);

INVx2_ASAP7_75t_L g14111 ( 
.A(n_12726),
.Y(n_14111)
);

INVx2_ASAP7_75t_L g14112 ( 
.A(n_12737),
.Y(n_14112)
);

AND2x2_ASAP7_75t_L g14113 ( 
.A(n_13111),
.B(n_8053),
.Y(n_14113)
);

INVx2_ASAP7_75t_L g14114 ( 
.A(n_12708),
.Y(n_14114)
);

INVx1_ASAP7_75t_L g14115 ( 
.A(n_12979),
.Y(n_14115)
);

INVx1_ASAP7_75t_L g14116 ( 
.A(n_12984),
.Y(n_14116)
);

AND2x2_ASAP7_75t_L g14117 ( 
.A(n_13113),
.B(n_8053),
.Y(n_14117)
);

INVx1_ASAP7_75t_L g14118 ( 
.A(n_12991),
.Y(n_14118)
);

AND2x2_ASAP7_75t_L g14119 ( 
.A(n_13119),
.B(n_8053),
.Y(n_14119)
);

INVx1_ASAP7_75t_L g14120 ( 
.A(n_12819),
.Y(n_14120)
);

INVx1_ASAP7_75t_L g14121 ( 
.A(n_13089),
.Y(n_14121)
);

AOI22xp33_ASAP7_75t_L g14122 ( 
.A1(n_13372),
.A2(n_8036),
.B1(n_8037),
.B2(n_8005),
.Y(n_14122)
);

HB1xp67_ASAP7_75t_L g14123 ( 
.A(n_13005),
.Y(n_14123)
);

AND2x2_ASAP7_75t_L g14124 ( 
.A(n_13120),
.B(n_8068),
.Y(n_14124)
);

NAND2xp5_ASAP7_75t_L g14125 ( 
.A(n_12709),
.B(n_9799),
.Y(n_14125)
);

INVx1_ASAP7_75t_L g14126 ( 
.A(n_13094),
.Y(n_14126)
);

AND2x2_ASAP7_75t_L g14127 ( 
.A(n_13251),
.B(n_8068),
.Y(n_14127)
);

INVx1_ASAP7_75t_L g14128 ( 
.A(n_13102),
.Y(n_14128)
);

AND2x4_ASAP7_75t_L g14129 ( 
.A(n_12710),
.B(n_10827),
.Y(n_14129)
);

INVx1_ASAP7_75t_L g14130 ( 
.A(n_13127),
.Y(n_14130)
);

AND2x2_ASAP7_75t_L g14131 ( 
.A(n_13123),
.B(n_8068),
.Y(n_14131)
);

OR2x2_ASAP7_75t_L g14132 ( 
.A(n_13302),
.B(n_8094),
.Y(n_14132)
);

AND2x4_ASAP7_75t_L g14133 ( 
.A(n_12716),
.B(n_10827),
.Y(n_14133)
);

INVx1_ASAP7_75t_L g14134 ( 
.A(n_13139),
.Y(n_14134)
);

INVx1_ASAP7_75t_L g14135 ( 
.A(n_13141),
.Y(n_14135)
);

HB1xp67_ASAP7_75t_L g14136 ( 
.A(n_13005),
.Y(n_14136)
);

AND2x2_ASAP7_75t_L g14137 ( 
.A(n_13126),
.B(n_8068),
.Y(n_14137)
);

INVx1_ASAP7_75t_L g14138 ( 
.A(n_12818),
.Y(n_14138)
);

AND2x2_ASAP7_75t_L g14139 ( 
.A(n_13047),
.B(n_8068),
.Y(n_14139)
);

NAND2xp5_ASAP7_75t_L g14140 ( 
.A(n_12719),
.B(n_9800),
.Y(n_14140)
);

BUFx6f_ASAP7_75t_L g14141 ( 
.A(n_12950),
.Y(n_14141)
);

INVx3_ASAP7_75t_L g14142 ( 
.A(n_12951),
.Y(n_14142)
);

BUFx6f_ASAP7_75t_L g14143 ( 
.A(n_12953),
.Y(n_14143)
);

AOI22xp33_ASAP7_75t_L g14144 ( 
.A1(n_13385),
.A2(n_8037),
.B1(n_8098),
.B2(n_8005),
.Y(n_14144)
);

INVx2_ASAP7_75t_L g14145 ( 
.A(n_13122),
.Y(n_14145)
);

INVx1_ASAP7_75t_L g14146 ( 
.A(n_12805),
.Y(n_14146)
);

HB1xp67_ASAP7_75t_L g14147 ( 
.A(n_13022),
.Y(n_14147)
);

OAI22xp5_ASAP7_75t_L g14148 ( 
.A1(n_12725),
.A2(n_7749),
.B1(n_7823),
.B2(n_7792),
.Y(n_14148)
);

AND2x2_ASAP7_75t_L g14149 ( 
.A(n_13055),
.B(n_8083),
.Y(n_14149)
);

BUFx2_ASAP7_75t_L g14150 ( 
.A(n_13022),
.Y(n_14150)
);

OR2x2_ASAP7_75t_L g14151 ( 
.A(n_12877),
.B(n_8196),
.Y(n_14151)
);

HB1xp67_ASAP7_75t_L g14152 ( 
.A(n_13024),
.Y(n_14152)
);

BUFx2_ASAP7_75t_L g14153 ( 
.A(n_13024),
.Y(n_14153)
);

INVx1_ASAP7_75t_L g14154 ( 
.A(n_13011),
.Y(n_14154)
);

AOI22xp33_ASAP7_75t_L g14155 ( 
.A1(n_12832),
.A2(n_8098),
.B1(n_8005),
.B2(n_8156),
.Y(n_14155)
);

INVx1_ASAP7_75t_L g14156 ( 
.A(n_13012),
.Y(n_14156)
);

OR2x2_ASAP7_75t_L g14157 ( 
.A(n_13299),
.B(n_8196),
.Y(n_14157)
);

BUFx2_ASAP7_75t_L g14158 ( 
.A(n_13087),
.Y(n_14158)
);

AND2x2_ASAP7_75t_L g14159 ( 
.A(n_13153),
.B(n_8083),
.Y(n_14159)
);

INVx2_ASAP7_75t_L g14160 ( 
.A(n_12854),
.Y(n_14160)
);

INVx2_ASAP7_75t_L g14161 ( 
.A(n_12856),
.Y(n_14161)
);

BUFx3_ASAP7_75t_L g14162 ( 
.A(n_12956),
.Y(n_14162)
);

INVx2_ASAP7_75t_SL g14163 ( 
.A(n_12960),
.Y(n_14163)
);

AND2x2_ASAP7_75t_L g14164 ( 
.A(n_12901),
.B(n_8083),
.Y(n_14164)
);

INVx2_ASAP7_75t_L g14165 ( 
.A(n_12778),
.Y(n_14165)
);

OAI22xp33_ASAP7_75t_L g14166 ( 
.A1(n_13142),
.A2(n_8329),
.B1(n_8340),
.B2(n_8282),
.Y(n_14166)
);

INVx1_ASAP7_75t_L g14167 ( 
.A(n_13025),
.Y(n_14167)
);

INVx1_ASAP7_75t_L g14168 ( 
.A(n_12878),
.Y(n_14168)
);

INVx2_ASAP7_75t_L g14169 ( 
.A(n_13110),
.Y(n_14169)
);

AND2x2_ASAP7_75t_L g14170 ( 
.A(n_13178),
.B(n_8083),
.Y(n_14170)
);

INVx1_ASAP7_75t_L g14171 ( 
.A(n_12883),
.Y(n_14171)
);

BUFx3_ASAP7_75t_L g14172 ( 
.A(n_12962),
.Y(n_14172)
);

INVx2_ASAP7_75t_L g14173 ( 
.A(n_12970),
.Y(n_14173)
);

INVx2_ASAP7_75t_SL g14174 ( 
.A(n_12975),
.Y(n_14174)
);

INVxp67_ASAP7_75t_L g14175 ( 
.A(n_13382),
.Y(n_14175)
);

NAND2xp5_ASAP7_75t_L g14176 ( 
.A(n_13036),
.B(n_9800),
.Y(n_14176)
);

INVx1_ASAP7_75t_L g14177 ( 
.A(n_12649),
.Y(n_14177)
);

INVx2_ASAP7_75t_L g14178 ( 
.A(n_12872),
.Y(n_14178)
);

INVx2_ASAP7_75t_L g14179 ( 
.A(n_12879),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13397),
.B(n_13014),
.Y(n_14180)
);

INVx2_ASAP7_75t_L g14181 ( 
.A(n_12886),
.Y(n_14181)
);

BUFx2_ASAP7_75t_L g14182 ( 
.A(n_13087),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_13017),
.B(n_8083),
.Y(n_14183)
);

AOI22xp33_ASAP7_75t_L g14184 ( 
.A1(n_13400),
.A2(n_8098),
.B1(n_8161),
.B2(n_8156),
.Y(n_14184)
);

AND2x4_ASAP7_75t_L g14185 ( 
.A(n_13036),
.B(n_11112),
.Y(n_14185)
);

INVx1_ASAP7_75t_L g14186 ( 
.A(n_12657),
.Y(n_14186)
);

BUFx2_ASAP7_75t_L g14187 ( 
.A(n_13406),
.Y(n_14187)
);

INVx3_ASAP7_75t_L g14188 ( 
.A(n_13069),
.Y(n_14188)
);

AND2x4_ASAP7_75t_L g14189 ( 
.A(n_13082),
.B(n_11112),
.Y(n_14189)
);

AND2x2_ASAP7_75t_L g14190 ( 
.A(n_13272),
.B(n_8099),
.Y(n_14190)
);

BUFx3_ASAP7_75t_L g14191 ( 
.A(n_12993),
.Y(n_14191)
);

AND2x2_ASAP7_75t_L g14192 ( 
.A(n_13250),
.B(n_8099),
.Y(n_14192)
);

HB1xp67_ASAP7_75t_L g14193 ( 
.A(n_13130),
.Y(n_14193)
);

OR2x2_ASAP7_75t_L g14194 ( 
.A(n_12944),
.B(n_13322),
.Y(n_14194)
);

INVx1_ASAP7_75t_L g14195 ( 
.A(n_12660),
.Y(n_14195)
);

AOI22xp33_ASAP7_75t_L g14196 ( 
.A1(n_13400),
.A2(n_8098),
.B1(n_8161),
.B2(n_8156),
.Y(n_14196)
);

NAND2xp5_ASAP7_75t_L g14197 ( 
.A(n_13128),
.B(n_9806),
.Y(n_14197)
);

AND2x2_ASAP7_75t_L g14198 ( 
.A(n_13252),
.B(n_8099),
.Y(n_14198)
);

INVx1_ASAP7_75t_L g14199 ( 
.A(n_12721),
.Y(n_14199)
);

CKINVDCx6p67_ASAP7_75t_R g14200 ( 
.A(n_13422),
.Y(n_14200)
);

OR2x2_ASAP7_75t_L g14201 ( 
.A(n_12804),
.B(n_8196),
.Y(n_14201)
);

INVx2_ASAP7_75t_L g14202 ( 
.A(n_12888),
.Y(n_14202)
);

NOR3xp33_ASAP7_75t_SL g14203 ( 
.A(n_12697),
.B(n_6976),
.C(n_6970),
.Y(n_14203)
);

INVx1_ASAP7_75t_L g14204 ( 
.A(n_12728),
.Y(n_14204)
);

INVx1_ASAP7_75t_L g14205 ( 
.A(n_12731),
.Y(n_14205)
);

INVx1_ASAP7_75t_L g14206 ( 
.A(n_13104),
.Y(n_14206)
);

INVx1_ASAP7_75t_L g14207 ( 
.A(n_13104),
.Y(n_14207)
);

NAND2xp5_ASAP7_75t_L g14208 ( 
.A(n_13319),
.B(n_9806),
.Y(n_14208)
);

OR2x2_ASAP7_75t_L g14209 ( 
.A(n_12907),
.B(n_8198),
.Y(n_14209)
);

INVx3_ASAP7_75t_L g14210 ( 
.A(n_13084),
.Y(n_14210)
);

HB1xp67_ASAP7_75t_L g14211 ( 
.A(n_13204),
.Y(n_14211)
);

AND2x2_ASAP7_75t_L g14212 ( 
.A(n_13258),
.B(n_8099),
.Y(n_14212)
);

INVx2_ASAP7_75t_L g14213 ( 
.A(n_12889),
.Y(n_14213)
);

AND2x2_ASAP7_75t_L g14214 ( 
.A(n_13261),
.B(n_13262),
.Y(n_14214)
);

OR2x2_ASAP7_75t_L g14215 ( 
.A(n_13286),
.B(n_13386),
.Y(n_14215)
);

INVx1_ASAP7_75t_L g14216 ( 
.A(n_13105),
.Y(n_14216)
);

INVx1_ASAP7_75t_L g14217 ( 
.A(n_13105),
.Y(n_14217)
);

NAND2xp5_ASAP7_75t_L g14218 ( 
.A(n_13319),
.B(n_9810),
.Y(n_14218)
);

AND2x2_ASAP7_75t_L g14219 ( 
.A(n_13369),
.B(n_8099),
.Y(n_14219)
);

INVx1_ASAP7_75t_L g14220 ( 
.A(n_13106),
.Y(n_14220)
);

INVx2_ASAP7_75t_L g14221 ( 
.A(n_12892),
.Y(n_14221)
);

OAI221xp5_ASAP7_75t_L g14222 ( 
.A1(n_13495),
.A2(n_13507),
.B1(n_13586),
.B2(n_13516),
.C(n_13453),
.Y(n_14222)
);

OR2x2_ASAP7_75t_L g14223 ( 
.A(n_14072),
.B(n_13330),
.Y(n_14223)
);

HB1xp67_ASAP7_75t_L g14224 ( 
.A(n_14150),
.Y(n_14224)
);

INVx2_ASAP7_75t_L g14225 ( 
.A(n_13478),
.Y(n_14225)
);

NOR2xp33_ASAP7_75t_L g14226 ( 
.A(n_13691),
.B(n_13008),
.Y(n_14226)
);

OAI22xp5_ASAP7_75t_L g14227 ( 
.A1(n_13708),
.A2(n_12824),
.B1(n_13436),
.B2(n_13193),
.Y(n_14227)
);

INVx1_ASAP7_75t_L g14228 ( 
.A(n_13761),
.Y(n_14228)
);

AOI22xp5_ASAP7_75t_L g14229 ( 
.A1(n_13668),
.A2(n_13364),
.B1(n_12674),
.B2(n_13441),
.Y(n_14229)
);

BUFx2_ASAP7_75t_L g14230 ( 
.A(n_13562),
.Y(n_14230)
);

HB1xp67_ASAP7_75t_L g14231 ( 
.A(n_14150),
.Y(n_14231)
);

AND2x2_ASAP7_75t_L g14232 ( 
.A(n_13489),
.B(n_13196),
.Y(n_14232)
);

INVx2_ASAP7_75t_L g14233 ( 
.A(n_13478),
.Y(n_14233)
);

INVx1_ASAP7_75t_L g14234 ( 
.A(n_13761),
.Y(n_14234)
);

NOR2xp33_ASAP7_75t_L g14235 ( 
.A(n_13489),
.B(n_13348),
.Y(n_14235)
);

INVx4_ASAP7_75t_L g14236 ( 
.A(n_13483),
.Y(n_14236)
);

AND2x2_ASAP7_75t_L g14237 ( 
.A(n_13471),
.B(n_13600),
.Y(n_14237)
);

INVx2_ASAP7_75t_L g14238 ( 
.A(n_13513),
.Y(n_14238)
);

INVx5_ASAP7_75t_L g14239 ( 
.A(n_13730),
.Y(n_14239)
);

INVx1_ASAP7_75t_L g14240 ( 
.A(n_13846),
.Y(n_14240)
);

NAND2x1_ASAP7_75t_L g14241 ( 
.A(n_13544),
.B(n_13331),
.Y(n_14241)
);

AND2x2_ASAP7_75t_L g14242 ( 
.A(n_13472),
.B(n_13284),
.Y(n_14242)
);

AND2x4_ASAP7_75t_L g14243 ( 
.A(n_13455),
.B(n_13093),
.Y(n_14243)
);

OR2x2_ASAP7_75t_L g14244 ( 
.A(n_13991),
.B(n_13201),
.Y(n_14244)
);

AND2x2_ASAP7_75t_L g14245 ( 
.A(n_13537),
.B(n_13320),
.Y(n_14245)
);

OR2x2_ASAP7_75t_L g14246 ( 
.A(n_13462),
.B(n_13340),
.Y(n_14246)
);

AND2x2_ASAP7_75t_L g14247 ( 
.A(n_13568),
.B(n_13320),
.Y(n_14247)
);

AO31x2_ASAP7_75t_L g14248 ( 
.A1(n_13846),
.A2(n_13364),
.A3(n_13109),
.B(n_13114),
.Y(n_14248)
);

INVx1_ASAP7_75t_L g14249 ( 
.A(n_13852),
.Y(n_14249)
);

NOR2x1p5_ASAP7_75t_L g14250 ( 
.A(n_13800),
.B(n_13351),
.Y(n_14250)
);

INVx2_ASAP7_75t_L g14251 ( 
.A(n_13513),
.Y(n_14251)
);

INVx1_ASAP7_75t_L g14252 ( 
.A(n_13852),
.Y(n_14252)
);

INVx1_ASAP7_75t_L g14253 ( 
.A(n_13456),
.Y(n_14253)
);

OR2x2_ASAP7_75t_L g14254 ( 
.A(n_13554),
.B(n_12828),
.Y(n_14254)
);

INVx2_ASAP7_75t_L g14255 ( 
.A(n_14153),
.Y(n_14255)
);

AND2x2_ASAP7_75t_L g14256 ( 
.A(n_13579),
.B(n_13327),
.Y(n_14256)
);

AND2x2_ASAP7_75t_L g14257 ( 
.A(n_13710),
.B(n_13910),
.Y(n_14257)
);

BUFx2_ASAP7_75t_L g14258 ( 
.A(n_13562),
.Y(n_14258)
);

INVx1_ASAP7_75t_L g14259 ( 
.A(n_13576),
.Y(n_14259)
);

NOR2x1_ASAP7_75t_L g14260 ( 
.A(n_14071),
.B(n_12751),
.Y(n_14260)
);

INVx1_ASAP7_75t_L g14261 ( 
.A(n_13527),
.Y(n_14261)
);

NAND4xp25_ASAP7_75t_L g14262 ( 
.A(n_14070),
.B(n_12588),
.C(n_13430),
.D(n_13434),
.Y(n_14262)
);

HB1xp67_ASAP7_75t_L g14263 ( 
.A(n_14153),
.Y(n_14263)
);

INVx2_ASAP7_75t_L g14264 ( 
.A(n_14158),
.Y(n_14264)
);

INVx2_ASAP7_75t_L g14265 ( 
.A(n_14158),
.Y(n_14265)
);

BUFx2_ASAP7_75t_L g14266 ( 
.A(n_14071),
.Y(n_14266)
);

INVx1_ASAP7_75t_L g14267 ( 
.A(n_13542),
.Y(n_14267)
);

INVx1_ASAP7_75t_L g14268 ( 
.A(n_13830),
.Y(n_14268)
);

AND2x4_ASAP7_75t_SL g14269 ( 
.A(n_13793),
.B(n_13099),
.Y(n_14269)
);

AOI22xp5_ASAP7_75t_L g14270 ( 
.A1(n_13864),
.A2(n_13408),
.B1(n_13425),
.B2(n_13407),
.Y(n_14270)
);

AND2x2_ASAP7_75t_L g14271 ( 
.A(n_13479),
.B(n_13327),
.Y(n_14271)
);

INVx1_ASAP7_75t_L g14272 ( 
.A(n_13878),
.Y(n_14272)
);

INVx2_ASAP7_75t_L g14273 ( 
.A(n_14182),
.Y(n_14273)
);

BUFx6f_ASAP7_75t_L g14274 ( 
.A(n_13693),
.Y(n_14274)
);

BUFx2_ASAP7_75t_L g14275 ( 
.A(n_14075),
.Y(n_14275)
);

AND2x2_ASAP7_75t_L g14276 ( 
.A(n_13539),
.B(n_13285),
.Y(n_14276)
);

NAND2xp5_ASAP7_75t_SL g14277 ( 
.A(n_13641),
.B(n_13331),
.Y(n_14277)
);

NAND2xp5_ASAP7_75t_L g14278 ( 
.A(n_13445),
.B(n_13437),
.Y(n_14278)
);

AOI22xp33_ASAP7_75t_SL g14279 ( 
.A1(n_13630),
.A2(n_13406),
.B1(n_13311),
.B2(n_13306),
.Y(n_14279)
);

INVx1_ASAP7_75t_L g14280 ( 
.A(n_13881),
.Y(n_14280)
);

INVx2_ASAP7_75t_L g14281 ( 
.A(n_14182),
.Y(n_14281)
);

AND2x2_ASAP7_75t_L g14282 ( 
.A(n_13726),
.B(n_13288),
.Y(n_14282)
);

INVx1_ASAP7_75t_L g14283 ( 
.A(n_13903),
.Y(n_14283)
);

OR2x2_ASAP7_75t_L g14284 ( 
.A(n_14012),
.B(n_12887),
.Y(n_14284)
);

AND2x2_ASAP7_75t_L g14285 ( 
.A(n_13684),
.B(n_13291),
.Y(n_14285)
);

BUFx3_ASAP7_75t_L g14286 ( 
.A(n_13502),
.Y(n_14286)
);

OR2x2_ASAP7_75t_L g14287 ( 
.A(n_13820),
.B(n_12909),
.Y(n_14287)
);

HB1xp67_ASAP7_75t_L g14288 ( 
.A(n_14123),
.Y(n_14288)
);

NOR2x1_ASAP7_75t_L g14289 ( 
.A(n_14075),
.B(n_13877),
.Y(n_14289)
);

AND2x2_ASAP7_75t_L g14290 ( 
.A(n_13660),
.B(n_13300),
.Y(n_14290)
);

INVx1_ASAP7_75t_L g14291 ( 
.A(n_14136),
.Y(n_14291)
);

AO21x2_ASAP7_75t_L g14292 ( 
.A1(n_13959),
.A2(n_13190),
.B(n_13167),
.Y(n_14292)
);

INVx3_ASAP7_75t_L g14293 ( 
.A(n_13544),
.Y(n_14293)
);

AND2x2_ASAP7_75t_L g14294 ( 
.A(n_13474),
.B(n_13307),
.Y(n_14294)
);

OR2x2_ASAP7_75t_L g14295 ( 
.A(n_13971),
.B(n_12919),
.Y(n_14295)
);

INVx2_ASAP7_75t_L g14296 ( 
.A(n_13809),
.Y(n_14296)
);

INVx2_ASAP7_75t_L g14297 ( 
.A(n_13545),
.Y(n_14297)
);

INVx2_ASAP7_75t_L g14298 ( 
.A(n_13582),
.Y(n_14298)
);

INVx1_ASAP7_75t_L g14299 ( 
.A(n_14147),
.Y(n_14299)
);

AND2x2_ASAP7_75t_L g14300 ( 
.A(n_13514),
.B(n_13629),
.Y(n_14300)
);

HB1xp67_ASAP7_75t_L g14301 ( 
.A(n_14152),
.Y(n_14301)
);

AND2x2_ASAP7_75t_L g14302 ( 
.A(n_13650),
.B(n_13314),
.Y(n_14302)
);

OR2x2_ASAP7_75t_L g14303 ( 
.A(n_13448),
.B(n_12945),
.Y(n_14303)
);

INVx1_ASAP7_75t_L g14304 ( 
.A(n_13512),
.Y(n_14304)
);

OR2x2_ASAP7_75t_L g14305 ( 
.A(n_13899),
.B(n_14078),
.Y(n_14305)
);

AND2x2_ASAP7_75t_L g14306 ( 
.A(n_13653),
.B(n_13281),
.Y(n_14306)
);

HB1xp67_ASAP7_75t_L g14307 ( 
.A(n_13734),
.Y(n_14307)
);

INVx1_ASAP7_75t_SL g14308 ( 
.A(n_13636),
.Y(n_14308)
);

BUFx2_ASAP7_75t_L g14309 ( 
.A(n_13636),
.Y(n_14309)
);

INVx1_ASAP7_75t_SL g14310 ( 
.A(n_13640),
.Y(n_14310)
);

INVx2_ASAP7_75t_L g14311 ( 
.A(n_13655),
.Y(n_14311)
);

AND2x2_ASAP7_75t_L g14312 ( 
.A(n_13656),
.B(n_13417),
.Y(n_14312)
);

INVx2_ASAP7_75t_L g14313 ( 
.A(n_13707),
.Y(n_14313)
);

INVx1_ASAP7_75t_L g14314 ( 
.A(n_13558),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_13590),
.Y(n_14315)
);

OR2x2_ASAP7_75t_L g14316 ( 
.A(n_14083),
.B(n_13996),
.Y(n_14316)
);

AOI21xp33_ASAP7_75t_L g14317 ( 
.A1(n_13461),
.A2(n_13408),
.B(n_13407),
.Y(n_14317)
);

BUFx2_ASAP7_75t_L g14318 ( 
.A(n_13640),
.Y(n_14318)
);

INVx2_ASAP7_75t_L g14319 ( 
.A(n_14076),
.Y(n_14319)
);

AOI22xp33_ASAP7_75t_L g14320 ( 
.A1(n_13574),
.A2(n_13394),
.B1(n_13431),
.B2(n_13433),
.Y(n_14320)
);

INVxp67_ASAP7_75t_L g14321 ( 
.A(n_13553),
.Y(n_14321)
);

AND2x2_ASAP7_75t_L g14322 ( 
.A(n_13855),
.B(n_13419),
.Y(n_14322)
);

INVxp67_ASAP7_75t_L g14323 ( 
.A(n_13695),
.Y(n_14323)
);

INVx1_ASAP7_75t_L g14324 ( 
.A(n_14211),
.Y(n_14324)
);

INVx2_ASAP7_75t_L g14325 ( 
.A(n_13747),
.Y(n_14325)
);

AND2x4_ASAP7_75t_L g14326 ( 
.A(n_13454),
.B(n_13135),
.Y(n_14326)
);

AND2x2_ASAP7_75t_L g14327 ( 
.A(n_13588),
.B(n_13424),
.Y(n_14327)
);

BUFx6f_ASAP7_75t_L g14328 ( 
.A(n_13693),
.Y(n_14328)
);

BUFx3_ASAP7_75t_L g14329 ( 
.A(n_13818),
.Y(n_14329)
);

NAND2xp5_ASAP7_75t_L g14330 ( 
.A(n_13695),
.B(n_13112),
.Y(n_14330)
);

INVx2_ASAP7_75t_SL g14331 ( 
.A(n_13497),
.Y(n_14331)
);

NAND2xp5_ASAP7_75t_L g14332 ( 
.A(n_13926),
.B(n_13112),
.Y(n_14332)
);

AO21x2_ASAP7_75t_L g14333 ( 
.A1(n_13968),
.A2(n_13109),
.B(n_13106),
.Y(n_14333)
);

AND2x2_ASAP7_75t_L g14334 ( 
.A(n_13596),
.B(n_13334),
.Y(n_14334)
);

NAND2xp5_ASAP7_75t_L g14335 ( 
.A(n_13926),
.B(n_13135),
.Y(n_14335)
);

INVx1_ASAP7_75t_L g14336 ( 
.A(n_13624),
.Y(n_14336)
);

INVx2_ASAP7_75t_SL g14337 ( 
.A(n_13538),
.Y(n_14337)
);

INVx2_ASAP7_75t_L g14338 ( 
.A(n_13768),
.Y(n_14338)
);

INVx3_ASAP7_75t_L g14339 ( 
.A(n_13518),
.Y(n_14339)
);

HB1xp67_ASAP7_75t_L g14340 ( 
.A(n_13802),
.Y(n_14340)
);

BUFx3_ASAP7_75t_L g14341 ( 
.A(n_13860),
.Y(n_14341)
);

INVx2_ASAP7_75t_L g14342 ( 
.A(n_13797),
.Y(n_14342)
);

INVxp67_ASAP7_75t_SL g14343 ( 
.A(n_13645),
.Y(n_14343)
);

INVx1_ASAP7_75t_L g14344 ( 
.A(n_13773),
.Y(n_14344)
);

INVx1_ASAP7_75t_L g14345 ( 
.A(n_13785),
.Y(n_14345)
);

NAND2xp5_ASAP7_75t_L g14346 ( 
.A(n_13677),
.B(n_13027),
.Y(n_14346)
);

INVx1_ASAP7_75t_L g14347 ( 
.A(n_13904),
.Y(n_14347)
);

AND2x2_ASAP7_75t_L g14348 ( 
.A(n_13535),
.B(n_13349),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_13985),
.Y(n_14349)
);

HB1xp67_ASAP7_75t_L g14350 ( 
.A(n_13790),
.Y(n_14350)
);

BUFx3_ASAP7_75t_L g14351 ( 
.A(n_13676),
.Y(n_14351)
);

BUFx2_ASAP7_75t_L g14352 ( 
.A(n_13532),
.Y(n_14352)
);

INVx5_ASAP7_75t_L g14353 ( 
.A(n_13602),
.Y(n_14353)
);

AND2x2_ASAP7_75t_L g14354 ( 
.A(n_13561),
.B(n_13352),
.Y(n_14354)
);

HB1xp67_ASAP7_75t_L g14355 ( 
.A(n_13804),
.Y(n_14355)
);

INVx2_ASAP7_75t_L g14356 ( 
.A(n_13805),
.Y(n_14356)
);

INVx2_ASAP7_75t_L g14357 ( 
.A(n_13825),
.Y(n_14357)
);

BUFx2_ASAP7_75t_L g14358 ( 
.A(n_13470),
.Y(n_14358)
);

AND2x4_ASAP7_75t_L g14359 ( 
.A(n_13972),
.B(n_12981),
.Y(n_14359)
);

AND2x4_ASAP7_75t_L g14360 ( 
.A(n_14043),
.B(n_12982),
.Y(n_14360)
);

OAI22xp5_ASAP7_75t_L g14361 ( 
.A1(n_13557),
.A2(n_13321),
.B1(n_13426),
.B2(n_13425),
.Y(n_14361)
);

NAND2xp5_ASAP7_75t_L g14362 ( 
.A(n_13897),
.B(n_13034),
.Y(n_14362)
);

INVx2_ASAP7_75t_L g14363 ( 
.A(n_13970),
.Y(n_14363)
);

OA21x2_ASAP7_75t_L g14364 ( 
.A1(n_13877),
.A2(n_13212),
.B(n_13198),
.Y(n_14364)
);

AND2x2_ASAP7_75t_L g14365 ( 
.A(n_13778),
.B(n_13289),
.Y(n_14365)
);

OAI21xp5_ASAP7_75t_SL g14366 ( 
.A1(n_13547),
.A2(n_13216),
.B(n_13426),
.Y(n_14366)
);

BUFx2_ASAP7_75t_L g14367 ( 
.A(n_13896),
.Y(n_14367)
);

BUFx2_ASAP7_75t_L g14368 ( 
.A(n_13896),
.Y(n_14368)
);

BUFx6f_ASAP7_75t_L g14369 ( 
.A(n_13604),
.Y(n_14369)
);

INVx3_ASAP7_75t_L g14370 ( 
.A(n_13518),
.Y(n_14370)
);

AND2x2_ASAP7_75t_L g14371 ( 
.A(n_13634),
.B(n_13449),
.Y(n_14371)
);

AND2x4_ASAP7_75t_L g14372 ( 
.A(n_13491),
.B(n_12986),
.Y(n_14372)
);

INVx2_ASAP7_75t_L g14373 ( 
.A(n_13998),
.Y(n_14373)
);

AND2x2_ASAP7_75t_L g14374 ( 
.A(n_13550),
.B(n_13248),
.Y(n_14374)
);

AND2x2_ASAP7_75t_L g14375 ( 
.A(n_13567),
.B(n_13463),
.Y(n_14375)
);

INVx2_ASAP7_75t_SL g14376 ( 
.A(n_14141),
.Y(n_14376)
);

INVx1_ASAP7_75t_L g14377 ( 
.A(n_14206),
.Y(n_14377)
);

INVxp67_ASAP7_75t_L g14378 ( 
.A(n_13827),
.Y(n_14378)
);

AND2x2_ASAP7_75t_L g14379 ( 
.A(n_13680),
.B(n_13387),
.Y(n_14379)
);

BUFx6f_ASAP7_75t_L g14380 ( 
.A(n_13861),
.Y(n_14380)
);

AND2x2_ASAP7_75t_L g14381 ( 
.A(n_13446),
.B(n_13387),
.Y(n_14381)
);

INVx2_ASAP7_75t_L g14382 ( 
.A(n_14141),
.Y(n_14382)
);

INVx2_ASAP7_75t_L g14383 ( 
.A(n_14141),
.Y(n_14383)
);

INVx2_ASAP7_75t_L g14384 ( 
.A(n_13451),
.Y(n_14384)
);

INVx1_ASAP7_75t_L g14385 ( 
.A(n_14207),
.Y(n_14385)
);

NAND2xp5_ASAP7_75t_L g14386 ( 
.A(n_13505),
.B(n_13037),
.Y(n_14386)
);

OR2x6_ASAP7_75t_L g14387 ( 
.A(n_13599),
.B(n_13001),
.Y(n_14387)
);

AND2x2_ASAP7_75t_L g14388 ( 
.A(n_13667),
.B(n_13202),
.Y(n_14388)
);

HB1xp67_ASAP7_75t_L g14389 ( 
.A(n_13821),
.Y(n_14389)
);

BUFx3_ASAP7_75t_L g14390 ( 
.A(n_13676),
.Y(n_14390)
);

INVx1_ASAP7_75t_L g14391 ( 
.A(n_14216),
.Y(n_14391)
);

HB1xp67_ASAP7_75t_L g14392 ( 
.A(n_14187),
.Y(n_14392)
);

NAND2xp5_ASAP7_75t_L g14393 ( 
.A(n_13944),
.B(n_13044),
.Y(n_14393)
);

OR2x2_ASAP7_75t_L g14394 ( 
.A(n_14031),
.B(n_12957),
.Y(n_14394)
);

INVx2_ASAP7_75t_L g14395 ( 
.A(n_13451),
.Y(n_14395)
);

OR2x2_ASAP7_75t_L g14396 ( 
.A(n_13964),
.B(n_12992),
.Y(n_14396)
);

AND2x2_ASAP7_75t_L g14397 ( 
.A(n_13499),
.B(n_13203),
.Y(n_14397)
);

AO21x2_ASAP7_75t_L g14398 ( 
.A1(n_13564),
.A2(n_13118),
.B(n_13114),
.Y(n_14398)
);

INVxp67_ASAP7_75t_L g14399 ( 
.A(n_13757),
.Y(n_14399)
);

AND2x2_ASAP7_75t_L g14400 ( 
.A(n_13812),
.B(n_13218),
.Y(n_14400)
);

INVx2_ASAP7_75t_L g14401 ( 
.A(n_13460),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_14217),
.Y(n_14402)
);

HB1xp67_ASAP7_75t_L g14403 ( 
.A(n_14187),
.Y(n_14403)
);

INVx2_ASAP7_75t_L g14404 ( 
.A(n_13460),
.Y(n_14404)
);

OAI211xp5_ASAP7_75t_L g14405 ( 
.A1(n_13493),
.A2(n_13435),
.B(n_13145),
.C(n_13393),
.Y(n_14405)
);

NOR2x1_ASAP7_75t_SL g14406 ( 
.A(n_13662),
.B(n_13209),
.Y(n_14406)
);

OAI31xp33_ASAP7_75t_L g14407 ( 
.A1(n_13523),
.A2(n_13435),
.A3(n_12754),
.B(n_13393),
.Y(n_14407)
);

INVx2_ASAP7_75t_L g14408 ( 
.A(n_13526),
.Y(n_14408)
);

INVx2_ASAP7_75t_L g14409 ( 
.A(n_13533),
.Y(n_14409)
);

NAND2xp5_ASAP7_75t_L g14410 ( 
.A(n_13952),
.B(n_13046),
.Y(n_14410)
);

INVx2_ASAP7_75t_L g14411 ( 
.A(n_13819),
.Y(n_14411)
);

AOI22xp5_ASAP7_75t_L g14412 ( 
.A1(n_13628),
.A2(n_13386),
.B1(n_13398),
.B2(n_13341),
.Y(n_14412)
);

AND2x2_ASAP7_75t_L g14413 ( 
.A(n_13601),
.B(n_13383),
.Y(n_14413)
);

INVx1_ASAP7_75t_L g14414 ( 
.A(n_14220),
.Y(n_14414)
);

NAND2xp5_ASAP7_75t_L g14415 ( 
.A(n_13501),
.B(n_13052),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_13443),
.Y(n_14416)
);

AND2x2_ASAP7_75t_L g14417 ( 
.A(n_13608),
.B(n_13232),
.Y(n_14417)
);

AND2x2_ASAP7_75t_L g14418 ( 
.A(n_13694),
.B(n_13234),
.Y(n_14418)
);

AND2x2_ASAP7_75t_L g14419 ( 
.A(n_13698),
.B(n_13347),
.Y(n_14419)
);

OR2x2_ASAP7_75t_L g14420 ( 
.A(n_13457),
.B(n_13013),
.Y(n_14420)
);

INVx2_ASAP7_75t_L g14421 ( 
.A(n_13617),
.Y(n_14421)
);

HB1xp67_ASAP7_75t_L g14422 ( 
.A(n_13757),
.Y(n_14422)
);

AND2x2_ASAP7_75t_L g14423 ( 
.A(n_13701),
.B(n_13350),
.Y(n_14423)
);

AOI22xp33_ASAP7_75t_L g14424 ( 
.A1(n_13465),
.A2(n_13398),
.B1(n_13376),
.B2(n_13374),
.Y(n_14424)
);

NAND2x1_ASAP7_75t_L g14425 ( 
.A(n_13999),
.B(n_13124),
.Y(n_14425)
);

INVx3_ASAP7_75t_L g14426 ( 
.A(n_13609),
.Y(n_14426)
);

INVx1_ASAP7_75t_L g14427 ( 
.A(n_13444),
.Y(n_14427)
);

INVx2_ASAP7_75t_SL g14428 ( 
.A(n_13584),
.Y(n_14428)
);

INVxp67_ASAP7_75t_SL g14429 ( 
.A(n_13988),
.Y(n_14429)
);

INVx3_ASAP7_75t_L g14430 ( 
.A(n_14143),
.Y(n_14430)
);

INVxp67_ASAP7_75t_SL g14431 ( 
.A(n_13799),
.Y(n_14431)
);

INVx1_ASAP7_75t_L g14432 ( 
.A(n_13447),
.Y(n_14432)
);

INVx4_ASAP7_75t_L g14433 ( 
.A(n_13496),
.Y(n_14433)
);

INVx1_ASAP7_75t_L g14434 ( 
.A(n_14154),
.Y(n_14434)
);

CKINVDCx6p67_ASAP7_75t_R g14435 ( 
.A(n_13829),
.Y(n_14435)
);

INVx1_ASAP7_75t_L g14436 ( 
.A(n_14156),
.Y(n_14436)
);

HB1xp67_ASAP7_75t_L g14437 ( 
.A(n_14193),
.Y(n_14437)
);

NOR2x1_ASAP7_75t_L g14438 ( 
.A(n_14004),
.B(n_12571),
.Y(n_14438)
);

INVx1_ASAP7_75t_L g14439 ( 
.A(n_14167),
.Y(n_14439)
);

INVx1_ASAP7_75t_L g14440 ( 
.A(n_13464),
.Y(n_14440)
);

INVx1_ASAP7_75t_L g14441 ( 
.A(n_13466),
.Y(n_14441)
);

AND2x4_ASAP7_75t_L g14442 ( 
.A(n_13543),
.B(n_12995),
.Y(n_14442)
);

INVx3_ASAP7_75t_L g14443 ( 
.A(n_14143),
.Y(n_14443)
);

INVx1_ASAP7_75t_L g14444 ( 
.A(n_13468),
.Y(n_14444)
);

AO21x2_ASAP7_75t_L g14445 ( 
.A1(n_13521),
.A2(n_13121),
.B(n_13118),
.Y(n_14445)
);

NAND2xp5_ASAP7_75t_L g14446 ( 
.A(n_13832),
.B(n_13054),
.Y(n_14446)
);

CKINVDCx16_ASAP7_75t_R g14447 ( 
.A(n_13610),
.Y(n_14447)
);

AND2x4_ASAP7_75t_L g14448 ( 
.A(n_13560),
.B(n_12996),
.Y(n_14448)
);

AOI221xp5_ASAP7_75t_L g14449 ( 
.A1(n_13801),
.A2(n_13341),
.B1(n_12563),
.B2(n_13057),
.C(n_12618),
.Y(n_14449)
);

INVx1_ASAP7_75t_L g14450 ( 
.A(n_13473),
.Y(n_14450)
);

AND2x2_ASAP7_75t_L g14451 ( 
.A(n_13504),
.B(n_13355),
.Y(n_14451)
);

OR2x2_ASAP7_75t_L g14452 ( 
.A(n_13593),
.B(n_12999),
.Y(n_14452)
);

INVx1_ASAP7_75t_L g14453 ( 
.A(n_13476),
.Y(n_14453)
);

OAI31xp33_ASAP7_75t_L g14454 ( 
.A1(n_13791),
.A2(n_13401),
.A3(n_13371),
.B(n_13370),
.Y(n_14454)
);

INVx1_ASAP7_75t_L g14455 ( 
.A(n_13477),
.Y(n_14455)
);

AND2x2_ASAP7_75t_L g14456 ( 
.A(n_13498),
.B(n_13186),
.Y(n_14456)
);

INVx2_ASAP7_75t_L g14457 ( 
.A(n_13748),
.Y(n_14457)
);

AND2x2_ASAP7_75t_L g14458 ( 
.A(n_13888),
.B(n_13194),
.Y(n_14458)
);

HB1xp67_ASAP7_75t_L g14459 ( 
.A(n_14069),
.Y(n_14459)
);

INVx1_ASAP7_75t_L g14460 ( 
.A(n_13480),
.Y(n_14460)
);

INVx1_ASAP7_75t_L g14461 ( 
.A(n_13481),
.Y(n_14461)
);

AND2x2_ASAP7_75t_L g14462 ( 
.A(n_13647),
.B(n_12940),
.Y(n_14462)
);

INVx2_ASAP7_75t_L g14463 ( 
.A(n_13750),
.Y(n_14463)
);

OR2x2_ASAP7_75t_L g14464 ( 
.A(n_13743),
.B(n_13006),
.Y(n_14464)
);

AOI221xp5_ASAP7_75t_L g14465 ( 
.A1(n_13876),
.A2(n_13292),
.B1(n_13010),
.B2(n_13020),
.C(n_13016),
.Y(n_14465)
);

INVx1_ASAP7_75t_L g14466 ( 
.A(n_13482),
.Y(n_14466)
);

AND2x2_ASAP7_75t_L g14467 ( 
.A(n_13719),
.B(n_12955),
.Y(n_14467)
);

INVx3_ASAP7_75t_L g14468 ( 
.A(n_14081),
.Y(n_14468)
);

INVx3_ASAP7_75t_L g14469 ( 
.A(n_14102),
.Y(n_14469)
);

NAND2xp5_ASAP7_75t_L g14470 ( 
.A(n_13729),
.B(n_13007),
.Y(n_14470)
);

NOR2x1_ASAP7_75t_L g14471 ( 
.A(n_14004),
.B(n_13075),
.Y(n_14471)
);

AND2x2_ASAP7_75t_L g14472 ( 
.A(n_13733),
.B(n_12961),
.Y(n_14472)
);

HB1xp67_ASAP7_75t_L g14473 ( 
.A(n_14095),
.Y(n_14473)
);

CKINVDCx16_ASAP7_75t_R g14474 ( 
.A(n_14017),
.Y(n_14474)
);

OAI211xp5_ASAP7_75t_L g14475 ( 
.A1(n_13681),
.A2(n_13138),
.B(n_13206),
.C(n_13028),
.Y(n_14475)
);

AND2x2_ASAP7_75t_L g14476 ( 
.A(n_13737),
.B(n_12963),
.Y(n_14476)
);

INVx1_ASAP7_75t_L g14477 ( 
.A(n_13485),
.Y(n_14477)
);

INVx1_ASAP7_75t_L g14478 ( 
.A(n_13486),
.Y(n_14478)
);

INVx2_ASAP7_75t_L g14479 ( 
.A(n_13769),
.Y(n_14479)
);

INVx1_ASAP7_75t_L g14480 ( 
.A(n_13490),
.Y(n_14480)
);

INVx2_ASAP7_75t_L g14481 ( 
.A(n_13861),
.Y(n_14481)
);

HB1xp67_ASAP7_75t_L g14482 ( 
.A(n_14162),
.Y(n_14482)
);

INVx1_ASAP7_75t_L g14483 ( 
.A(n_13492),
.Y(n_14483)
);

INVx1_ASAP7_75t_L g14484 ( 
.A(n_13500),
.Y(n_14484)
);

INVx2_ASAP7_75t_L g14485 ( 
.A(n_13977),
.Y(n_14485)
);

HB1xp67_ASAP7_75t_L g14486 ( 
.A(n_14172),
.Y(n_14486)
);

NAND2xp5_ASAP7_75t_L g14487 ( 
.A(n_13909),
.B(n_13045),
.Y(n_14487)
);

AND2x2_ASAP7_75t_L g14488 ( 
.A(n_13975),
.B(n_12964),
.Y(n_14488)
);

BUFx3_ASAP7_75t_L g14489 ( 
.A(n_13977),
.Y(n_14489)
);

AND2x2_ASAP7_75t_L g14490 ( 
.A(n_13674),
.B(n_12965),
.Y(n_14490)
);

INVx1_ASAP7_75t_L g14491 ( 
.A(n_13509),
.Y(n_14491)
);

INVx2_ASAP7_75t_L g14492 ( 
.A(n_14030),
.Y(n_14492)
);

NOR2xp33_ASAP7_75t_L g14493 ( 
.A(n_13475),
.B(n_12928),
.Y(n_14493)
);

INVx4_ASAP7_75t_L g14494 ( 
.A(n_14030),
.Y(n_14494)
);

HB1xp67_ASAP7_75t_L g14495 ( 
.A(n_14003),
.Y(n_14495)
);

AND2x2_ASAP7_75t_L g14496 ( 
.A(n_13563),
.B(n_12930),
.Y(n_14496)
);

OR2x2_ASAP7_75t_L g14497 ( 
.A(n_14093),
.B(n_13048),
.Y(n_14497)
);

AOI21xp5_ASAP7_75t_SL g14498 ( 
.A1(n_13487),
.A2(n_13276),
.B(n_13158),
.Y(n_14498)
);

INVx2_ASAP7_75t_L g14499 ( 
.A(n_14080),
.Y(n_14499)
);

NAND2x1p5_ASAP7_75t_L g14500 ( 
.A(n_13978),
.B(n_13051),
.Y(n_14500)
);

NAND2xp5_ASAP7_75t_L g14501 ( 
.A(n_13847),
.B(n_13061),
.Y(n_14501)
);

NAND2xp5_ASAP7_75t_L g14502 ( 
.A(n_13936),
.B(n_13067),
.Y(n_14502)
);

INVx2_ASAP7_75t_L g14503 ( 
.A(n_14080),
.Y(n_14503)
);

AND2x2_ASAP7_75t_L g14504 ( 
.A(n_14200),
.B(n_12933),
.Y(n_14504)
);

INVx2_ASAP7_75t_L g14505 ( 
.A(n_13828),
.Y(n_14505)
);

AO21x2_ASAP7_75t_L g14506 ( 
.A1(n_13506),
.A2(n_13131),
.B(n_13121),
.Y(n_14506)
);

INVx1_ASAP7_75t_L g14507 ( 
.A(n_13511),
.Y(n_14507)
);

AND2x2_ASAP7_75t_L g14508 ( 
.A(n_13786),
.B(n_12990),
.Y(n_14508)
);

NAND2xp5_ASAP7_75t_L g14509 ( 
.A(n_13936),
.B(n_14175),
.Y(n_14509)
);

INVx1_ASAP7_75t_L g14510 ( 
.A(n_13515),
.Y(n_14510)
);

AND2x2_ASAP7_75t_L g14511 ( 
.A(n_13746),
.B(n_13156),
.Y(n_14511)
);

NOR2xp33_ASAP7_75t_L g14512 ( 
.A(n_13503),
.B(n_13418),
.Y(n_14512)
);

HB1xp67_ASAP7_75t_L g14513 ( 
.A(n_13669),
.Y(n_14513)
);

INVx1_ASAP7_75t_SL g14514 ( 
.A(n_13943),
.Y(n_14514)
);

AND2x4_ASAP7_75t_L g14515 ( 
.A(n_13678),
.B(n_13399),
.Y(n_14515)
);

INVx2_ASAP7_75t_L g14516 ( 
.A(n_13844),
.Y(n_14516)
);

AND2x2_ASAP7_75t_L g14517 ( 
.A(n_13555),
.B(n_13160),
.Y(n_14517)
);

AND2x2_ASAP7_75t_L g14518 ( 
.A(n_13638),
.B(n_13164),
.Y(n_14518)
);

INVx1_ASAP7_75t_L g14519 ( 
.A(n_13519),
.Y(n_14519)
);

INVx3_ASAP7_75t_L g14520 ( 
.A(n_13584),
.Y(n_14520)
);

INVx2_ASAP7_75t_L g14521 ( 
.A(n_13863),
.Y(n_14521)
);

AND2x2_ASAP7_75t_L g14522 ( 
.A(n_13643),
.B(n_13467),
.Y(n_14522)
);

INVx1_ASAP7_75t_L g14523 ( 
.A(n_13520),
.Y(n_14523)
);

INVx1_ASAP7_75t_L g14524 ( 
.A(n_13522),
.Y(n_14524)
);

AND2x4_ASAP7_75t_L g14525 ( 
.A(n_13954),
.B(n_13384),
.Y(n_14525)
);

NAND2xp5_ASAP7_75t_L g14526 ( 
.A(n_14142),
.B(n_14163),
.Y(n_14526)
);

HB1xp67_ASAP7_75t_L g14527 ( 
.A(n_13569),
.Y(n_14527)
);

INVx2_ASAP7_75t_L g14528 ( 
.A(n_13866),
.Y(n_14528)
);

INVx3_ASAP7_75t_L g14529 ( 
.A(n_13720),
.Y(n_14529)
);

HB1xp67_ASAP7_75t_L g14530 ( 
.A(n_13581),
.Y(n_14530)
);

AND2x4_ASAP7_75t_L g14531 ( 
.A(n_13956),
.B(n_13396),
.Y(n_14531)
);

INVx1_ASAP7_75t_L g14532 ( 
.A(n_13524),
.Y(n_14532)
);

INVx1_ASAP7_75t_SL g14533 ( 
.A(n_13851),
.Y(n_14533)
);

OR2x2_ASAP7_75t_L g14534 ( 
.A(n_13450),
.B(n_12654),
.Y(n_14534)
);

AND2x2_ASAP7_75t_L g14535 ( 
.A(n_13459),
.B(n_13429),
.Y(n_14535)
);

INVx1_ASAP7_75t_L g14536 ( 
.A(n_13528),
.Y(n_14536)
);

BUFx2_ASAP7_75t_L g14537 ( 
.A(n_13874),
.Y(n_14537)
);

INVx1_ASAP7_75t_L g14538 ( 
.A(n_13529),
.Y(n_14538)
);

AND2x2_ASAP7_75t_L g14539 ( 
.A(n_14061),
.B(n_13432),
.Y(n_14539)
);

NOR2xp33_ASAP7_75t_L g14540 ( 
.A(n_13664),
.B(n_13337),
.Y(n_14540)
);

AND2x4_ASAP7_75t_L g14541 ( 
.A(n_13587),
.B(n_13155),
.Y(n_14541)
);

AND2x2_ASAP7_75t_L g14542 ( 
.A(n_13709),
.B(n_13713),
.Y(n_14542)
);

OR2x2_ASAP7_75t_L g14543 ( 
.A(n_14157),
.B(n_12690),
.Y(n_14543)
);

AND2x2_ASAP7_75t_L g14544 ( 
.A(n_13714),
.B(n_13338),
.Y(n_14544)
);

AND2x2_ASAP7_75t_L g14545 ( 
.A(n_13442),
.B(n_13342),
.Y(n_14545)
);

INVx3_ASAP7_75t_L g14546 ( 
.A(n_13720),
.Y(n_14546)
);

INVx2_ASAP7_75t_L g14547 ( 
.A(n_13880),
.Y(n_14547)
);

NAND2xp5_ASAP7_75t_SL g14548 ( 
.A(n_13731),
.B(n_13292),
.Y(n_14548)
);

OR2x2_ASAP7_75t_L g14549 ( 
.A(n_13559),
.B(n_12707),
.Y(n_14549)
);

INVx2_ASAP7_75t_L g14550 ( 
.A(n_13902),
.Y(n_14550)
);

INVx1_ASAP7_75t_L g14551 ( 
.A(n_13531),
.Y(n_14551)
);

INVx1_ASAP7_75t_L g14552 ( 
.A(n_13540),
.Y(n_14552)
);

INVx2_ASAP7_75t_L g14553 ( 
.A(n_13770),
.Y(n_14553)
);

NOR2x1_ASAP7_75t_SL g14554 ( 
.A(n_13536),
.B(n_13235),
.Y(n_14554)
);

HB1xp67_ASAP7_75t_L g14555 ( 
.A(n_13795),
.Y(n_14555)
);

AND2x2_ASAP7_75t_L g14556 ( 
.A(n_14180),
.B(n_13343),
.Y(n_14556)
);

INVxp67_ASAP7_75t_SL g14557 ( 
.A(n_13918),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_13541),
.Y(n_14558)
);

NAND2xp5_ASAP7_75t_L g14559 ( 
.A(n_14174),
.B(n_13229),
.Y(n_14559)
);

INVx2_ASAP7_75t_SL g14560 ( 
.A(n_14007),
.Y(n_14560)
);

INVx2_ASAP7_75t_L g14561 ( 
.A(n_13803),
.Y(n_14561)
);

INVx5_ASAP7_75t_SL g14562 ( 
.A(n_14114),
.Y(n_14562)
);

INVx1_ASAP7_75t_L g14563 ( 
.A(n_13546),
.Y(n_14563)
);

HB1xp67_ASAP7_75t_L g14564 ( 
.A(n_13894),
.Y(n_14564)
);

INVx3_ASAP7_75t_L g14565 ( 
.A(n_13721),
.Y(n_14565)
);

INVx1_ASAP7_75t_L g14566 ( 
.A(n_13552),
.Y(n_14566)
);

INVx2_ASAP7_75t_L g14567 ( 
.A(n_13920),
.Y(n_14567)
);

NAND2xp5_ASAP7_75t_L g14568 ( 
.A(n_14188),
.B(n_13229),
.Y(n_14568)
);

HB1xp67_ASAP7_75t_L g14569 ( 
.A(n_13848),
.Y(n_14569)
);

NAND2xp5_ASAP7_75t_L g14570 ( 
.A(n_14210),
.B(n_13224),
.Y(n_14570)
);

INVx1_ASAP7_75t_L g14571 ( 
.A(n_13565),
.Y(n_14571)
);

INVx1_ASAP7_75t_L g14572 ( 
.A(n_13571),
.Y(n_14572)
);

AND2x2_ASAP7_75t_L g14573 ( 
.A(n_14098),
.B(n_13344),
.Y(n_14573)
);

AND2x2_ASAP7_75t_L g14574 ( 
.A(n_13597),
.B(n_13583),
.Y(n_14574)
);

NOR2xp67_ASAP7_75t_L g14575 ( 
.A(n_13774),
.B(n_13147),
.Y(n_14575)
);

AOI22xp33_ASAP7_75t_L g14576 ( 
.A1(n_13510),
.A2(n_13228),
.B1(n_13381),
.B2(n_13379),
.Y(n_14576)
);

OR2x2_ASAP7_75t_L g14577 ( 
.A(n_13753),
.B(n_12713),
.Y(n_14577)
);

INVx1_ASAP7_75t_L g14578 ( 
.A(n_13572),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_13573),
.Y(n_14579)
);

INVx3_ASAP7_75t_L g14580 ( 
.A(n_13721),
.Y(n_14580)
);

INVx1_ASAP7_75t_L g14581 ( 
.A(n_13577),
.Y(n_14581)
);

INVx1_ASAP7_75t_L g14582 ( 
.A(n_13585),
.Y(n_14582)
);

INVx1_ASAP7_75t_L g14583 ( 
.A(n_13589),
.Y(n_14583)
);

INVx1_ASAP7_75t_SL g14584 ( 
.A(n_14094),
.Y(n_14584)
);

INVx4_ASAP7_75t_L g14585 ( 
.A(n_14191),
.Y(n_14585)
);

INVx1_ASAP7_75t_L g14586 ( 
.A(n_13591),
.Y(n_14586)
);

INVx2_ASAP7_75t_L g14587 ( 
.A(n_13932),
.Y(n_14587)
);

INVx2_ASAP7_75t_L g14588 ( 
.A(n_13623),
.Y(n_14588)
);

AND2x2_ASAP7_75t_L g14589 ( 
.A(n_13941),
.B(n_13409),
.Y(n_14589)
);

INVx1_ASAP7_75t_L g14590 ( 
.A(n_13594),
.Y(n_14590)
);

INVx1_ASAP7_75t_L g14591 ( 
.A(n_13595),
.Y(n_14591)
);

NOR2xp33_ASAP7_75t_L g14592 ( 
.A(n_13689),
.B(n_13293),
.Y(n_14592)
);

INVx2_ASAP7_75t_L g14593 ( 
.A(n_13623),
.Y(n_14593)
);

HB1xp67_ASAP7_75t_L g14594 ( 
.A(n_13900),
.Y(n_14594)
);

INVx1_ASAP7_75t_L g14595 ( 
.A(n_13598),
.Y(n_14595)
);

AND2x4_ASAP7_75t_L g14596 ( 
.A(n_13711),
.B(n_12858),
.Y(n_14596)
);

OR2x2_ASAP7_75t_L g14597 ( 
.A(n_13764),
.B(n_12745),
.Y(n_14597)
);

AND2x2_ASAP7_75t_L g14598 ( 
.A(n_13962),
.B(n_13648),
.Y(n_14598)
);

NAND2xp5_ASAP7_75t_L g14599 ( 
.A(n_13622),
.B(n_13175),
.Y(n_14599)
);

INVx1_ASAP7_75t_L g14600 ( 
.A(n_13606),
.Y(n_14600)
);

INVx1_ASAP7_75t_L g14601 ( 
.A(n_13612),
.Y(n_14601)
);

INVx1_ASAP7_75t_L g14602 ( 
.A(n_13615),
.Y(n_14602)
);

INVx2_ASAP7_75t_L g14603 ( 
.A(n_13663),
.Y(n_14603)
);

INVx1_ASAP7_75t_L g14604 ( 
.A(n_13616),
.Y(n_14604)
);

HB1xp67_ASAP7_75t_L g14605 ( 
.A(n_13699),
.Y(n_14605)
);

AND2x2_ASAP7_75t_L g14606 ( 
.A(n_13974),
.B(n_13211),
.Y(n_14606)
);

NAND2xp5_ASAP7_75t_L g14607 ( 
.A(n_14214),
.B(n_13223),
.Y(n_14607)
);

INVx2_ASAP7_75t_L g14608 ( 
.A(n_13663),
.Y(n_14608)
);

OR2x2_ASAP7_75t_L g14609 ( 
.A(n_13566),
.B(n_12758),
.Y(n_14609)
);

AND2x2_ASAP7_75t_L g14610 ( 
.A(n_13993),
.B(n_13297),
.Y(n_14610)
);

INVx1_ASAP7_75t_L g14611 ( 
.A(n_13618),
.Y(n_14611)
);

AND2x2_ASAP7_75t_L g14612 ( 
.A(n_13994),
.B(n_13298),
.Y(n_14612)
);

INVx1_ASAP7_75t_L g14613 ( 
.A(n_13619),
.Y(n_14613)
);

NOR2xp33_ASAP7_75t_L g14614 ( 
.A(n_13921),
.B(n_13303),
.Y(n_14614)
);

BUFx2_ASAP7_75t_L g14615 ( 
.A(n_13487),
.Y(n_14615)
);

AND2x2_ASAP7_75t_L g14616 ( 
.A(n_14006),
.B(n_13313),
.Y(n_14616)
);

INVx1_ASAP7_75t_L g14617 ( 
.A(n_13620),
.Y(n_14617)
);

AND2x2_ASAP7_75t_L g14618 ( 
.A(n_14018),
.B(n_13318),
.Y(n_14618)
);

INVx1_ASAP7_75t_L g14619 ( 
.A(n_13621),
.Y(n_14619)
);

INVx1_ASAP7_75t_L g14620 ( 
.A(n_13626),
.Y(n_14620)
);

AND2x4_ASAP7_75t_L g14621 ( 
.A(n_13717),
.B(n_12859),
.Y(n_14621)
);

NOR2xp33_ASAP7_75t_L g14622 ( 
.A(n_14194),
.B(n_13325),
.Y(n_14622)
);

INVxp67_ASAP7_75t_SL g14623 ( 
.A(n_13787),
.Y(n_14623)
);

BUFx2_ASAP7_75t_L g14624 ( 
.A(n_14048),
.Y(n_14624)
);

OAI221xp5_ASAP7_75t_SL g14625 ( 
.A1(n_13644),
.A2(n_13551),
.B1(n_13672),
.B2(n_13530),
.C(n_13611),
.Y(n_14625)
);

BUFx2_ASAP7_75t_L g14626 ( 
.A(n_13934),
.Y(n_14626)
);

HB1xp67_ASAP7_75t_L g14627 ( 
.A(n_13798),
.Y(n_14627)
);

NAND2xp5_ASAP7_75t_L g14628 ( 
.A(n_13735),
.B(n_13225),
.Y(n_14628)
);

AND2x4_ASAP7_75t_L g14629 ( 
.A(n_13718),
.B(n_14173),
.Y(n_14629)
);

BUFx2_ASAP7_75t_SL g14630 ( 
.A(n_14145),
.Y(n_14630)
);

INVx1_ASAP7_75t_SL g14631 ( 
.A(n_13690),
.Y(n_14631)
);

INVx2_ASAP7_75t_L g14632 ( 
.A(n_13732),
.Y(n_14632)
);

OR2x2_ASAP7_75t_L g14633 ( 
.A(n_14132),
.B(n_12760),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_13635),
.Y(n_14634)
);

NAND2xp5_ASAP7_75t_L g14635 ( 
.A(n_13917),
.B(n_13040),
.Y(n_14635)
);

AND2x2_ASAP7_75t_L g14636 ( 
.A(n_14026),
.B(n_13270),
.Y(n_14636)
);

AND2x2_ASAP7_75t_L g14637 ( 
.A(n_14035),
.B(n_13274),
.Y(n_14637)
);

AND2x2_ASAP7_75t_L g14638 ( 
.A(n_14037),
.B(n_13282),
.Y(n_14638)
);

HB1xp67_ASAP7_75t_L g14639 ( 
.A(n_13796),
.Y(n_14639)
);

BUFx6f_ASAP7_75t_L g14640 ( 
.A(n_13934),
.Y(n_14640)
);

OR2x2_ASAP7_75t_L g14641 ( 
.A(n_13836),
.B(n_12766),
.Y(n_14641)
);

NAND2xp5_ASAP7_75t_L g14642 ( 
.A(n_13923),
.B(n_12978),
.Y(n_14642)
);

HB1xp67_ASAP7_75t_L g14643 ( 
.A(n_13756),
.Y(n_14643)
);

NAND2xp5_ASAP7_75t_L g14644 ( 
.A(n_13924),
.B(n_12980),
.Y(n_14644)
);

AND2x2_ASAP7_75t_L g14645 ( 
.A(n_14038),
.B(n_13129),
.Y(n_14645)
);

INVx1_ASAP7_75t_L g14646 ( 
.A(n_13637),
.Y(n_14646)
);

INVx2_ASAP7_75t_L g14647 ( 
.A(n_13732),
.Y(n_14647)
);

BUFx2_ASAP7_75t_L g14648 ( 
.A(n_13940),
.Y(n_14648)
);

INVxp67_ASAP7_75t_SL g14649 ( 
.A(n_13914),
.Y(n_14649)
);

AND2x2_ASAP7_75t_L g14650 ( 
.A(n_14045),
.B(n_13143),
.Y(n_14650)
);

INVx1_ASAP7_75t_L g14651 ( 
.A(n_13642),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_13649),
.Y(n_14652)
);

BUFx3_ASAP7_75t_L g14653 ( 
.A(n_13857),
.Y(n_14653)
);

NAND2xp5_ASAP7_75t_L g14654 ( 
.A(n_13886),
.B(n_13332),
.Y(n_14654)
);

AND2x2_ASAP7_75t_L g14655 ( 
.A(n_14049),
.B(n_12870),
.Y(n_14655)
);

INVxp67_ASAP7_75t_SL g14656 ( 
.A(n_13919),
.Y(n_14656)
);

INVx2_ASAP7_75t_L g14657 ( 
.A(n_13736),
.Y(n_14657)
);

NAND2xp5_ASAP7_75t_L g14658 ( 
.A(n_13889),
.B(n_13157),
.Y(n_14658)
);

CKINVDCx14_ASAP7_75t_R g14659 ( 
.A(n_14215),
.Y(n_14659)
);

INVx1_ASAP7_75t_L g14660 ( 
.A(n_13652),
.Y(n_14660)
);

BUFx3_ASAP7_75t_L g14661 ( 
.A(n_14160),
.Y(n_14661)
);

OR2x2_ASAP7_75t_L g14662 ( 
.A(n_13671),
.B(n_13162),
.Y(n_14662)
);

AND2x2_ASAP7_75t_L g14663 ( 
.A(n_14057),
.B(n_13404),
.Y(n_14663)
);

INVx1_ASAP7_75t_L g14664 ( 
.A(n_13654),
.Y(n_14664)
);

HB1xp67_ASAP7_75t_L g14665 ( 
.A(n_13756),
.Y(n_14665)
);

BUFx2_ASAP7_75t_L g14666 ( 
.A(n_13940),
.Y(n_14666)
);

AO21x2_ASAP7_75t_L g14667 ( 
.A1(n_13580),
.A2(n_13132),
.B(n_13131),
.Y(n_14667)
);

INVx1_ASAP7_75t_L g14668 ( 
.A(n_13673),
.Y(n_14668)
);

AND2x4_ASAP7_75t_L g14669 ( 
.A(n_14161),
.B(n_13134),
.Y(n_14669)
);

OAI21x1_ASAP7_75t_L g14670 ( 
.A1(n_13939),
.A2(n_13144),
.B(n_13137),
.Y(n_14670)
);

OR2x6_ASAP7_75t_L g14671 ( 
.A(n_13613),
.B(n_13214),
.Y(n_14671)
);

INVx1_ASAP7_75t_L g14672 ( 
.A(n_13679),
.Y(n_14672)
);

AND2x4_ASAP7_75t_L g14673 ( 
.A(n_13776),
.B(n_14120),
.Y(n_14673)
);

INVx1_ASAP7_75t_L g14674 ( 
.A(n_13685),
.Y(n_14674)
);

BUFx3_ASAP7_75t_L g14675 ( 
.A(n_13517),
.Y(n_14675)
);

OR2x2_ASAP7_75t_L g14676 ( 
.A(n_14121),
.B(n_13179),
.Y(n_14676)
);

AND2x2_ASAP7_75t_L g14677 ( 
.A(n_14097),
.B(n_13136),
.Y(n_14677)
);

AOI222xp33_ASAP7_75t_L g14678 ( 
.A1(n_13494),
.A2(n_13217),
.B1(n_13294),
.B2(n_13287),
.C1(n_13101),
.C2(n_13079),
.Y(n_14678)
);

AND2x4_ASAP7_75t_L g14679 ( 
.A(n_14126),
.B(n_13161),
.Y(n_14679)
);

NAND2xp5_ASAP7_75t_L g14680 ( 
.A(n_13875),
.B(n_13182),
.Y(n_14680)
);

AND2x2_ASAP7_75t_L g14681 ( 
.A(n_14111),
.B(n_13230),
.Y(n_14681)
);

NAND2xp5_ASAP7_75t_L g14682 ( 
.A(n_13879),
.B(n_13207),
.Y(n_14682)
);

BUFx3_ASAP7_75t_L g14683 ( 
.A(n_13814),
.Y(n_14683)
);

INVx1_ASAP7_75t_L g14684 ( 
.A(n_13692),
.Y(n_14684)
);

INVx2_ASAP7_75t_L g14685 ( 
.A(n_13736),
.Y(n_14685)
);

NAND2xp5_ASAP7_75t_L g14686 ( 
.A(n_13883),
.B(n_13241),
.Y(n_14686)
);

INVx4_ASAP7_75t_L g14687 ( 
.A(n_13967),
.Y(n_14687)
);

AND2x2_ASAP7_75t_L g14688 ( 
.A(n_14112),
.B(n_13244),
.Y(n_14688)
);

INVxp67_ASAP7_75t_SL g14689 ( 
.A(n_13749),
.Y(n_14689)
);

NAND2xp5_ASAP7_75t_L g14690 ( 
.A(n_13885),
.B(n_13265),
.Y(n_14690)
);

BUFx2_ASAP7_75t_L g14691 ( 
.A(n_13967),
.Y(n_14691)
);

INVxp67_ASAP7_75t_SL g14692 ( 
.A(n_13716),
.Y(n_14692)
);

AND2x2_ASAP7_75t_L g14693 ( 
.A(n_14165),
.B(n_13268),
.Y(n_14693)
);

INVx1_ASAP7_75t_L g14694 ( 
.A(n_13696),
.Y(n_14694)
);

AOI33xp33_ASAP7_75t_L g14695 ( 
.A1(n_13811),
.A2(n_13294),
.A3(n_13287),
.B1(n_13075),
.B2(n_13092),
.B3(n_13146),
.Y(n_14695)
);

NAND2xp5_ASAP7_75t_SL g14696 ( 
.A(n_13783),
.B(n_13079),
.Y(n_14696)
);

AND2x2_ASAP7_75t_L g14697 ( 
.A(n_13979),
.B(n_13092),
.Y(n_14697)
);

INVx2_ASAP7_75t_SL g14698 ( 
.A(n_13913),
.Y(n_14698)
);

HB1xp67_ASAP7_75t_L g14699 ( 
.A(n_13767),
.Y(n_14699)
);

OR2x2_ASAP7_75t_L g14700 ( 
.A(n_14128),
.B(n_13101),
.Y(n_14700)
);

HB1xp67_ASAP7_75t_L g14701 ( 
.A(n_14130),
.Y(n_14701)
);

OAI22xp5_ASAP7_75t_L g14702 ( 
.A1(n_14105),
.A2(n_13171),
.B1(n_13174),
.B2(n_13146),
.Y(n_14702)
);

INVx2_ASAP7_75t_L g14703 ( 
.A(n_14052),
.Y(n_14703)
);

INVx2_ASAP7_75t_L g14704 ( 
.A(n_13913),
.Y(n_14704)
);

INVx1_ASAP7_75t_L g14705 ( 
.A(n_13697),
.Y(n_14705)
);

INVx5_ASAP7_75t_SL g14706 ( 
.A(n_13922),
.Y(n_14706)
);

HB1xp67_ASAP7_75t_L g14707 ( 
.A(n_14134),
.Y(n_14707)
);

AND2x2_ASAP7_75t_L g14708 ( 
.A(n_14019),
.B(n_13171),
.Y(n_14708)
);

AND2x2_ASAP7_75t_L g14709 ( 
.A(n_14178),
.B(n_13174),
.Y(n_14709)
);

AND2x2_ASAP7_75t_L g14710 ( 
.A(n_14179),
.B(n_13177),
.Y(n_14710)
);

AND2x2_ASAP7_75t_L g14711 ( 
.A(n_14192),
.B(n_13177),
.Y(n_14711)
);

BUFx2_ASAP7_75t_L g14712 ( 
.A(n_13922),
.Y(n_14712)
);

INVx2_ASAP7_75t_SL g14713 ( 
.A(n_13895),
.Y(n_14713)
);

AND2x4_ASAP7_75t_SL g14714 ( 
.A(n_13682),
.B(n_13683),
.Y(n_14714)
);

INVx2_ASAP7_75t_L g14715 ( 
.A(n_13946),
.Y(n_14715)
);

AO21x2_ASAP7_75t_L g14716 ( 
.A1(n_13488),
.A2(n_13140),
.B(n_13132),
.Y(n_14716)
);

AND2x2_ASAP7_75t_L g14717 ( 
.A(n_14198),
.B(n_13185),
.Y(n_14717)
);

NAND2xp5_ASAP7_75t_L g14718 ( 
.A(n_13837),
.B(n_13928),
.Y(n_14718)
);

BUFx6f_ASAP7_75t_L g14719 ( 
.A(n_14079),
.Y(n_14719)
);

INVxp67_ASAP7_75t_L g14720 ( 
.A(n_13925),
.Y(n_14720)
);

INVx2_ASAP7_75t_L g14721 ( 
.A(n_13948),
.Y(n_14721)
);

INVx1_ASAP7_75t_L g14722 ( 
.A(n_13702),
.Y(n_14722)
);

INVx2_ASAP7_75t_L g14723 ( 
.A(n_14127),
.Y(n_14723)
);

AND2x4_ASAP7_75t_L g14724 ( 
.A(n_14135),
.B(n_13185),
.Y(n_14724)
);

AND2x4_ASAP7_75t_L g14725 ( 
.A(n_14138),
.B(n_13189),
.Y(n_14725)
);

AND2x2_ASAP7_75t_L g14726 ( 
.A(n_14212),
.B(n_13189),
.Y(n_14726)
);

NAND2xp5_ASAP7_75t_L g14727 ( 
.A(n_13982),
.B(n_13192),
.Y(n_14727)
);

INVx1_ASAP7_75t_L g14728 ( 
.A(n_13703),
.Y(n_14728)
);

INVx1_ASAP7_75t_SL g14729 ( 
.A(n_13458),
.Y(n_14729)
);

INVx1_ASAP7_75t_L g14730 ( 
.A(n_13705),
.Y(n_14730)
);

AND2x2_ASAP7_75t_L g14731 ( 
.A(n_14219),
.B(n_13192),
.Y(n_14731)
);

OR2x2_ASAP7_75t_L g14732 ( 
.A(n_13906),
.B(n_13195),
.Y(n_14732)
);

AND2x4_ASAP7_75t_L g14733 ( 
.A(n_14146),
.B(n_13195),
.Y(n_14733)
);

OAI321xp33_ASAP7_75t_L g14734 ( 
.A1(n_13892),
.A2(n_13140),
.A3(n_13181),
.B1(n_13173),
.B2(n_13163),
.C(n_13198),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_13706),
.Y(n_14735)
);

AND2x2_ASAP7_75t_L g14736 ( 
.A(n_13607),
.B(n_13059),
.Y(n_14736)
);

AND2x2_ASAP7_75t_SL g14737 ( 
.A(n_13525),
.B(n_13212),
.Y(n_14737)
);

BUFx2_ASAP7_75t_L g14738 ( 
.A(n_13807),
.Y(n_14738)
);

HB1xp67_ASAP7_75t_L g14739 ( 
.A(n_13833),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_13712),
.Y(n_14740)
);

INVx1_ASAP7_75t_L g14741 ( 
.A(n_13722),
.Y(n_14741)
);

INVx1_ASAP7_75t_L g14742 ( 
.A(n_13728),
.Y(n_14742)
);

INVx1_ASAP7_75t_L g14743 ( 
.A(n_13738),
.Y(n_14743)
);

INVx1_ASAP7_75t_L g14744 ( 
.A(n_13740),
.Y(n_14744)
);

AND2x2_ASAP7_75t_L g14745 ( 
.A(n_14221),
.B(n_13059),
.Y(n_14745)
);

NAND2xp5_ASAP7_75t_L g14746 ( 
.A(n_13815),
.B(n_13823),
.Y(n_14746)
);

AND2x2_ASAP7_75t_L g14747 ( 
.A(n_14181),
.B(n_13063),
.Y(n_14747)
);

INVx2_ASAP7_75t_L g14748 ( 
.A(n_14190),
.Y(n_14748)
);

INVx2_ASAP7_75t_L g14749 ( 
.A(n_13949),
.Y(n_14749)
);

AND2x2_ASAP7_75t_L g14750 ( 
.A(n_14202),
.B(n_13063),
.Y(n_14750)
);

BUFx3_ASAP7_75t_L g14751 ( 
.A(n_13842),
.Y(n_14751)
);

AND2x2_ASAP7_75t_L g14752 ( 
.A(n_14213),
.B(n_13071),
.Y(n_14752)
);

INVx2_ASAP7_75t_L g14753 ( 
.A(n_14068),
.Y(n_14753)
);

AND2x4_ASAP7_75t_L g14754 ( 
.A(n_13792),
.B(n_8199),
.Y(n_14754)
);

INVx2_ASAP7_75t_L g14755 ( 
.A(n_14009),
.Y(n_14755)
);

NOR3xp33_ASAP7_75t_SL g14756 ( 
.A(n_13625),
.B(n_13071),
.C(n_6976),
.Y(n_14756)
);

AND2x2_ASAP7_75t_L g14757 ( 
.A(n_13508),
.B(n_10522),
.Y(n_14757)
);

INVx1_ASAP7_75t_SL g14758 ( 
.A(n_13849),
.Y(n_14758)
);

NAND2xp5_ASAP7_75t_L g14759 ( 
.A(n_13781),
.B(n_10522),
.Y(n_14759)
);

INVxp67_ASAP7_75t_SL g14760 ( 
.A(n_13739),
.Y(n_14760)
);

AND2x2_ASAP7_75t_L g14761 ( 
.A(n_14063),
.B(n_13570),
.Y(n_14761)
);

INVx1_ASAP7_75t_L g14762 ( 
.A(n_13751),
.Y(n_14762)
);

INVx2_ASAP7_75t_L g14763 ( 
.A(n_14013),
.Y(n_14763)
);

AND2x2_ASAP7_75t_L g14764 ( 
.A(n_14029),
.B(n_10526),
.Y(n_14764)
);

HB1xp67_ASAP7_75t_L g14765 ( 
.A(n_13675),
.Y(n_14765)
);

AND2x2_ASAP7_75t_L g14766 ( 
.A(n_14034),
.B(n_14046),
.Y(n_14766)
);

NOR2x1_ASAP7_75t_L g14767 ( 
.A(n_13752),
.B(n_10526),
.Y(n_14767)
);

NOR2xp33_ASAP7_75t_L g14768 ( 
.A(n_14168),
.B(n_8812),
.Y(n_14768)
);

AND2x2_ASAP7_75t_L g14769 ( 
.A(n_14020),
.B(n_10531),
.Y(n_14769)
);

AND2x2_ASAP7_75t_L g14770 ( 
.A(n_14024),
.B(n_10531),
.Y(n_14770)
);

INVx2_ASAP7_75t_L g14771 ( 
.A(n_14164),
.Y(n_14771)
);

OR2x2_ASAP7_75t_L g14772 ( 
.A(n_13670),
.B(n_10539),
.Y(n_14772)
);

INVxp67_ASAP7_75t_SL g14773 ( 
.A(n_13556),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_13763),
.Y(n_14774)
);

HB1xp67_ASAP7_75t_L g14775 ( 
.A(n_13854),
.Y(n_14775)
);

INVx2_ASAP7_75t_L g14776 ( 
.A(n_14086),
.Y(n_14776)
);

AND2x2_ASAP7_75t_L g14777 ( 
.A(n_14025),
.B(n_10539),
.Y(n_14777)
);

OR2x2_ASAP7_75t_L g14778 ( 
.A(n_13633),
.B(n_10540),
.Y(n_14778)
);

AND2x2_ASAP7_75t_L g14779 ( 
.A(n_14028),
.B(n_10540),
.Y(n_14779)
);

BUFx2_ASAP7_75t_L g14780 ( 
.A(n_13766),
.Y(n_14780)
);

INVx1_ASAP7_75t_L g14781 ( 
.A(n_13772),
.Y(n_14781)
);

NOR2xp33_ASAP7_75t_R g14782 ( 
.A(n_14171),
.B(n_6648),
.Y(n_14782)
);

AND2x2_ASAP7_75t_L g14783 ( 
.A(n_13548),
.B(n_13549),
.Y(n_14783)
);

HB1xp67_ASAP7_75t_L g14784 ( 
.A(n_13871),
.Y(n_14784)
);

OR2x2_ASAP7_75t_L g14785 ( 
.A(n_13775),
.B(n_10541),
.Y(n_14785)
);

NAND2xp5_ASAP7_75t_L g14786 ( 
.A(n_13788),
.B(n_10541),
.Y(n_14786)
);

HB1xp67_ASAP7_75t_L g14787 ( 
.A(n_14109),
.Y(n_14787)
);

BUFx2_ASAP7_75t_L g14788 ( 
.A(n_14169),
.Y(n_14788)
);

INVx2_ASAP7_75t_L g14789 ( 
.A(n_14090),
.Y(n_14789)
);

INVx1_ASAP7_75t_L g14790 ( 
.A(n_13651),
.Y(n_14790)
);

INVx2_ASAP7_75t_L g14791 ( 
.A(n_14092),
.Y(n_14791)
);

INVx2_ASAP7_75t_L g14792 ( 
.A(n_14099),
.Y(n_14792)
);

AND2x2_ASAP7_75t_L g14793 ( 
.A(n_13755),
.B(n_10545),
.Y(n_14793)
);

BUFx3_ASAP7_75t_L g14794 ( 
.A(n_13841),
.Y(n_14794)
);

INVxp67_ASAP7_75t_SL g14795 ( 
.A(n_14014),
.Y(n_14795)
);

INVx2_ASAP7_75t_L g14796 ( 
.A(n_14110),
.Y(n_14796)
);

AND2x2_ASAP7_75t_L g14797 ( 
.A(n_13758),
.B(n_10545),
.Y(n_14797)
);

AND2x4_ASAP7_75t_L g14798 ( 
.A(n_13933),
.B(n_8199),
.Y(n_14798)
);

INVx3_ASAP7_75t_L g14799 ( 
.A(n_13744),
.Y(n_14799)
);

AND2x2_ASAP7_75t_L g14800 ( 
.A(n_13760),
.B(n_10550),
.Y(n_14800)
);

NAND2xp5_ASAP7_75t_L g14801 ( 
.A(n_14177),
.B(n_10550),
.Y(n_14801)
);

NAND2xp5_ASAP7_75t_L g14802 ( 
.A(n_14186),
.B(n_10556),
.Y(n_14802)
);

AND2x4_ASAP7_75t_L g14803 ( 
.A(n_13725),
.B(n_8199),
.Y(n_14803)
);

AND2x2_ASAP7_75t_L g14804 ( 
.A(n_13765),
.B(n_10556),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_13657),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_13575),
.Y(n_14806)
);

AND2x2_ASAP7_75t_L g14807 ( 
.A(n_13578),
.B(n_10559),
.Y(n_14807)
);

INVx1_ASAP7_75t_L g14808 ( 
.A(n_13639),
.Y(n_14808)
);

BUFx2_ASAP7_75t_L g14809 ( 
.A(n_13452),
.Y(n_14809)
);

AND2x2_ASAP7_75t_L g14810 ( 
.A(n_14058),
.B(n_10559),
.Y(n_14810)
);

INVx2_ASAP7_75t_SL g14811 ( 
.A(n_13870),
.Y(n_14811)
);

INVx2_ASAP7_75t_L g14812 ( 
.A(n_14113),
.Y(n_14812)
);

AND2x4_ASAP7_75t_L g14813 ( 
.A(n_13727),
.B(n_8199),
.Y(n_14813)
);

OR2x6_ASAP7_75t_L g14814 ( 
.A(n_14195),
.B(n_5898),
.Y(n_14814)
);

INVx4_ASAP7_75t_L g14815 ( 
.A(n_13782),
.Y(n_14815)
);

AOI21xp33_ASAP7_75t_L g14816 ( 
.A1(n_13484),
.A2(n_10227),
.B(n_10098),
.Y(n_14816)
);

INVx2_ASAP7_75t_L g14817 ( 
.A(n_14117),
.Y(n_14817)
);

INVxp67_ASAP7_75t_SL g14818 ( 
.A(n_13631),
.Y(n_14818)
);

HB1xp67_ASAP7_75t_L g14819 ( 
.A(n_13905),
.Y(n_14819)
);

INVxp67_ASAP7_75t_SL g14820 ( 
.A(n_13665),
.Y(n_14820)
);

INVx1_ASAP7_75t_L g14821 ( 
.A(n_13839),
.Y(n_14821)
);

INVx2_ASAP7_75t_L g14822 ( 
.A(n_14119),
.Y(n_14822)
);

AND2x2_ASAP7_75t_L g14823 ( 
.A(n_13771),
.B(n_10563),
.Y(n_14823)
);

AND2x2_ASAP7_75t_L g14824 ( 
.A(n_13603),
.B(n_10563),
.Y(n_14824)
);

INVx1_ASAP7_75t_L g14825 ( 
.A(n_13666),
.Y(n_14825)
);

BUFx2_ASAP7_75t_L g14826 ( 
.A(n_13688),
.Y(n_14826)
);

INVx1_ASAP7_75t_L g14827 ( 
.A(n_13704),
.Y(n_14827)
);

AND2x2_ASAP7_75t_L g14828 ( 
.A(n_13843),
.B(n_13930),
.Y(n_14828)
);

INVx2_ASAP7_75t_L g14829 ( 
.A(n_14124),
.Y(n_14829)
);

INVx1_ASAP7_75t_L g14830 ( 
.A(n_13715),
.Y(n_14830)
);

AND2x2_ASAP7_75t_L g14831 ( 
.A(n_13911),
.B(n_13794),
.Y(n_14831)
);

AND2x2_ASAP7_75t_L g14832 ( 
.A(n_13935),
.B(n_10564),
.Y(n_14832)
);

OR2x2_ASAP7_75t_L g14833 ( 
.A(n_13658),
.B(n_10564),
.Y(n_14833)
);

BUFx2_ASAP7_75t_L g14834 ( 
.A(n_13723),
.Y(n_14834)
);

AO21x2_ASAP7_75t_L g14835 ( 
.A1(n_13646),
.A2(n_10453),
.B(n_10445),
.Y(n_14835)
);

INVx1_ASAP7_75t_L g14836 ( 
.A(n_13884),
.Y(n_14836)
);

NAND2xp5_ASAP7_75t_L g14837 ( 
.A(n_14199),
.B(n_10569),
.Y(n_14837)
);

AND2x2_ASAP7_75t_L g14838 ( 
.A(n_13614),
.B(n_10569),
.Y(n_14838)
);

INVx2_ASAP7_75t_L g14839 ( 
.A(n_14131),
.Y(n_14839)
);

AND2x2_ASAP7_75t_L g14840 ( 
.A(n_13632),
.B(n_10574),
.Y(n_14840)
);

NOR2x1p5_ASAP7_75t_L g14841 ( 
.A(n_13882),
.B(n_8282),
.Y(n_14841)
);

INVx2_ASAP7_75t_L g14842 ( 
.A(n_14137),
.Y(n_14842)
);

NOR2x1_ASAP7_75t_SL g14843 ( 
.A(n_13862),
.B(n_9134),
.Y(n_14843)
);

INVx1_ASAP7_75t_L g14844 ( 
.A(n_13887),
.Y(n_14844)
);

HB1xp67_ASAP7_75t_L g14845 ( 
.A(n_14176),
.Y(n_14845)
);

INVx2_ASAP7_75t_L g14846 ( 
.A(n_14139),
.Y(n_14846)
);

INVx2_ASAP7_75t_SL g14847 ( 
.A(n_13724),
.Y(n_14847)
);

INVx2_ASAP7_75t_L g14848 ( 
.A(n_14149),
.Y(n_14848)
);

INVx1_ASAP7_75t_L g14849 ( 
.A(n_14054),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_14056),
.Y(n_14850)
);

INVx2_ASAP7_75t_L g14851 ( 
.A(n_14066),
.Y(n_14851)
);

AND2x4_ASAP7_75t_SL g14852 ( 
.A(n_14059),
.B(n_6760),
.Y(n_14852)
);

BUFx3_ASAP7_75t_L g14853 ( 
.A(n_13741),
.Y(n_14853)
);

INVx2_ASAP7_75t_L g14854 ( 
.A(n_14067),
.Y(n_14854)
);

BUFx5_ASAP7_75t_L g14855 ( 
.A(n_13784),
.Y(n_14855)
);

AND2x2_ASAP7_75t_L g14856 ( 
.A(n_13686),
.B(n_10574),
.Y(n_14856)
);

INVx1_ASAP7_75t_L g14857 ( 
.A(n_14088),
.Y(n_14857)
);

AND2x2_ASAP7_75t_L g14858 ( 
.A(n_14183),
.B(n_10593),
.Y(n_14858)
);

NAND2xp5_ASAP7_75t_L g14859 ( 
.A(n_14204),
.B(n_10593),
.Y(n_14859)
);

OR2x2_ASAP7_75t_L g14860 ( 
.A(n_13661),
.B(n_10601),
.Y(n_14860)
);

INVx1_ASAP7_75t_L g14861 ( 
.A(n_14096),
.Y(n_14861)
);

NOR2x1_ASAP7_75t_SL g14862 ( 
.A(n_13627),
.B(n_9134),
.Y(n_14862)
);

OR2x2_ASAP7_75t_L g14863 ( 
.A(n_13938),
.B(n_10601),
.Y(n_14863)
);

INVx4_ASAP7_75t_L g14864 ( 
.A(n_13806),
.Y(n_14864)
);

AND2x2_ASAP7_75t_L g14865 ( 
.A(n_14159),
.B(n_10606),
.Y(n_14865)
);

INVx2_ASAP7_75t_L g14866 ( 
.A(n_14074),
.Y(n_14866)
);

INVxp67_ASAP7_75t_SL g14867 ( 
.A(n_14016),
.Y(n_14867)
);

AND2x2_ASAP7_75t_L g14868 ( 
.A(n_13865),
.B(n_10606),
.Y(n_14868)
);

HB1xp67_ASAP7_75t_L g14869 ( 
.A(n_14023),
.Y(n_14869)
);

AND2x2_ASAP7_75t_L g14870 ( 
.A(n_14011),
.B(n_10610),
.Y(n_14870)
);

INVx1_ASAP7_75t_L g14871 ( 
.A(n_14107),
.Y(n_14871)
);

BUFx3_ASAP7_75t_L g14872 ( 
.A(n_13742),
.Y(n_14872)
);

INVx1_ASAP7_75t_L g14873 ( 
.A(n_14108),
.Y(n_14873)
);

INVx4_ASAP7_75t_R g14874 ( 
.A(n_14205),
.Y(n_14874)
);

INVx4_ASAP7_75t_L g14875 ( 
.A(n_13808),
.Y(n_14875)
);

INVx3_ASAP7_75t_L g14876 ( 
.A(n_14185),
.Y(n_14876)
);

AND2x2_ASAP7_75t_L g14877 ( 
.A(n_14084),
.B(n_14170),
.Y(n_14877)
);

OR2x2_ASAP7_75t_L g14878 ( 
.A(n_13976),
.B(n_10610),
.Y(n_14878)
);

OR2x2_ASAP7_75t_L g14879 ( 
.A(n_13950),
.B(n_10611),
.Y(n_14879)
);

HB1xp67_ASAP7_75t_L g14880 ( 
.A(n_14015),
.Y(n_14880)
);

AND2x4_ASAP7_75t_L g14881 ( 
.A(n_13810),
.B(n_8199),
.Y(n_14881)
);

BUFx2_ASAP7_75t_L g14882 ( 
.A(n_14002),
.Y(n_14882)
);

INVx2_ASAP7_75t_L g14883 ( 
.A(n_14185),
.Y(n_14883)
);

HB1xp67_ASAP7_75t_L g14884 ( 
.A(n_13816),
.Y(n_14884)
);

INVx1_ASAP7_75t_L g14885 ( 
.A(n_14125),
.Y(n_14885)
);

BUFx2_ASAP7_75t_L g14886 ( 
.A(n_13534),
.Y(n_14886)
);

AND2x2_ASAP7_75t_L g14887 ( 
.A(n_13992),
.B(n_10611),
.Y(n_14887)
);

NOR2xp67_ASAP7_75t_L g14888 ( 
.A(n_13961),
.B(n_10625),
.Y(n_14888)
);

NAND2xp5_ASAP7_75t_L g14889 ( 
.A(n_13469),
.B(n_10625),
.Y(n_14889)
);

OAI22xp5_ASAP7_75t_SL g14890 ( 
.A1(n_13780),
.A2(n_6987),
.B1(n_10452),
.B2(n_10508),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_14140),
.Y(n_14891)
);

AND2x2_ASAP7_75t_L g14892 ( 
.A(n_14106),
.B(n_10630),
.Y(n_14892)
);

AND2x2_ASAP7_75t_L g14893 ( 
.A(n_13659),
.B(n_10630),
.Y(n_14893)
);

INVx3_ASAP7_75t_L g14894 ( 
.A(n_14151),
.Y(n_14894)
);

INVx2_ASAP7_75t_L g14895 ( 
.A(n_14201),
.Y(n_14895)
);

OR2x2_ASAP7_75t_L g14896 ( 
.A(n_13858),
.B(n_10631),
.Y(n_14896)
);

INVx3_ASAP7_75t_L g14897 ( 
.A(n_14209),
.Y(n_14897)
);

INVx2_ASAP7_75t_L g14898 ( 
.A(n_14053),
.Y(n_14898)
);

AND2x2_ASAP7_75t_L g14899 ( 
.A(n_13853),
.B(n_10631),
.Y(n_14899)
);

OR2x2_ASAP7_75t_L g14900 ( 
.A(n_13687),
.B(n_10638),
.Y(n_14900)
);

INVx1_ASAP7_75t_L g14901 ( 
.A(n_13745),
.Y(n_14901)
);

INVx2_ASAP7_75t_L g14902 ( 
.A(n_14189),
.Y(n_14902)
);

INVx1_ASAP7_75t_L g14903 ( 
.A(n_13754),
.Y(n_14903)
);

INVx1_ASAP7_75t_L g14904 ( 
.A(n_13759),
.Y(n_14904)
);

AOI22xp33_ASAP7_75t_L g14905 ( 
.A1(n_13951),
.A2(n_10227),
.B1(n_10228),
.B2(n_9994),
.Y(n_14905)
);

AND2x4_ASAP7_75t_L g14906 ( 
.A(n_13813),
.B(n_8396),
.Y(n_14906)
);

AND2x2_ASAP7_75t_L g14907 ( 
.A(n_14474),
.B(n_13840),
.Y(n_14907)
);

INVx1_ASAP7_75t_L g14908 ( 
.A(n_14266),
.Y(n_14908)
);

INVx1_ASAP7_75t_L g14909 ( 
.A(n_14266),
.Y(n_14909)
);

AND2x2_ASAP7_75t_L g14910 ( 
.A(n_14237),
.B(n_13873),
.Y(n_14910)
);

INVx2_ASAP7_75t_L g14911 ( 
.A(n_14351),
.Y(n_14911)
);

AND2x4_ASAP7_75t_L g14912 ( 
.A(n_14390),
.B(n_13817),
.Y(n_14912)
);

INVx2_ASAP7_75t_L g14913 ( 
.A(n_14309),
.Y(n_14913)
);

NAND2xp5_ASAP7_75t_L g14914 ( 
.A(n_14308),
.B(n_13908),
.Y(n_14914)
);

OR2x2_ASAP7_75t_L g14915 ( 
.A(n_14305),
.B(n_13963),
.Y(n_14915)
);

INVxp67_ASAP7_75t_L g14916 ( 
.A(n_14367),
.Y(n_14916)
);

AND2x2_ASAP7_75t_L g14917 ( 
.A(n_14257),
.B(n_13856),
.Y(n_14917)
);

OR2x2_ASAP7_75t_L g14918 ( 
.A(n_14310),
.B(n_13984),
.Y(n_14918)
);

BUFx2_ASAP7_75t_L g14919 ( 
.A(n_14289),
.Y(n_14919)
);

NAND2xp5_ASAP7_75t_SL g14920 ( 
.A(n_14447),
.B(n_14166),
.Y(n_14920)
);

AND2x2_ASAP7_75t_L g14921 ( 
.A(n_14232),
.B(n_14371),
.Y(n_14921)
);

OAI21xp5_ASAP7_75t_L g14922 ( 
.A1(n_14366),
.A2(n_13605),
.B(n_13592),
.Y(n_14922)
);

OR2x2_ASAP7_75t_L g14923 ( 
.A(n_14225),
.B(n_13987),
.Y(n_14923)
);

AND2x2_ASAP7_75t_L g14924 ( 
.A(n_14245),
.B(n_14379),
.Y(n_14924)
);

NOR2xp33_ASAP7_75t_L g14925 ( 
.A(n_14236),
.B(n_13822),
.Y(n_14925)
);

AND2x2_ASAP7_75t_L g14926 ( 
.A(n_14247),
.B(n_13824),
.Y(n_14926)
);

AND2x2_ASAP7_75t_L g14927 ( 
.A(n_14256),
.B(n_13826),
.Y(n_14927)
);

INVx1_ASAP7_75t_L g14928 ( 
.A(n_14275),
.Y(n_14928)
);

AND2x4_ASAP7_75t_L g14929 ( 
.A(n_14341),
.B(n_13831),
.Y(n_14929)
);

INVx2_ASAP7_75t_L g14930 ( 
.A(n_14309),
.Y(n_14930)
);

NAND2xp5_ASAP7_75t_L g14931 ( 
.A(n_14233),
.B(n_13762),
.Y(n_14931)
);

OR2x2_ASAP7_75t_L g14932 ( 
.A(n_14238),
.B(n_13937),
.Y(n_14932)
);

AND2x2_ASAP7_75t_L g14933 ( 
.A(n_14271),
.B(n_13834),
.Y(n_14933)
);

AND2x4_ASAP7_75t_SL g14934 ( 
.A(n_14435),
.B(n_13835),
.Y(n_14934)
);

INVx1_ASAP7_75t_L g14935 ( 
.A(n_14275),
.Y(n_14935)
);

AND2x2_ASAP7_75t_L g14936 ( 
.A(n_14365),
.B(n_14352),
.Y(n_14936)
);

HB1xp67_ASAP7_75t_L g14937 ( 
.A(n_14367),
.Y(n_14937)
);

AND2x2_ASAP7_75t_L g14938 ( 
.A(n_14322),
.B(n_14242),
.Y(n_14938)
);

INVx1_ASAP7_75t_L g14939 ( 
.A(n_14224),
.Y(n_14939)
);

OR2x2_ASAP7_75t_L g14940 ( 
.A(n_14251),
.B(n_13942),
.Y(n_14940)
);

AND2x2_ASAP7_75t_L g14941 ( 
.A(n_14458),
.B(n_14388),
.Y(n_14941)
);

NAND2xp5_ASAP7_75t_L g14942 ( 
.A(n_14564),
.B(n_13777),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_14231),
.Y(n_14943)
);

OR2x2_ASAP7_75t_L g14944 ( 
.A(n_14509),
.B(n_13779),
.Y(n_14944)
);

INVx1_ASAP7_75t_L g14945 ( 
.A(n_14263),
.Y(n_14945)
);

HB1xp67_ASAP7_75t_L g14946 ( 
.A(n_14368),
.Y(n_14946)
);

INVx1_ASAP7_75t_L g14947 ( 
.A(n_14368),
.Y(n_14947)
);

INVx1_ASAP7_75t_L g14948 ( 
.A(n_14318),
.Y(n_14948)
);

NAND3xp33_ASAP7_75t_L g14949 ( 
.A(n_14317),
.B(n_14087),
.C(n_13845),
.Y(n_14949)
);

INVx4_ASAP7_75t_L g14950 ( 
.A(n_14239),
.Y(n_14950)
);

INVx1_ASAP7_75t_L g14951 ( 
.A(n_14318),
.Y(n_14951)
);

NAND2xp5_ASAP7_75t_L g14952 ( 
.A(n_14343),
.B(n_14036),
.Y(n_14952)
);

INVx1_ASAP7_75t_L g14953 ( 
.A(n_14392),
.Y(n_14953)
);

OR2x2_ASAP7_75t_L g14954 ( 
.A(n_14533),
.B(n_13955),
.Y(n_14954)
);

NOR2x1p5_ASAP7_75t_L g14955 ( 
.A(n_14330),
.B(n_14208),
.Y(n_14955)
);

AND2x2_ASAP7_75t_L g14956 ( 
.A(n_14329),
.B(n_13838),
.Y(n_14956)
);

AND2x2_ASAP7_75t_L g14957 ( 
.A(n_14400),
.B(n_13850),
.Y(n_14957)
);

OR2x2_ASAP7_75t_L g14958 ( 
.A(n_14605),
.B(n_14197),
.Y(n_14958)
);

OR2x2_ASAP7_75t_L g14959 ( 
.A(n_14809),
.B(n_14218),
.Y(n_14959)
);

OR2x2_ASAP7_75t_L g14960 ( 
.A(n_14809),
.B(n_13859),
.Y(n_14960)
);

INVx2_ASAP7_75t_L g14961 ( 
.A(n_14626),
.Y(n_14961)
);

INVx1_ASAP7_75t_L g14962 ( 
.A(n_14403),
.Y(n_14962)
);

NAND2xp5_ASAP7_75t_L g14963 ( 
.A(n_14331),
.B(n_13867),
.Y(n_14963)
);

NAND2xp5_ASAP7_75t_L g14964 ( 
.A(n_14337),
.B(n_14323),
.Y(n_14964)
);

AND2x2_ASAP7_75t_L g14965 ( 
.A(n_14504),
.B(n_13868),
.Y(n_14965)
);

AND2x2_ASAP7_75t_L g14966 ( 
.A(n_14522),
.B(n_14574),
.Y(n_14966)
);

INVxp67_ASAP7_75t_L g14967 ( 
.A(n_14537),
.Y(n_14967)
);

AND2x2_ASAP7_75t_L g14968 ( 
.A(n_14358),
.B(n_13869),
.Y(n_14968)
);

NOR3xp33_ASAP7_75t_L g14969 ( 
.A(n_14222),
.B(n_13890),
.C(n_13872),
.Y(n_14969)
);

INVx2_ASAP7_75t_L g14970 ( 
.A(n_14626),
.Y(n_14970)
);

NAND2xp5_ASAP7_75t_L g14971 ( 
.A(n_14623),
.B(n_13891),
.Y(n_14971)
);

NAND2xp5_ASAP7_75t_L g14972 ( 
.A(n_14659),
.B(n_13893),
.Y(n_14972)
);

AND2x2_ASAP7_75t_L g14973 ( 
.A(n_14375),
.B(n_13898),
.Y(n_14973)
);

AND2x2_ASAP7_75t_L g14974 ( 
.A(n_14374),
.B(n_13901),
.Y(n_14974)
);

AND2x2_ASAP7_75t_L g14975 ( 
.A(n_14508),
.B(n_13907),
.Y(n_14975)
);

NAND2xp5_ASAP7_75t_L g14976 ( 
.A(n_14737),
.B(n_13915),
.Y(n_14976)
);

OR2x2_ASAP7_75t_L g14977 ( 
.A(n_14787),
.B(n_13916),
.Y(n_14977)
);

AND2x2_ASAP7_75t_L g14978 ( 
.A(n_14556),
.B(n_13927),
.Y(n_14978)
);

INVx1_ASAP7_75t_L g14979 ( 
.A(n_14288),
.Y(n_14979)
);

AND2x2_ASAP7_75t_L g14980 ( 
.A(n_14269),
.B(n_14381),
.Y(n_14980)
);

INVx1_ASAP7_75t_L g14981 ( 
.A(n_14301),
.Y(n_14981)
);

INVx1_ASAP7_75t_L g14982 ( 
.A(n_14228),
.Y(n_14982)
);

NAND2xp67_ASAP7_75t_L g14983 ( 
.A(n_14300),
.B(n_13929),
.Y(n_14983)
);

HB1xp67_ASAP7_75t_L g14984 ( 
.A(n_14615),
.Y(n_14984)
);

AND2x2_ASAP7_75t_L g14985 ( 
.A(n_14326),
.B(n_13931),
.Y(n_14985)
);

INVx2_ASAP7_75t_L g14986 ( 
.A(n_14691),
.Y(n_14986)
);

INVx2_ASAP7_75t_L g14987 ( 
.A(n_14691),
.Y(n_14987)
);

INVx1_ASAP7_75t_L g14988 ( 
.A(n_14234),
.Y(n_14988)
);

AND2x2_ASAP7_75t_L g14989 ( 
.A(n_14573),
.B(n_14511),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14240),
.Y(n_14990)
);

AND2x2_ASAP7_75t_L g14991 ( 
.A(n_14451),
.B(n_13947),
.Y(n_14991)
);

NAND2xp5_ASAP7_75t_L g14992 ( 
.A(n_14648),
.B(n_13953),
.Y(n_14992)
);

NAND2xp5_ASAP7_75t_SL g14993 ( 
.A(n_14353),
.B(n_13700),
.Y(n_14993)
);

AND2x2_ASAP7_75t_L g14994 ( 
.A(n_14482),
.B(n_13957),
.Y(n_14994)
);

INVx2_ASAP7_75t_SL g14995 ( 
.A(n_14353),
.Y(n_14995)
);

AND2x2_ASAP7_75t_L g14996 ( 
.A(n_14486),
.B(n_13958),
.Y(n_14996)
);

AND2x2_ASAP7_75t_L g14997 ( 
.A(n_14426),
.B(n_13960),
.Y(n_14997)
);

AND2x2_ASAP7_75t_L g14998 ( 
.A(n_14462),
.B(n_13966),
.Y(n_14998)
);

AND2x2_ASAP7_75t_L g14999 ( 
.A(n_14363),
.B(n_13973),
.Y(n_14999)
);

AND2x4_ASAP7_75t_L g15000 ( 
.A(n_14653),
.B(n_13983),
.Y(n_15000)
);

AND2x2_ASAP7_75t_L g15001 ( 
.A(n_14495),
.B(n_13986),
.Y(n_15001)
);

INVx2_ASAP7_75t_L g15002 ( 
.A(n_14241),
.Y(n_15002)
);

AND2x4_ASAP7_75t_SL g15003 ( 
.A(n_14585),
.B(n_13989),
.Y(n_15003)
);

AND2x2_ASAP7_75t_L g15004 ( 
.A(n_14468),
.B(n_14001),
.Y(n_15004)
);

OR2x2_ASAP7_75t_L g15005 ( 
.A(n_14594),
.B(n_14005),
.Y(n_15005)
);

OR2x2_ASAP7_75t_L g15006 ( 
.A(n_14264),
.B(n_14008),
.Y(n_15006)
);

INVx1_ASAP7_75t_L g15007 ( 
.A(n_14249),
.Y(n_15007)
);

INVx2_ASAP7_75t_L g15008 ( 
.A(n_14353),
.Y(n_15008)
);

INVx2_ASAP7_75t_L g15009 ( 
.A(n_14239),
.Y(n_15009)
);

AND2x4_ASAP7_75t_L g15010 ( 
.A(n_14286),
.B(n_14010),
.Y(n_15010)
);

NAND3xp33_ASAP7_75t_L g15011 ( 
.A(n_14615),
.B(n_14032),
.C(n_14027),
.Y(n_15011)
);

INVx1_ASAP7_75t_SL g15012 ( 
.A(n_14537),
.Y(n_15012)
);

AND2x2_ASAP7_75t_L g15013 ( 
.A(n_14469),
.B(n_14039),
.Y(n_15013)
);

OR2x2_ASAP7_75t_L g15014 ( 
.A(n_14265),
.B(n_14040),
.Y(n_15014)
);

INVx1_ASAP7_75t_L g15015 ( 
.A(n_14252),
.Y(n_15015)
);

NOR2xp33_ASAP7_75t_L g15016 ( 
.A(n_14321),
.B(n_14041),
.Y(n_15016)
);

NAND2xp5_ASAP7_75t_L g15017 ( 
.A(n_14666),
.B(n_14044),
.Y(n_15017)
);

AND2x2_ASAP7_75t_L g15018 ( 
.A(n_14285),
.B(n_14050),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14437),
.Y(n_15019)
);

AND2x2_ASAP7_75t_L g15020 ( 
.A(n_14418),
.B(n_14055),
.Y(n_15020)
);

NAND2xp5_ASAP7_75t_L g15021 ( 
.A(n_14712),
.B(n_14376),
.Y(n_15021)
);

AND2x4_ASAP7_75t_L g15022 ( 
.A(n_14243),
.B(n_14060),
.Y(n_15022)
);

AND2x2_ASAP7_75t_L g15023 ( 
.A(n_14282),
.B(n_14062),
.Y(n_15023)
);

INVx2_ASAP7_75t_L g15024 ( 
.A(n_14239),
.Y(n_15024)
);

OR2x2_ASAP7_75t_L g15025 ( 
.A(n_14273),
.B(n_14064),
.Y(n_15025)
);

AND2x2_ASAP7_75t_L g15026 ( 
.A(n_14290),
.B(n_14065),
.Y(n_15026)
);

AND2x2_ASAP7_75t_L g15027 ( 
.A(n_14313),
.B(n_14077),
.Y(n_15027)
);

NOR3xp33_ASAP7_75t_L g15028 ( 
.A(n_14734),
.B(n_14085),
.C(n_14082),
.Y(n_15028)
);

AND2x4_ASAP7_75t_L g15029 ( 
.A(n_14714),
.B(n_14100),
.Y(n_15029)
);

NAND2xp5_ASAP7_75t_L g15030 ( 
.A(n_14643),
.B(n_14103),
.Y(n_15030)
);

AND2x4_ASAP7_75t_L g15031 ( 
.A(n_14683),
.B(n_14104),
.Y(n_15031)
);

OR2x2_ASAP7_75t_L g15032 ( 
.A(n_14281),
.B(n_14115),
.Y(n_15032)
);

AND2x2_ASAP7_75t_L g15033 ( 
.A(n_14325),
.B(n_14116),
.Y(n_15033)
);

INVx1_ASAP7_75t_L g15034 ( 
.A(n_14471),
.Y(n_15034)
);

INVx2_ASAP7_75t_L g15035 ( 
.A(n_14255),
.Y(n_15035)
);

NAND2xp5_ASAP7_75t_L g15036 ( 
.A(n_14665),
.B(n_14118),
.Y(n_15036)
);

AND2x2_ASAP7_75t_L g15037 ( 
.A(n_14338),
.B(n_14203),
.Y(n_15037)
);

INVx2_ASAP7_75t_L g15038 ( 
.A(n_14706),
.Y(n_15038)
);

NAND2xp5_ASAP7_75t_L g15039 ( 
.A(n_14783),
.B(n_13912),
.Y(n_15039)
);

AND2x2_ASAP7_75t_L g15040 ( 
.A(n_14342),
.B(n_14148),
.Y(n_15040)
);

OR2x2_ASAP7_75t_L g15041 ( 
.A(n_14386),
.B(n_14073),
.Y(n_15041)
);

NAND2x1p5_ASAP7_75t_L g15042 ( 
.A(n_14494),
.B(n_13990),
.Y(n_15042)
);

AND2x2_ASAP7_75t_L g15043 ( 
.A(n_14356),
.B(n_13981),
.Y(n_15043)
);

INVx1_ASAP7_75t_L g15044 ( 
.A(n_14230),
.Y(n_15044)
);

INVx2_ASAP7_75t_L g15045 ( 
.A(n_14706),
.Y(n_15045)
);

INVx2_ASAP7_75t_L g15046 ( 
.A(n_14293),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_14230),
.Y(n_15047)
);

AND2x2_ASAP7_75t_L g15048 ( 
.A(n_14467),
.B(n_14033),
.Y(n_15048)
);

NAND2xp5_ASAP7_75t_L g15049 ( 
.A(n_14698),
.B(n_14047),
.Y(n_15049)
);

AND2x2_ASAP7_75t_L g15050 ( 
.A(n_14472),
.B(n_14042),
.Y(n_15050)
);

INVx1_ASAP7_75t_L g15051 ( 
.A(n_14258),
.Y(n_15051)
);

OR2x2_ASAP7_75t_L g15052 ( 
.A(n_14246),
.B(n_13995),
.Y(n_15052)
);

NAND2x1_ASAP7_75t_SL g15053 ( 
.A(n_14260),
.B(n_14307),
.Y(n_15053)
);

AND2x2_ASAP7_75t_L g15054 ( 
.A(n_14476),
.B(n_13945),
.Y(n_15054)
);

OR2x2_ASAP7_75t_L g15055 ( 
.A(n_14254),
.B(n_14021),
.Y(n_15055)
);

NAND2xp5_ASAP7_75t_L g15056 ( 
.A(n_14428),
.B(n_13969),
.Y(n_15056)
);

AND2x2_ASAP7_75t_L g15057 ( 
.A(n_14518),
.B(n_13990),
.Y(n_15057)
);

INVx1_ASAP7_75t_L g15058 ( 
.A(n_14258),
.Y(n_15058)
);

INVx1_ASAP7_75t_L g15059 ( 
.A(n_14780),
.Y(n_15059)
);

NAND2xp5_ASAP7_75t_L g15060 ( 
.A(n_14397),
.B(n_13965),
.Y(n_15060)
);

NAND2xp5_ASAP7_75t_L g15061 ( 
.A(n_14350),
.B(n_14022),
.Y(n_15061)
);

NAND2xp5_ASAP7_75t_L g15062 ( 
.A(n_14355),
.B(n_14051),
.Y(n_15062)
);

NAND2xp5_ASAP7_75t_L g15063 ( 
.A(n_14389),
.B(n_14101),
.Y(n_15063)
);

BUFx3_ASAP7_75t_L g15064 ( 
.A(n_14500),
.Y(n_15064)
);

OR2x2_ASAP7_75t_L g15065 ( 
.A(n_14332),
.B(n_14155),
.Y(n_15065)
);

NAND2xp5_ASAP7_75t_L g15066 ( 
.A(n_14562),
.B(n_14089),
.Y(n_15066)
);

AND2x2_ASAP7_75t_L g15067 ( 
.A(n_14413),
.B(n_14189),
.Y(n_15067)
);

INVxp67_ASAP7_75t_L g15068 ( 
.A(n_14554),
.Y(n_15068)
);

INVx1_ASAP7_75t_L g15069 ( 
.A(n_14780),
.Y(n_15069)
);

AOI22xp33_ASAP7_75t_L g15070 ( 
.A1(n_14548),
.A2(n_13789),
.B1(n_14196),
.B2(n_14184),
.Y(n_15070)
);

AND2x4_ASAP7_75t_L g15071 ( 
.A(n_14751),
.B(n_13997),
.Y(n_15071)
);

INVx1_ASAP7_75t_L g15072 ( 
.A(n_14364),
.Y(n_15072)
);

AOI22xp33_ASAP7_75t_L g15073 ( 
.A1(n_14277),
.A2(n_14144),
.B1(n_14122),
.B2(n_14091),
.Y(n_15073)
);

INVx1_ASAP7_75t_L g15074 ( 
.A(n_14364),
.Y(n_15074)
);

INVx2_ASAP7_75t_L g15075 ( 
.A(n_14640),
.Y(n_15075)
);

AND2x4_ASAP7_75t_L g15076 ( 
.A(n_14489),
.B(n_13997),
.Y(n_15076)
);

INVx1_ASAP7_75t_L g15077 ( 
.A(n_14422),
.Y(n_15077)
);

AND2x4_ASAP7_75t_L g15078 ( 
.A(n_14319),
.B(n_14000),
.Y(n_15078)
);

INVx1_ASAP7_75t_L g15079 ( 
.A(n_14739),
.Y(n_15079)
);

AND2x2_ASAP7_75t_L g15080 ( 
.A(n_14761),
.B(n_14129),
.Y(n_15080)
);

OR2x2_ASAP7_75t_L g15081 ( 
.A(n_14316),
.B(n_14344),
.Y(n_15081)
);

INVx1_ASAP7_75t_L g15082 ( 
.A(n_14291),
.Y(n_15082)
);

INVx1_ASAP7_75t_L g15083 ( 
.A(n_14299),
.Y(n_15083)
);

INVx3_ASAP7_75t_L g15084 ( 
.A(n_14380),
.Y(n_15084)
);

NAND2xp5_ASAP7_75t_L g15085 ( 
.A(n_14562),
.B(n_14129),
.Y(n_15085)
);

NAND2xp5_ASAP7_75t_L g15086 ( 
.A(n_14297),
.B(n_14133),
.Y(n_15086)
);

NAND2xp5_ASAP7_75t_L g15087 ( 
.A(n_14298),
.B(n_14133),
.Y(n_15087)
);

NAND2xp5_ASAP7_75t_L g15088 ( 
.A(n_14311),
.B(n_13980),
.Y(n_15088)
);

AND2x2_ASAP7_75t_L g15089 ( 
.A(n_14545),
.B(n_14000),
.Y(n_15089)
);

INVxp67_ASAP7_75t_SL g15090 ( 
.A(n_14429),
.Y(n_15090)
);

INVx1_ASAP7_75t_L g15091 ( 
.A(n_14819),
.Y(n_15091)
);

NAND2xp5_ASAP7_75t_L g15092 ( 
.A(n_14345),
.B(n_10638),
.Y(n_15092)
);

NAND2xp5_ASAP7_75t_L g15093 ( 
.A(n_14359),
.B(n_10643),
.Y(n_15093)
);

AND2x2_ASAP7_75t_L g15094 ( 
.A(n_14417),
.B(n_10643),
.Y(n_15094)
);

INVx2_ASAP7_75t_L g15095 ( 
.A(n_14640),
.Y(n_15095)
);

NAND2xp5_ASAP7_75t_L g15096 ( 
.A(n_14360),
.B(n_10645),
.Y(n_15096)
);

AND2x2_ASAP7_75t_L g15097 ( 
.A(n_14517),
.B(n_10645),
.Y(n_15097)
);

INVx2_ASAP7_75t_L g15098 ( 
.A(n_14529),
.Y(n_15098)
);

AND2x2_ASAP7_75t_L g15099 ( 
.A(n_14419),
.B(n_14423),
.Y(n_15099)
);

AND2x2_ASAP7_75t_L g15100 ( 
.A(n_14828),
.B(n_10647),
.Y(n_15100)
);

INVx4_ASAP7_75t_L g15101 ( 
.A(n_14380),
.Y(n_15101)
);

AND2x2_ASAP7_75t_L g15102 ( 
.A(n_14488),
.B(n_10647),
.Y(n_15102)
);

AND2x2_ASAP7_75t_L g15103 ( 
.A(n_14766),
.B(n_10654),
.Y(n_15103)
);

OR2x2_ASAP7_75t_L g15104 ( 
.A(n_14335),
.B(n_10654),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_14765),
.Y(n_15105)
);

INVx1_ASAP7_75t_L g15106 ( 
.A(n_14624),
.Y(n_15106)
);

AND2x2_ASAP7_75t_L g15107 ( 
.A(n_14598),
.B(n_10673),
.Y(n_15107)
);

INVx2_ASAP7_75t_L g15108 ( 
.A(n_14546),
.Y(n_15108)
);

NAND2xp5_ASAP7_75t_L g15109 ( 
.A(n_14627),
.B(n_10673),
.Y(n_15109)
);

INVx2_ASAP7_75t_L g15110 ( 
.A(n_14565),
.Y(n_15110)
);

OR2x2_ASAP7_75t_L g15111 ( 
.A(n_14244),
.B(n_10681),
.Y(n_15111)
);

AND2x2_ASAP7_75t_L g15112 ( 
.A(n_14327),
.B(n_14312),
.Y(n_15112)
);

NAND2xp5_ASAP7_75t_L g15113 ( 
.A(n_14382),
.B(n_10681),
.Y(n_15113)
);

AND2x2_ASAP7_75t_L g15114 ( 
.A(n_14490),
.B(n_10688),
.Y(n_15114)
);

INVx1_ASAP7_75t_L g15115 ( 
.A(n_14624),
.Y(n_15115)
);

NOR2xp33_ASAP7_75t_L g15116 ( 
.A(n_14433),
.B(n_10688),
.Y(n_15116)
);

HB1xp67_ASAP7_75t_L g15117 ( 
.A(n_14340),
.Y(n_15117)
);

OR2x2_ASAP7_75t_L g15118 ( 
.A(n_14315),
.B(n_10690),
.Y(n_15118)
);

INVx2_ASAP7_75t_L g15119 ( 
.A(n_14580),
.Y(n_15119)
);

AND2x2_ASAP7_75t_L g15120 ( 
.A(n_14831),
.B(n_10690),
.Y(n_15120)
);

NAND2xp5_ASAP7_75t_SL g15121 ( 
.A(n_14369),
.B(n_8282),
.Y(n_15121)
);

NAND2xp5_ASAP7_75t_L g15122 ( 
.A(n_14383),
.B(n_10699),
.Y(n_15122)
);

NAND2x1_ASAP7_75t_L g15123 ( 
.A(n_14874),
.B(n_10508),
.Y(n_15123)
);

NAND2x1p5_ASAP7_75t_L g15124 ( 
.A(n_14369),
.B(n_8329),
.Y(n_15124)
);

INVx1_ASAP7_75t_L g15125 ( 
.A(n_14701),
.Y(n_15125)
);

NOR2xp67_ASAP7_75t_L g15126 ( 
.A(n_14399),
.B(n_10699),
.Y(n_15126)
);

OR2x2_ASAP7_75t_L g15127 ( 
.A(n_14336),
.B(n_14223),
.Y(n_15127)
);

INVx1_ASAP7_75t_L g15128 ( 
.A(n_14707),
.Y(n_15128)
);

AND2x4_ASAP7_75t_L g15129 ( 
.A(n_14373),
.B(n_8396),
.Y(n_15129)
);

INVx1_ASAP7_75t_L g15130 ( 
.A(n_14569),
.Y(n_15130)
);

INVx1_ASAP7_75t_L g15131 ( 
.A(n_14882),
.Y(n_15131)
);

NAND2xp5_ASAP7_75t_SL g15132 ( 
.A(n_14279),
.B(n_8329),
.Y(n_15132)
);

OR2x2_ASAP7_75t_L g15133 ( 
.A(n_14394),
.B(n_10704),
.Y(n_15133)
);

INVx2_ASAP7_75t_L g15134 ( 
.A(n_14876),
.Y(n_15134)
);

OR2x2_ASAP7_75t_L g15135 ( 
.A(n_14487),
.B(n_10704),
.Y(n_15135)
);

BUFx2_ASAP7_75t_L g15136 ( 
.A(n_14438),
.Y(n_15136)
);

AND2x4_ASAP7_75t_L g15137 ( 
.A(n_14713),
.B(n_8396),
.Y(n_15137)
);

INVx1_ASAP7_75t_L g15138 ( 
.A(n_14882),
.Y(n_15138)
);

AND2x4_ASAP7_75t_L g15139 ( 
.A(n_14296),
.B(n_8396),
.Y(n_15139)
);

INVx1_ASAP7_75t_L g15140 ( 
.A(n_14775),
.Y(n_15140)
);

AND2x2_ASAP7_75t_L g15141 ( 
.A(n_14276),
.B(n_10705),
.Y(n_15141)
);

INVx1_ASAP7_75t_L g15142 ( 
.A(n_14784),
.Y(n_15142)
);

OR2x2_ASAP7_75t_L g15143 ( 
.A(n_14446),
.B(n_14253),
.Y(n_15143)
);

OR2x2_ASAP7_75t_L g15144 ( 
.A(n_14324),
.B(n_10705),
.Y(n_15144)
);

OR2x2_ASAP7_75t_L g15145 ( 
.A(n_14729),
.B(n_14284),
.Y(n_15145)
);

AND2x2_ASAP7_75t_L g15146 ( 
.A(n_14456),
.B(n_10709),
.Y(n_15146)
);

INVx2_ASAP7_75t_L g15147 ( 
.A(n_14520),
.Y(n_15147)
);

NOR2x1_ASAP7_75t_L g15148 ( 
.A(n_14292),
.B(n_10709),
.Y(n_15148)
);

AOI211xp5_ASAP7_75t_L g15149 ( 
.A1(n_14625),
.A2(n_10383),
.B(n_10405),
.C(n_10393),
.Y(n_15149)
);

NAND2xp5_ASAP7_75t_L g15150 ( 
.A(n_14588),
.B(n_10710),
.Y(n_15150)
);

NAND2xp5_ASAP7_75t_L g15151 ( 
.A(n_14593),
.B(n_14603),
.Y(n_15151)
);

OR2x2_ASAP7_75t_L g15152 ( 
.A(n_14457),
.B(n_10710),
.Y(n_15152)
);

AND2x2_ASAP7_75t_L g15153 ( 
.A(n_14535),
.B(n_10713),
.Y(n_15153)
);

NAND2x1p5_ASAP7_75t_L g15154 ( 
.A(n_14687),
.B(n_8329),
.Y(n_15154)
);

AND2x2_ASAP7_75t_L g15155 ( 
.A(n_14539),
.B(n_10713),
.Y(n_15155)
);

OR2x2_ASAP7_75t_L g15156 ( 
.A(n_14463),
.B(n_10718),
.Y(n_15156)
);

HB1xp67_ASAP7_75t_L g15157 ( 
.A(n_14575),
.Y(n_15157)
);

NAND2xp5_ASAP7_75t_L g15158 ( 
.A(n_14608),
.B(n_10718),
.Y(n_15158)
);

NAND2xp5_ASAP7_75t_L g15159 ( 
.A(n_14699),
.B(n_10720),
.Y(n_15159)
);

AND2x2_ASAP7_75t_L g15160 ( 
.A(n_14430),
.B(n_10720),
.Y(n_15160)
);

NAND2xp5_ASAP7_75t_L g15161 ( 
.A(n_14339),
.B(n_10723),
.Y(n_15161)
);

AND2x2_ASAP7_75t_L g15162 ( 
.A(n_14443),
.B(n_14589),
.Y(n_15162)
);

AND2x4_ASAP7_75t_L g15163 ( 
.A(n_14704),
.B(n_11160),
.Y(n_15163)
);

AND2x2_ASAP7_75t_L g15164 ( 
.A(n_14348),
.B(n_14354),
.Y(n_15164)
);

OR2x2_ASAP7_75t_L g15165 ( 
.A(n_14304),
.B(n_14259),
.Y(n_15165)
);

AND2x2_ASAP7_75t_L g15166 ( 
.A(n_14596),
.B(n_10723),
.Y(n_15166)
);

NAND2xp5_ASAP7_75t_L g15167 ( 
.A(n_14370),
.B(n_10730),
.Y(n_15167)
);

NAND2xp5_ASAP7_75t_L g15168 ( 
.A(n_14270),
.B(n_10730),
.Y(n_15168)
);

INVx1_ASAP7_75t_L g15169 ( 
.A(n_14709),
.Y(n_15169)
);

NAND2xp5_ASAP7_75t_L g15170 ( 
.A(n_14514),
.B(n_10732),
.Y(n_15170)
);

AND2x2_ASAP7_75t_L g15171 ( 
.A(n_14621),
.B(n_10732),
.Y(n_15171)
);

AND2x2_ASAP7_75t_L g15172 ( 
.A(n_14334),
.B(n_10747),
.Y(n_15172)
);

INVx2_ASAP7_75t_SL g15173 ( 
.A(n_14274),
.Y(n_15173)
);

NAND2xp5_ASAP7_75t_L g15174 ( 
.A(n_14632),
.B(n_10747),
.Y(n_15174)
);

INVx1_ASAP7_75t_L g15175 ( 
.A(n_14710),
.Y(n_15175)
);

INVx1_ASAP7_75t_L g15176 ( 
.A(n_14248),
.Y(n_15176)
);

INVx2_ASAP7_75t_L g15177 ( 
.A(n_14387),
.Y(n_15177)
);

INVx2_ASAP7_75t_L g15178 ( 
.A(n_14387),
.Y(n_15178)
);

NOR2x1_ASAP7_75t_L g15179 ( 
.A(n_14667),
.B(n_10755),
.Y(n_15179)
);

AND2x2_ASAP7_75t_L g15180 ( 
.A(n_14481),
.B(n_10755),
.Y(n_15180)
);

AND2x2_ASAP7_75t_L g15181 ( 
.A(n_14485),
.B(n_10756),
.Y(n_15181)
);

NAND2xp5_ASAP7_75t_L g15182 ( 
.A(n_14647),
.B(n_10756),
.Y(n_15182)
);

INVx1_ASAP7_75t_L g15183 ( 
.A(n_14248),
.Y(n_15183)
);

INVx2_ASAP7_75t_L g15184 ( 
.A(n_14274),
.Y(n_15184)
);

AND2x2_ASAP7_75t_L g15185 ( 
.A(n_14306),
.B(n_14675),
.Y(n_15185)
);

OR2x2_ASAP7_75t_L g15186 ( 
.A(n_14295),
.B(n_10761),
.Y(n_15186)
);

INVx1_ASAP7_75t_L g15187 ( 
.A(n_14724),
.Y(n_15187)
);

NAND2xp5_ASAP7_75t_L g15188 ( 
.A(n_14657),
.B(n_10761),
.Y(n_15188)
);

INVx1_ASAP7_75t_L g15189 ( 
.A(n_14725),
.Y(n_15189)
);

INVx1_ASAP7_75t_L g15190 ( 
.A(n_14733),
.Y(n_15190)
);

NAND2xp5_ASAP7_75t_L g15191 ( 
.A(n_14685),
.B(n_10762),
.Y(n_15191)
);

INVx1_ASAP7_75t_L g15192 ( 
.A(n_14639),
.Y(n_15192)
);

AND2x2_ASAP7_75t_L g15193 ( 
.A(n_14544),
.B(n_10762),
.Y(n_15193)
);

INVx1_ASAP7_75t_L g15194 ( 
.A(n_14700),
.Y(n_15194)
);

NAND2xp5_ASAP7_75t_L g15195 ( 
.A(n_14513),
.B(n_10766),
.Y(n_15195)
);

INVx1_ASAP7_75t_L g15196 ( 
.A(n_14697),
.Y(n_15196)
);

INVx1_ASAP7_75t_L g15197 ( 
.A(n_14333),
.Y(n_15197)
);

AND2x4_ASAP7_75t_L g15198 ( 
.A(n_14384),
.B(n_11160),
.Y(n_15198)
);

INVx1_ASAP7_75t_L g15199 ( 
.A(n_14314),
.Y(n_15199)
);

INVx2_ASAP7_75t_L g15200 ( 
.A(n_14328),
.Y(n_15200)
);

AND2x4_ASAP7_75t_L g15201 ( 
.A(n_14395),
.B(n_11199),
.Y(n_15201)
);

INVx2_ASAP7_75t_L g15202 ( 
.A(n_14328),
.Y(n_15202)
);

HB1xp67_ASAP7_75t_L g15203 ( 
.A(n_14459),
.Y(n_15203)
);

NAND2xp5_ASAP7_75t_L g15204 ( 
.A(n_14788),
.B(n_10766),
.Y(n_15204)
);

INVx1_ASAP7_75t_L g15205 ( 
.A(n_14555),
.Y(n_15205)
);

AND2x2_ASAP7_75t_L g15206 ( 
.A(n_14302),
.B(n_10772),
.Y(n_15206)
);

OR2x2_ASAP7_75t_L g15207 ( 
.A(n_14642),
.B(n_10772),
.Y(n_15207)
);

INVx2_ASAP7_75t_L g15208 ( 
.A(n_14855),
.Y(n_15208)
);

BUFx2_ASAP7_75t_L g15209 ( 
.A(n_14557),
.Y(n_15209)
);

INVx1_ASAP7_75t_L g15210 ( 
.A(n_14689),
.Y(n_15210)
);

HB1xp67_ASAP7_75t_L g15211 ( 
.A(n_14473),
.Y(n_15211)
);

AND2x2_ASAP7_75t_L g15212 ( 
.A(n_14525),
.B(n_10777),
.Y(n_15212)
);

INVx1_ASAP7_75t_L g15213 ( 
.A(n_14692),
.Y(n_15213)
);

AND2x2_ASAP7_75t_L g15214 ( 
.A(n_14531),
.B(n_10777),
.Y(n_15214)
);

INVx2_ASAP7_75t_L g15215 ( 
.A(n_14855),
.Y(n_15215)
);

INVx2_ASAP7_75t_L g15216 ( 
.A(n_14855),
.Y(n_15216)
);

NAND2xp5_ASAP7_75t_L g15217 ( 
.A(n_14788),
.B(n_10779),
.Y(n_15217)
);

INVx1_ASAP7_75t_L g15218 ( 
.A(n_14261),
.Y(n_15218)
);

INVx1_ASAP7_75t_L g15219 ( 
.A(n_14267),
.Y(n_15219)
);

INVx2_ASAP7_75t_L g15220 ( 
.A(n_14855),
.Y(n_15220)
);

OR2x2_ASAP7_75t_L g15221 ( 
.A(n_14644),
.B(n_10779),
.Y(n_15221)
);

HB1xp67_ASAP7_75t_L g15222 ( 
.A(n_14671),
.Y(n_15222)
);

INVx1_ASAP7_75t_L g15223 ( 
.A(n_14527),
.Y(n_15223)
);

INVx1_ASAP7_75t_L g15224 ( 
.A(n_14530),
.Y(n_15224)
);

AND2x2_ASAP7_75t_L g15225 ( 
.A(n_14515),
.B(n_10796),
.Y(n_15225)
);

INVx2_ASAP7_75t_L g15226 ( 
.A(n_14401),
.Y(n_15226)
);

AND2x2_ASAP7_75t_L g15227 ( 
.A(n_14492),
.B(n_10796),
.Y(n_15227)
);

INVx2_ASAP7_75t_L g15228 ( 
.A(n_14404),
.Y(n_15228)
);

CKINVDCx14_ASAP7_75t_R g15229 ( 
.A(n_14294),
.Y(n_15229)
);

AND2x2_ASAP7_75t_L g15230 ( 
.A(n_14499),
.B(n_10799),
.Y(n_15230)
);

NAND2xp5_ASAP7_75t_L g15231 ( 
.A(n_14799),
.B(n_10799),
.Y(n_15231)
);

NAND2xp5_ASAP7_75t_L g15232 ( 
.A(n_14226),
.B(n_10817),
.Y(n_15232)
);

NAND2xp5_ASAP7_75t_SL g15233 ( 
.A(n_14719),
.B(n_8329),
.Y(n_15233)
);

AND2x2_ASAP7_75t_L g15234 ( 
.A(n_14503),
.B(n_10817),
.Y(n_15234)
);

INVx1_ASAP7_75t_L g15235 ( 
.A(n_14268),
.Y(n_15235)
);

INVx1_ASAP7_75t_L g15236 ( 
.A(n_14272),
.Y(n_15236)
);

INVx1_ASAP7_75t_L g15237 ( 
.A(n_14280),
.Y(n_15237)
);

AND2x2_ASAP7_75t_L g15238 ( 
.A(n_14655),
.B(n_14610),
.Y(n_15238)
);

OR2x2_ASAP7_75t_L g15239 ( 
.A(n_14408),
.B(n_10828),
.Y(n_15239)
);

INVx1_ASAP7_75t_L g15240 ( 
.A(n_14283),
.Y(n_15240)
);

NAND2xp5_ASAP7_75t_L g15241 ( 
.A(n_14811),
.B(n_10828),
.Y(n_15241)
);

INVx2_ASAP7_75t_L g15242 ( 
.A(n_14902),
.Y(n_15242)
);

CKINVDCx11_ASAP7_75t_R g15243 ( 
.A(n_14719),
.Y(n_15243)
);

AND2x4_ASAP7_75t_L g15244 ( 
.A(n_14629),
.B(n_11199),
.Y(n_15244)
);

AND2x2_ASAP7_75t_L g15245 ( 
.A(n_14612),
.B(n_10831),
.Y(n_15245)
);

HB1xp67_ASAP7_75t_L g15246 ( 
.A(n_14671),
.Y(n_15246)
);

AND2x2_ASAP7_75t_L g15247 ( 
.A(n_14616),
.B(n_14618),
.Y(n_15247)
);

INVx2_ASAP7_75t_L g15248 ( 
.A(n_14883),
.Y(n_15248)
);

INVx1_ASAP7_75t_L g15249 ( 
.A(n_14497),
.Y(n_15249)
);

OR2x2_ASAP7_75t_L g15250 ( 
.A(n_14409),
.B(n_10831),
.Y(n_15250)
);

AND2x4_ASAP7_75t_L g15251 ( 
.A(n_14661),
.B(n_8396),
.Y(n_15251)
);

AND2x4_ASAP7_75t_L g15252 ( 
.A(n_14442),
.B(n_8436),
.Y(n_15252)
);

NAND2xp5_ASAP7_75t_L g15253 ( 
.A(n_14250),
.B(n_10836),
.Y(n_15253)
);

AND2x2_ASAP7_75t_L g15254 ( 
.A(n_14636),
.B(n_10836),
.Y(n_15254)
);

INVx2_ASAP7_75t_L g15255 ( 
.A(n_14357),
.Y(n_15255)
);

NAND2xp5_ASAP7_75t_L g15256 ( 
.A(n_14448),
.B(n_10837),
.Y(n_15256)
);

AND2x4_ASAP7_75t_L g15257 ( 
.A(n_14567),
.B(n_8436),
.Y(n_15257)
);

INVx1_ASAP7_75t_L g15258 ( 
.A(n_14431),
.Y(n_15258)
);

AND2x4_ASAP7_75t_SL g15259 ( 
.A(n_14673),
.B(n_6760),
.Y(n_15259)
);

INVxp67_ASAP7_75t_SL g15260 ( 
.A(n_14406),
.Y(n_15260)
);

AND2x2_ASAP7_75t_L g15261 ( 
.A(n_14637),
.B(n_10837),
.Y(n_15261)
);

INVx2_ASAP7_75t_L g15262 ( 
.A(n_14425),
.Y(n_15262)
);

AND2x2_ASAP7_75t_L g15263 ( 
.A(n_14638),
.B(n_10841),
.Y(n_15263)
);

AND2x2_ASAP7_75t_L g15264 ( 
.A(n_14645),
.B(n_10841),
.Y(n_15264)
);

OR2x2_ASAP7_75t_L g15265 ( 
.A(n_14758),
.B(n_10843),
.Y(n_15265)
);

AND2x2_ASAP7_75t_L g15266 ( 
.A(n_14650),
.B(n_10843),
.Y(n_15266)
);

AND2x2_ASAP7_75t_L g15267 ( 
.A(n_14496),
.B(n_14542),
.Y(n_15267)
);

INVx1_ASAP7_75t_L g15268 ( 
.A(n_14362),
.Y(n_15268)
);

INVx1_ASAP7_75t_L g15269 ( 
.A(n_14745),
.Y(n_15269)
);

NOR2xp33_ASAP7_75t_L g15270 ( 
.A(n_14262),
.B(n_10848),
.Y(n_15270)
);

CKINVDCx5p33_ASAP7_75t_R g15271 ( 
.A(n_14630),
.Y(n_15271)
);

INVx2_ASAP7_75t_L g15272 ( 
.A(n_14843),
.Y(n_15272)
);

HB1xp67_ASAP7_75t_L g15273 ( 
.A(n_14894),
.Y(n_15273)
);

INVx1_ASAP7_75t_L g15274 ( 
.A(n_14747),
.Y(n_15274)
);

INVx1_ASAP7_75t_L g15275 ( 
.A(n_14750),
.Y(n_15275)
);

AND2x2_ASAP7_75t_L g15276 ( 
.A(n_14663),
.B(n_10848),
.Y(n_15276)
);

INVx1_ASAP7_75t_L g15277 ( 
.A(n_14752),
.Y(n_15277)
);

INVx3_ASAP7_75t_L g15278 ( 
.A(n_14372),
.Y(n_15278)
);

AND2x2_ASAP7_75t_L g15279 ( 
.A(n_14606),
.B(n_10852),
.Y(n_15279)
);

OAI21xp33_ASAP7_75t_L g15280 ( 
.A1(n_14229),
.A2(n_10854),
.B(n_10852),
.Y(n_15280)
);

INVx2_ASAP7_75t_L g15281 ( 
.A(n_14862),
.Y(n_15281)
);

NAND3xp33_ASAP7_75t_L g15282 ( 
.A(n_14449),
.B(n_14405),
.C(n_14227),
.Y(n_15282)
);

INVx1_ASAP7_75t_L g15283 ( 
.A(n_14347),
.Y(n_15283)
);

NAND2xp5_ASAP7_75t_L g15284 ( 
.A(n_14421),
.B(n_10854),
.Y(n_15284)
);

AND2x4_ASAP7_75t_SL g15285 ( 
.A(n_14541),
.B(n_6760),
.Y(n_15285)
);

OR2x6_ASAP7_75t_L g15286 ( 
.A(n_14278),
.B(n_6172),
.Y(n_15286)
);

OR2x2_ASAP7_75t_L g15287 ( 
.A(n_14654),
.B(n_10860),
.Y(n_15287)
);

NAND2xp5_ASAP7_75t_L g15288 ( 
.A(n_14679),
.B(n_10860),
.Y(n_15288)
);

BUFx4f_ASAP7_75t_L g15289 ( 
.A(n_14553),
.Y(n_15289)
);

INVx2_ASAP7_75t_L g15290 ( 
.A(n_14897),
.Y(n_15290)
);

INVx1_ASAP7_75t_L g15291 ( 
.A(n_14349),
.Y(n_15291)
);

INVx1_ASAP7_75t_L g15292 ( 
.A(n_14688),
.Y(n_15292)
);

OR2x2_ASAP7_75t_L g15293 ( 
.A(n_14570),
.B(n_10863),
.Y(n_15293)
);

AND2x2_ASAP7_75t_L g15294 ( 
.A(n_14235),
.B(n_10863),
.Y(n_15294)
);

INVx1_ASAP7_75t_L g15295 ( 
.A(n_14693),
.Y(n_15295)
);

OR2x6_ASAP7_75t_L g15296 ( 
.A(n_14378),
.B(n_6188),
.Y(n_15296)
);

OR2x2_ASAP7_75t_L g15297 ( 
.A(n_14587),
.B(n_10865),
.Y(n_15297)
);

OR2x2_ASAP7_75t_L g15298 ( 
.A(n_14346),
.B(n_10865),
.Y(n_15298)
);

OR2x2_ASAP7_75t_L g15299 ( 
.A(n_14411),
.B(n_10874),
.Y(n_15299)
);

NAND2xp5_ASAP7_75t_L g15300 ( 
.A(n_14424),
.B(n_10874),
.Y(n_15300)
);

HB1xp67_ASAP7_75t_L g15301 ( 
.A(n_14708),
.Y(n_15301)
);

AND2x2_ASAP7_75t_L g15302 ( 
.A(n_14715),
.B(n_14721),
.Y(n_15302)
);

NAND2x1p5_ASAP7_75t_L g15303 ( 
.A(n_14631),
.B(n_8329),
.Y(n_15303)
);

INVx1_ASAP7_75t_L g15304 ( 
.A(n_14559),
.Y(n_15304)
);

AND2x2_ASAP7_75t_L g15305 ( 
.A(n_14749),
.B(n_10878),
.Y(n_15305)
);

AND2x4_ASAP7_75t_L g15306 ( 
.A(n_14847),
.B(n_11208),
.Y(n_15306)
);

NAND2xp5_ASAP7_75t_L g15307 ( 
.A(n_14711),
.B(n_10878),
.Y(n_15307)
);

AND2x2_ASAP7_75t_L g15308 ( 
.A(n_14755),
.B(n_14771),
.Y(n_15308)
);

OR2x2_ASAP7_75t_L g15309 ( 
.A(n_14561),
.B(n_10882),
.Y(n_15309)
);

NAND2xp5_ASAP7_75t_L g15310 ( 
.A(n_14717),
.B(n_10882),
.Y(n_15310)
);

INVx1_ASAP7_75t_L g15311 ( 
.A(n_14795),
.Y(n_15311)
);

INVx2_ASAP7_75t_L g15312 ( 
.A(n_14877),
.Y(n_15312)
);

NAND2x1_ASAP7_75t_L g15313 ( 
.A(n_14498),
.B(n_10508),
.Y(n_15313)
);

INVx1_ASAP7_75t_L g15314 ( 
.A(n_14676),
.Y(n_15314)
);

INVx1_ASAP7_75t_L g15315 ( 
.A(n_14420),
.Y(n_15315)
);

INVx2_ASAP7_75t_L g15316 ( 
.A(n_14731),
.Y(n_15316)
);

AND2x2_ASAP7_75t_L g15317 ( 
.A(n_14763),
.B(n_10896),
.Y(n_15317)
);

HB1xp67_ASAP7_75t_L g15318 ( 
.A(n_14826),
.Y(n_15318)
);

AND2x2_ASAP7_75t_L g15319 ( 
.A(n_14703),
.B(n_10896),
.Y(n_15319)
);

INVx1_ASAP7_75t_L g15320 ( 
.A(n_14501),
.Y(n_15320)
);

INVx1_ASAP7_75t_L g15321 ( 
.A(n_14726),
.Y(n_15321)
);

AND2x2_ASAP7_75t_L g15322 ( 
.A(n_14723),
.B(n_10899),
.Y(n_15322)
);

AND2x2_ASAP7_75t_L g15323 ( 
.A(n_14895),
.B(n_10899),
.Y(n_15323)
);

OR2x2_ASAP7_75t_L g15324 ( 
.A(n_14534),
.B(n_10903),
.Y(n_15324)
);

AND2x2_ASAP7_75t_L g15325 ( 
.A(n_14753),
.B(n_10903),
.Y(n_15325)
);

OR2x2_ASAP7_75t_L g15326 ( 
.A(n_14658),
.B(n_10910),
.Y(n_15326)
);

AND2x4_ASAP7_75t_SL g15327 ( 
.A(n_14748),
.B(n_6907),
.Y(n_15327)
);

AND2x4_ASAP7_75t_L g15328 ( 
.A(n_14505),
.B(n_8436),
.Y(n_15328)
);

INVxp67_ASAP7_75t_L g15329 ( 
.A(n_14738),
.Y(n_15329)
);

AND2x2_ASAP7_75t_L g15330 ( 
.A(n_14776),
.B(n_10910),
.Y(n_15330)
);

INVx1_ASAP7_75t_L g15331 ( 
.A(n_14568),
.Y(n_15331)
);

INVx1_ASAP7_75t_L g15332 ( 
.A(n_14732),
.Y(n_15332)
);

NAND2xp5_ASAP7_75t_L g15333 ( 
.A(n_14736),
.B(n_10927),
.Y(n_15333)
);

INVx1_ASAP7_75t_L g15334 ( 
.A(n_14790),
.Y(n_15334)
);

AND2x2_ASAP7_75t_L g15335 ( 
.A(n_14789),
.B(n_10927),
.Y(n_15335)
);

INVx2_ASAP7_75t_L g15336 ( 
.A(n_14464),
.Y(n_15336)
);

INVx1_ASAP7_75t_L g15337 ( 
.A(n_14805),
.Y(n_15337)
);

OR2x2_ASAP7_75t_L g15338 ( 
.A(n_14680),
.B(n_10931),
.Y(n_15338)
);

NOR2x1_ASAP7_75t_L g15339 ( 
.A(n_14506),
.B(n_10931),
.Y(n_15339)
);

NOR2xp33_ASAP7_75t_L g15340 ( 
.A(n_14720),
.B(n_10932),
.Y(n_15340)
);

INVx2_ASAP7_75t_L g15341 ( 
.A(n_14479),
.Y(n_15341)
);

NAND2xp5_ASAP7_75t_L g15342 ( 
.A(n_14773),
.B(n_14412),
.Y(n_15342)
);

AND2x2_ASAP7_75t_L g15343 ( 
.A(n_14791),
.B(n_10932),
.Y(n_15343)
);

INVx1_ASAP7_75t_L g15344 ( 
.A(n_14836),
.Y(n_15344)
);

NAND2xp5_ASAP7_75t_L g15345 ( 
.A(n_14886),
.B(n_10935),
.Y(n_15345)
);

INVx1_ASAP7_75t_L g15346 ( 
.A(n_14844),
.Y(n_15346)
);

HB1xp67_ASAP7_75t_L g15347 ( 
.A(n_14826),
.Y(n_15347)
);

INVx1_ASAP7_75t_L g15348 ( 
.A(n_14577),
.Y(n_15348)
);

AND2x4_ASAP7_75t_SL g15349 ( 
.A(n_14560),
.B(n_6907),
.Y(n_15349)
);

BUFx2_ASAP7_75t_L g15350 ( 
.A(n_14738),
.Y(n_15350)
);

INVx2_ASAP7_75t_L g15351 ( 
.A(n_14669),
.Y(n_15351)
);

NAND2xp5_ASAP7_75t_L g15352 ( 
.A(n_14886),
.B(n_10935),
.Y(n_15352)
);

NOR2xp33_ASAP7_75t_L g15353 ( 
.A(n_14493),
.B(n_10939),
.Y(n_15353)
);

INVx2_ASAP7_75t_L g15354 ( 
.A(n_14516),
.Y(n_15354)
);

INVx1_ASAP7_75t_L g15355 ( 
.A(n_14597),
.Y(n_15355)
);

AND2x4_ASAP7_75t_L g15356 ( 
.A(n_14521),
.B(n_8436),
.Y(n_15356)
);

AND2x4_ASAP7_75t_SL g15357 ( 
.A(n_14815),
.B(n_6907),
.Y(n_15357)
);

NAND2xp5_ASAP7_75t_L g15358 ( 
.A(n_14576),
.B(n_10939),
.Y(n_15358)
);

AND2x4_ASAP7_75t_L g15359 ( 
.A(n_14528),
.B(n_8436),
.Y(n_15359)
);

OR2x2_ASAP7_75t_L g15360 ( 
.A(n_14682),
.B(n_10941),
.Y(n_15360)
);

AND2x2_ASAP7_75t_L g15361 ( 
.A(n_14792),
.B(n_10941),
.Y(n_15361)
);

INVx1_ASAP7_75t_L g15362 ( 
.A(n_14808),
.Y(n_15362)
);

INVxp67_ASAP7_75t_L g15363 ( 
.A(n_14614),
.Y(n_15363)
);

OAI21xp33_ASAP7_75t_L g15364 ( 
.A1(n_14320),
.A2(n_10946),
.B(n_10944),
.Y(n_15364)
);

INVx1_ASAP7_75t_L g15365 ( 
.A(n_14821),
.Y(n_15365)
);

INVx1_ASAP7_75t_L g15366 ( 
.A(n_14686),
.Y(n_15366)
);

AND2x4_ASAP7_75t_L g15367 ( 
.A(n_14547),
.B(n_8478),
.Y(n_15367)
);

NAND3xp33_ASAP7_75t_L g15368 ( 
.A(n_14407),
.B(n_11227),
.C(n_11156),
.Y(n_15368)
);

HB1xp67_ASAP7_75t_L g15369 ( 
.A(n_14834),
.Y(n_15369)
);

INVx1_ASAP7_75t_L g15370 ( 
.A(n_14690),
.Y(n_15370)
);

INVx1_ASAP7_75t_L g15371 ( 
.A(n_14393),
.Y(n_15371)
);

BUFx3_ASAP7_75t_L g15372 ( 
.A(n_14526),
.Y(n_15372)
);

AND2x4_ASAP7_75t_SL g15373 ( 
.A(n_14864),
.B(n_6907),
.Y(n_15373)
);

AND2x2_ASAP7_75t_L g15374 ( 
.A(n_14796),
.B(n_10944),
.Y(n_15374)
);

INVx2_ASAP7_75t_L g15375 ( 
.A(n_14550),
.Y(n_15375)
);

AND2x2_ASAP7_75t_L g15376 ( 
.A(n_14812),
.B(n_14817),
.Y(n_15376)
);

INVx2_ASAP7_75t_L g15377 ( 
.A(n_14677),
.Y(n_15377)
);

HB1xp67_ASAP7_75t_L g15378 ( 
.A(n_14834),
.Y(n_15378)
);

BUFx6f_ASAP7_75t_L g15379 ( 
.A(n_14502),
.Y(n_15379)
);

OAI221xp5_ASAP7_75t_SL g15380 ( 
.A1(n_14454),
.A2(n_9209),
.B1(n_9222),
.B2(n_9215),
.C(n_9189),
.Y(n_15380)
);

HB1xp67_ASAP7_75t_L g15381 ( 
.A(n_14835),
.Y(n_15381)
);

INVxp67_ASAP7_75t_SL g15382 ( 
.A(n_14746),
.Y(n_15382)
);

AND2x2_ASAP7_75t_L g15383 ( 
.A(n_14822),
.B(n_10946),
.Y(n_15383)
);

INVx1_ASAP7_75t_L g15384 ( 
.A(n_14410),
.Y(n_15384)
);

INVx1_ASAP7_75t_L g15385 ( 
.A(n_14806),
.Y(n_15385)
);

AOI22xp33_ASAP7_75t_L g15386 ( 
.A1(n_14361),
.A2(n_10228),
.B1(n_9994),
.B2(n_9753),
.Y(n_15386)
);

NAND2xp5_ASAP7_75t_L g15387 ( 
.A(n_14868),
.B(n_10950),
.Y(n_15387)
);

AND2x2_ASAP7_75t_L g15388 ( 
.A(n_14829),
.B(n_10950),
.Y(n_15388)
);

OR2x2_ASAP7_75t_L g15389 ( 
.A(n_14452),
.B(n_14470),
.Y(n_15389)
);

INVx1_ASAP7_75t_L g15390 ( 
.A(n_14416),
.Y(n_15390)
);

INVx2_ASAP7_75t_L g15391 ( 
.A(n_14681),
.Y(n_15391)
);

AND2x4_ASAP7_75t_L g15392 ( 
.A(n_14584),
.B(n_8478),
.Y(n_15392)
);

INVx1_ASAP7_75t_L g15393 ( 
.A(n_14427),
.Y(n_15393)
);

NAND2x1p5_ASAP7_75t_L g15394 ( 
.A(n_14875),
.B(n_8329),
.Y(n_15394)
);

AND2x2_ASAP7_75t_L g15395 ( 
.A(n_14839),
.B(n_10951),
.Y(n_15395)
);

OR2x2_ASAP7_75t_L g15396 ( 
.A(n_14396),
.B(n_10951),
.Y(n_15396)
);

AND2x2_ASAP7_75t_L g15397 ( 
.A(n_14842),
.B(n_10952),
.Y(n_15397)
);

AND2x2_ASAP7_75t_L g15398 ( 
.A(n_14846),
.B(n_10952),
.Y(n_15398)
);

INVx1_ASAP7_75t_L g15399 ( 
.A(n_14432),
.Y(n_15399)
);

AND2x2_ASAP7_75t_L g15400 ( 
.A(n_14848),
.B(n_10961),
.Y(n_15400)
);

OR2x2_ASAP7_75t_L g15401 ( 
.A(n_14599),
.B(n_10961),
.Y(n_15401)
);

INVx2_ASAP7_75t_L g15402 ( 
.A(n_14807),
.Y(n_15402)
);

AND2x2_ASAP7_75t_L g15403 ( 
.A(n_14851),
.B(n_10963),
.Y(n_15403)
);

OR2x2_ASAP7_75t_L g15404 ( 
.A(n_14549),
.B(n_10963),
.Y(n_15404)
);

NAND2xp5_ASAP7_75t_L g15405 ( 
.A(n_14622),
.B(n_10965),
.Y(n_15405)
);

HB1xp67_ASAP7_75t_L g15406 ( 
.A(n_14670),
.Y(n_15406)
);

NAND2xp5_ASAP7_75t_L g15407 ( 
.A(n_14465),
.B(n_10965),
.Y(n_15407)
);

INVxp67_ASAP7_75t_SL g15408 ( 
.A(n_14696),
.Y(n_15408)
);

INVx1_ASAP7_75t_L g15409 ( 
.A(n_14532),
.Y(n_15409)
);

AND2x2_ASAP7_75t_SL g15410 ( 
.A(n_14303),
.B(n_8923),
.Y(n_15410)
);

AND2x2_ASAP7_75t_L g15411 ( 
.A(n_14854),
.B(n_10979),
.Y(n_15411)
);

NAND3xp33_ASAP7_75t_L g15412 ( 
.A(n_14678),
.B(n_11227),
.C(n_11156),
.Y(n_15412)
);

AND2x2_ASAP7_75t_L g15413 ( 
.A(n_14866),
.B(n_14540),
.Y(n_15413)
);

INVx2_ASAP7_75t_L g15414 ( 
.A(n_14754),
.Y(n_15414)
);

INVx1_ASAP7_75t_L g15415 ( 
.A(n_14536),
.Y(n_15415)
);

INVx2_ASAP7_75t_L g15416 ( 
.A(n_14757),
.Y(n_15416)
);

AND2x2_ASAP7_75t_L g15417 ( 
.A(n_14512),
.B(n_10979),
.Y(n_15417)
);

INVx3_ASAP7_75t_L g15418 ( 
.A(n_14803),
.Y(n_15418)
);

OR2x2_ASAP7_75t_L g15419 ( 
.A(n_14287),
.B(n_10987),
.Y(n_15419)
);

INVx1_ASAP7_75t_L g15420 ( 
.A(n_14695),
.Y(n_15420)
);

INVx2_ASAP7_75t_L g15421 ( 
.A(n_14813),
.Y(n_15421)
);

NAND2x1_ASAP7_75t_L g15422 ( 
.A(n_14814),
.B(n_10517),
.Y(n_15422)
);

AND2x2_ASAP7_75t_L g15423 ( 
.A(n_14592),
.B(n_10987),
.Y(n_15423)
);

INVx1_ASAP7_75t_L g15424 ( 
.A(n_14662),
.Y(n_15424)
);

NAND2xp5_ASAP7_75t_L g15425 ( 
.A(n_14649),
.B(n_10988),
.Y(n_15425)
);

AND4x1_ASAP7_75t_L g15426 ( 
.A(n_14718),
.B(n_7402),
.C(n_7643),
.D(n_7589),
.Y(n_15426)
);

INVx1_ASAP7_75t_L g15427 ( 
.A(n_14398),
.Y(n_15427)
);

OR2x2_ASAP7_75t_L g15428 ( 
.A(n_14609),
.B(n_10988),
.Y(n_15428)
);

AND2x2_ASAP7_75t_L g15429 ( 
.A(n_14794),
.B(n_14853),
.Y(n_15429)
);

AND2x2_ASAP7_75t_L g15430 ( 
.A(n_14872),
.B(n_10989),
.Y(n_15430)
);

INVx1_ASAP7_75t_L g15431 ( 
.A(n_14377),
.Y(n_15431)
);

INVx1_ASAP7_75t_L g15432 ( 
.A(n_14385),
.Y(n_15432)
);

INVx2_ASAP7_75t_L g15433 ( 
.A(n_14798),
.Y(n_15433)
);

NAND2xp5_ASAP7_75t_SL g15434 ( 
.A(n_14756),
.B(n_8329),
.Y(n_15434)
);

INVx1_ASAP7_75t_L g15435 ( 
.A(n_14391),
.Y(n_15435)
);

INVxp67_ASAP7_75t_SL g15436 ( 
.A(n_14884),
.Y(n_15436)
);

NAND2xp5_ASAP7_75t_L g15437 ( 
.A(n_14656),
.B(n_10989),
.Y(n_15437)
);

OR2x2_ASAP7_75t_L g15438 ( 
.A(n_14543),
.B(n_10992),
.Y(n_15438)
);

NAND2xp5_ASAP7_75t_SL g15439 ( 
.A(n_14888),
.B(n_8340),
.Y(n_15439)
);

AND2x2_ASAP7_75t_L g15440 ( 
.A(n_14824),
.B(n_10992),
.Y(n_15440)
);

INVx2_ASAP7_75t_L g15441 ( 
.A(n_14841),
.Y(n_15441)
);

AND2x2_ASAP7_75t_L g15442 ( 
.A(n_14898),
.B(n_11002),
.Y(n_15442)
);

INVx2_ASAP7_75t_L g15443 ( 
.A(n_14823),
.Y(n_15443)
);

OR2x2_ASAP7_75t_L g15444 ( 
.A(n_14607),
.B(n_11002),
.Y(n_15444)
);

INVx1_ASAP7_75t_L g15445 ( 
.A(n_14402),
.Y(n_15445)
);

NAND2xp5_ASAP7_75t_L g15446 ( 
.A(n_14867),
.B(n_11005),
.Y(n_15446)
);

INVx1_ASAP7_75t_L g15447 ( 
.A(n_14414),
.Y(n_15447)
);

INVx1_ASAP7_75t_L g15448 ( 
.A(n_14444),
.Y(n_15448)
);

OR2x2_ASAP7_75t_L g15449 ( 
.A(n_14415),
.B(n_11005),
.Y(n_15449)
);

INVx1_ASAP7_75t_L g15450 ( 
.A(n_14450),
.Y(n_15450)
);

AND2x2_ASAP7_75t_L g15451 ( 
.A(n_14899),
.B(n_11013),
.Y(n_15451)
);

HB1xp67_ASAP7_75t_L g15452 ( 
.A(n_14767),
.Y(n_15452)
);

NAND2xp5_ASAP7_75t_L g15453 ( 
.A(n_14880),
.B(n_11013),
.Y(n_15453)
);

INVxp67_ASAP7_75t_SL g15454 ( 
.A(n_14628),
.Y(n_15454)
);

HB1xp67_ASAP7_75t_L g15455 ( 
.A(n_14869),
.Y(n_15455)
);

INVx2_ASAP7_75t_L g15456 ( 
.A(n_14878),
.Y(n_15456)
);

OR2x2_ASAP7_75t_L g15457 ( 
.A(n_14727),
.B(n_14889),
.Y(n_15457)
);

INVx1_ASAP7_75t_L g15458 ( 
.A(n_14440),
.Y(n_15458)
);

INVx1_ASAP7_75t_SL g15459 ( 
.A(n_14633),
.Y(n_15459)
);

NAND2xp5_ASAP7_75t_L g15460 ( 
.A(n_14760),
.B(n_11014),
.Y(n_15460)
);

INVx1_ASAP7_75t_L g15461 ( 
.A(n_14441),
.Y(n_15461)
);

AND2x4_ASAP7_75t_L g15462 ( 
.A(n_14818),
.B(n_8478),
.Y(n_15462)
);

INVxp67_ASAP7_75t_L g15463 ( 
.A(n_14845),
.Y(n_15463)
);

OR2x2_ASAP7_75t_L g15464 ( 
.A(n_14635),
.B(n_11014),
.Y(n_15464)
);

OR2x2_ASAP7_75t_L g15465 ( 
.A(n_14641),
.B(n_11032),
.Y(n_15465)
);

NAND2xp5_ASAP7_75t_L g15466 ( 
.A(n_14820),
.B(n_11032),
.Y(n_15466)
);

AND2x2_ASAP7_75t_L g15467 ( 
.A(n_14893),
.B(n_11034),
.Y(n_15467)
);

NAND2xp5_ASAP7_75t_L g15468 ( 
.A(n_14901),
.B(n_11034),
.Y(n_15468)
);

AND2x2_ASAP7_75t_L g15469 ( 
.A(n_14838),
.B(n_11040),
.Y(n_15469)
);

AND2x2_ASAP7_75t_L g15470 ( 
.A(n_14840),
.B(n_11040),
.Y(n_15470)
);

INVx1_ASAP7_75t_L g15471 ( 
.A(n_14453),
.Y(n_15471)
);

INVx1_ASAP7_75t_L g15472 ( 
.A(n_14455),
.Y(n_15472)
);

INVx2_ASAP7_75t_L g15473 ( 
.A(n_14778),
.Y(n_15473)
);

AND2x2_ASAP7_75t_L g15474 ( 
.A(n_14825),
.B(n_14827),
.Y(n_15474)
);

OR2x2_ASAP7_75t_L g15475 ( 
.A(n_14702),
.B(n_11042),
.Y(n_15475)
);

AND2x2_ASAP7_75t_L g15476 ( 
.A(n_14830),
.B(n_14903),
.Y(n_15476)
);

AND2x4_ASAP7_75t_L g15477 ( 
.A(n_14460),
.B(n_14461),
.Y(n_15477)
);

INVx2_ASAP7_75t_L g15478 ( 
.A(n_14900),
.Y(n_15478)
);

AND2x2_ASAP7_75t_L g15479 ( 
.A(n_14904),
.B(n_11042),
.Y(n_15479)
);

INVx1_ASAP7_75t_L g15480 ( 
.A(n_14466),
.Y(n_15480)
);

AND2x2_ASAP7_75t_L g15481 ( 
.A(n_14892),
.B(n_11044),
.Y(n_15481)
);

INVx1_ASAP7_75t_L g15482 ( 
.A(n_14477),
.Y(n_15482)
);

BUFx2_ASAP7_75t_L g15483 ( 
.A(n_14716),
.Y(n_15483)
);

AND2x2_ASAP7_75t_L g15484 ( 
.A(n_14881),
.B(n_14906),
.Y(n_15484)
);

INVx1_ASAP7_75t_L g15485 ( 
.A(n_14478),
.Y(n_15485)
);

OR2x2_ASAP7_75t_L g15486 ( 
.A(n_14759),
.B(n_11044),
.Y(n_15486)
);

NAND2xp5_ASAP7_75t_L g15487 ( 
.A(n_14849),
.B(n_11045),
.Y(n_15487)
);

NAND2xp5_ASAP7_75t_L g15488 ( 
.A(n_14850),
.B(n_11045),
.Y(n_15488)
);

OR2x2_ASAP7_75t_L g15489 ( 
.A(n_14786),
.B(n_14863),
.Y(n_15489)
);

INVx1_ASAP7_75t_L g15490 ( 
.A(n_14480),
.Y(n_15490)
);

NAND2xp5_ASAP7_75t_L g15491 ( 
.A(n_14857),
.B(n_11046),
.Y(n_15491)
);

NAND2x1_ASAP7_75t_L g15492 ( 
.A(n_14814),
.B(n_10517),
.Y(n_15492)
);

AND2x2_ASAP7_75t_L g15493 ( 
.A(n_14764),
.B(n_11046),
.Y(n_15493)
);

NAND2xp5_ASAP7_75t_L g15494 ( 
.A(n_14861),
.B(n_11047),
.Y(n_15494)
);

INVx1_ASAP7_75t_L g15495 ( 
.A(n_14483),
.Y(n_15495)
);

INVx1_ASAP7_75t_SL g15496 ( 
.A(n_14782),
.Y(n_15496)
);

INVx2_ASAP7_75t_L g15497 ( 
.A(n_14793),
.Y(n_15497)
);

AND2x2_ASAP7_75t_L g15498 ( 
.A(n_14769),
.B(n_11047),
.Y(n_15498)
);

INVx2_ASAP7_75t_L g15499 ( 
.A(n_14797),
.Y(n_15499)
);

AND2x2_ASAP7_75t_L g15500 ( 
.A(n_14770),
.B(n_11050),
.Y(n_15500)
);

AND2x2_ASAP7_75t_L g15501 ( 
.A(n_14777),
.B(n_11050),
.Y(n_15501)
);

AND2x2_ASAP7_75t_L g15502 ( 
.A(n_14779),
.B(n_11052),
.Y(n_15502)
);

AND2x4_ASAP7_75t_L g15503 ( 
.A(n_14484),
.B(n_8478),
.Y(n_15503)
);

AND2x2_ASAP7_75t_L g15504 ( 
.A(n_14858),
.B(n_11052),
.Y(n_15504)
);

INVx1_ASAP7_75t_L g15505 ( 
.A(n_14491),
.Y(n_15505)
);

INVx1_ASAP7_75t_L g15506 ( 
.A(n_14507),
.Y(n_15506)
);

NAND2xp5_ASAP7_75t_L g15507 ( 
.A(n_14871),
.B(n_11056),
.Y(n_15507)
);

INVx1_ASAP7_75t_L g15508 ( 
.A(n_14510),
.Y(n_15508)
);

INVx2_ASAP7_75t_L g15509 ( 
.A(n_14800),
.Y(n_15509)
);

INVx1_ASAP7_75t_SL g15510 ( 
.A(n_14879),
.Y(n_15510)
);

AND2x2_ASAP7_75t_L g15511 ( 
.A(n_14768),
.B(n_11056),
.Y(n_15511)
);

AND2x4_ASAP7_75t_L g15512 ( 
.A(n_14519),
.B(n_14523),
.Y(n_15512)
);

INVx1_ASAP7_75t_L g15513 ( 
.A(n_14524),
.Y(n_15513)
);

AND2x2_ASAP7_75t_L g15514 ( 
.A(n_14865),
.B(n_11059),
.Y(n_15514)
);

NAND2xp5_ASAP7_75t_L g15515 ( 
.A(n_14873),
.B(n_11059),
.Y(n_15515)
);

AND2x2_ASAP7_75t_L g15516 ( 
.A(n_14885),
.B(n_11064),
.Y(n_15516)
);

INVx1_ASAP7_75t_L g15517 ( 
.A(n_14434),
.Y(n_15517)
);

INVx2_ASAP7_75t_L g15518 ( 
.A(n_14804),
.Y(n_15518)
);

INVx1_ASAP7_75t_L g15519 ( 
.A(n_14436),
.Y(n_15519)
);

AND2x4_ASAP7_75t_SL g15520 ( 
.A(n_14891),
.B(n_6907),
.Y(n_15520)
);

INVx1_ASAP7_75t_L g15521 ( 
.A(n_14439),
.Y(n_15521)
);

INVx2_ASAP7_75t_L g15522 ( 
.A(n_14785),
.Y(n_15522)
);

INVx1_ASAP7_75t_L g15523 ( 
.A(n_15483),
.Y(n_15523)
);

AND2x4_ASAP7_75t_L g15524 ( 
.A(n_14980),
.B(n_14936),
.Y(n_15524)
);

AND2x2_ASAP7_75t_L g15525 ( 
.A(n_14921),
.B(n_14445),
.Y(n_15525)
);

OR2x2_ASAP7_75t_L g15526 ( 
.A(n_15012),
.B(n_14860),
.Y(n_15526)
);

INVx1_ASAP7_75t_L g15527 ( 
.A(n_15483),
.Y(n_15527)
);

AND2x2_ASAP7_75t_L g15528 ( 
.A(n_14966),
.B(n_14832),
.Y(n_15528)
);

NAND2xp5_ASAP7_75t_L g15529 ( 
.A(n_14941),
.B(n_14538),
.Y(n_15529)
);

NAND2xp5_ASAP7_75t_L g15530 ( 
.A(n_15090),
.B(n_14551),
.Y(n_15530)
);

NAND2xp5_ASAP7_75t_L g15531 ( 
.A(n_14907),
.B(n_14552),
.Y(n_15531)
);

NAND2xp5_ASAP7_75t_L g15532 ( 
.A(n_14989),
.B(n_14558),
.Y(n_15532)
);

HB1xp67_ASAP7_75t_L g15533 ( 
.A(n_14984),
.Y(n_15533)
);

INVx2_ASAP7_75t_L g15534 ( 
.A(n_14950),
.Y(n_15534)
);

AND2x2_ASAP7_75t_L g15535 ( 
.A(n_14924),
.B(n_14856),
.Y(n_15535)
);

AND2x2_ASAP7_75t_L g15536 ( 
.A(n_14938),
.B(n_15099),
.Y(n_15536)
);

NOR2xp33_ASAP7_75t_L g15537 ( 
.A(n_15229),
.B(n_15243),
.Y(n_15537)
);

OR2x2_ASAP7_75t_L g15538 ( 
.A(n_14961),
.B(n_14833),
.Y(n_15538)
);

AND2x2_ASAP7_75t_L g15539 ( 
.A(n_15089),
.B(n_14852),
.Y(n_15539)
);

INVx1_ASAP7_75t_L g15540 ( 
.A(n_14937),
.Y(n_15540)
);

INVx2_ASAP7_75t_L g15541 ( 
.A(n_14995),
.Y(n_15541)
);

AND2x4_ASAP7_75t_L g15542 ( 
.A(n_15064),
.B(n_14563),
.Y(n_15542)
);

NOR2xp33_ASAP7_75t_L g15543 ( 
.A(n_15101),
.B(n_14475),
.Y(n_15543)
);

OAI33xp33_ASAP7_75t_L g15544 ( 
.A1(n_15420),
.A2(n_14578),
.A3(n_14571),
.B1(n_14579),
.B2(n_14572),
.B3(n_14566),
.Y(n_15544)
);

INVx2_ASAP7_75t_L g15545 ( 
.A(n_15042),
.Y(n_15545)
);

AND2x2_ASAP7_75t_L g15546 ( 
.A(n_15080),
.B(n_14581),
.Y(n_15546)
);

INVx1_ASAP7_75t_L g15547 ( 
.A(n_14946),
.Y(n_15547)
);

AND2x2_ASAP7_75t_L g15548 ( 
.A(n_15238),
.B(n_14582),
.Y(n_15548)
);

AND2x4_ASAP7_75t_L g15549 ( 
.A(n_14934),
.B(n_14583),
.Y(n_15549)
);

NAND2xp5_ASAP7_75t_L g15550 ( 
.A(n_15408),
.B(n_14586),
.Y(n_15550)
);

OAI21xp33_ASAP7_75t_L g15551 ( 
.A1(n_15282),
.A2(n_14802),
.B(n_14801),
.Y(n_15551)
);

INVx1_ASAP7_75t_L g15552 ( 
.A(n_15350),
.Y(n_15552)
);

INVx2_ASAP7_75t_L g15553 ( 
.A(n_15350),
.Y(n_15553)
);

NAND2x1_ASAP7_75t_L g15554 ( 
.A(n_14919),
.B(n_14590),
.Y(n_15554)
);

AND2x2_ASAP7_75t_L g15555 ( 
.A(n_15247),
.B(n_14591),
.Y(n_15555)
);

OR2x2_ASAP7_75t_L g15556 ( 
.A(n_14970),
.B(n_14896),
.Y(n_15556)
);

NOR2xp33_ASAP7_75t_L g15557 ( 
.A(n_15271),
.B(n_14595),
.Y(n_15557)
);

AND2x2_ASAP7_75t_L g15558 ( 
.A(n_15112),
.B(n_14600),
.Y(n_15558)
);

AND2x2_ASAP7_75t_L g15559 ( 
.A(n_15162),
.B(n_15185),
.Y(n_15559)
);

AND2x2_ASAP7_75t_L g15560 ( 
.A(n_15267),
.B(n_14601),
.Y(n_15560)
);

INVxp67_ASAP7_75t_L g15561 ( 
.A(n_15318),
.Y(n_15561)
);

AND2x2_ASAP7_75t_L g15562 ( 
.A(n_14910),
.B(n_14602),
.Y(n_15562)
);

INVx1_ASAP7_75t_L g15563 ( 
.A(n_15197),
.Y(n_15563)
);

OR2x2_ASAP7_75t_L g15564 ( 
.A(n_14986),
.B(n_14772),
.Y(n_15564)
);

AND2x2_ASAP7_75t_L g15565 ( 
.A(n_15038),
.B(n_14604),
.Y(n_15565)
);

BUFx3_ASAP7_75t_L g15566 ( 
.A(n_15278),
.Y(n_15566)
);

INVx2_ASAP7_75t_L g15567 ( 
.A(n_14913),
.Y(n_15567)
);

AND2x2_ASAP7_75t_L g15568 ( 
.A(n_15045),
.B(n_14611),
.Y(n_15568)
);

INVx1_ASAP7_75t_L g15569 ( 
.A(n_15347),
.Y(n_15569)
);

INVx1_ASAP7_75t_L g15570 ( 
.A(n_15369),
.Y(n_15570)
);

INVxp33_ASAP7_75t_L g15571 ( 
.A(n_15273),
.Y(n_15571)
);

AND2x2_ASAP7_75t_L g15572 ( 
.A(n_15057),
.B(n_14613),
.Y(n_15572)
);

INVx2_ASAP7_75t_L g15573 ( 
.A(n_14930),
.Y(n_15573)
);

INVx2_ASAP7_75t_L g15574 ( 
.A(n_15209),
.Y(n_15574)
);

OR2x2_ASAP7_75t_L g15575 ( 
.A(n_14987),
.B(n_14837),
.Y(n_15575)
);

HB1xp67_ASAP7_75t_L g15576 ( 
.A(n_14919),
.Y(n_15576)
);

INVx2_ASAP7_75t_L g15577 ( 
.A(n_15209),
.Y(n_15577)
);

INVx1_ASAP7_75t_L g15578 ( 
.A(n_15378),
.Y(n_15578)
);

OR2x2_ASAP7_75t_L g15579 ( 
.A(n_15301),
.B(n_14959),
.Y(n_15579)
);

AND2x2_ASAP7_75t_L g15580 ( 
.A(n_15164),
.B(n_14617),
.Y(n_15580)
);

INVx1_ASAP7_75t_L g15581 ( 
.A(n_14908),
.Y(n_15581)
);

INVx2_ASAP7_75t_SL g15582 ( 
.A(n_15003),
.Y(n_15582)
);

AND2x4_ASAP7_75t_L g15583 ( 
.A(n_15046),
.B(n_14619),
.Y(n_15583)
);

INVx1_ASAP7_75t_L g15584 ( 
.A(n_14909),
.Y(n_15584)
);

AND2x2_ASAP7_75t_L g15585 ( 
.A(n_14991),
.B(n_15048),
.Y(n_15585)
);

INVx1_ASAP7_75t_L g15586 ( 
.A(n_14928),
.Y(n_15586)
);

AND2x2_ASAP7_75t_L g15587 ( 
.A(n_15312),
.B(n_14620),
.Y(n_15587)
);

INVx2_ASAP7_75t_L g15588 ( 
.A(n_14948),
.Y(n_15588)
);

NOR4xp25_ASAP7_75t_SL g15589 ( 
.A(n_15136),
.B(n_14646),
.C(n_14651),
.D(n_14634),
.Y(n_15589)
);

AND2x2_ASAP7_75t_L g15590 ( 
.A(n_14965),
.B(n_14973),
.Y(n_15590)
);

AND2x2_ASAP7_75t_L g15591 ( 
.A(n_15098),
.B(n_14652),
.Y(n_15591)
);

INVx2_ASAP7_75t_L g15592 ( 
.A(n_14951),
.Y(n_15592)
);

INVx1_ASAP7_75t_L g15593 ( 
.A(n_14935),
.Y(n_15593)
);

INVx2_ASAP7_75t_L g15594 ( 
.A(n_15262),
.Y(n_15594)
);

INVx3_ASAP7_75t_L g15595 ( 
.A(n_14912),
.Y(n_15595)
);

OR2x2_ASAP7_75t_L g15596 ( 
.A(n_15145),
.B(n_14859),
.Y(n_15596)
);

AND2x2_ASAP7_75t_L g15597 ( 
.A(n_15108),
.B(n_14660),
.Y(n_15597)
);

OR2x2_ASAP7_75t_L g15598 ( 
.A(n_14960),
.B(n_14664),
.Y(n_15598)
);

BUFx2_ASAP7_75t_L g15599 ( 
.A(n_15136),
.Y(n_15599)
);

INVx1_ASAP7_75t_L g15600 ( 
.A(n_15072),
.Y(n_15600)
);

NAND2xp5_ASAP7_75t_L g15601 ( 
.A(n_15222),
.B(n_14668),
.Y(n_15601)
);

INVx2_ASAP7_75t_L g15602 ( 
.A(n_14947),
.Y(n_15602)
);

INVx2_ASAP7_75t_L g15603 ( 
.A(n_15008),
.Y(n_15603)
);

NAND2xp5_ASAP7_75t_L g15604 ( 
.A(n_15246),
.B(n_14672),
.Y(n_15604)
);

NAND2xp5_ASAP7_75t_L g15605 ( 
.A(n_14967),
.B(n_14674),
.Y(n_15605)
);

INVx1_ASAP7_75t_L g15606 ( 
.A(n_15074),
.Y(n_15606)
);

AND2x2_ASAP7_75t_L g15607 ( 
.A(n_15110),
.B(n_14684),
.Y(n_15607)
);

INVx1_ASAP7_75t_L g15608 ( 
.A(n_15452),
.Y(n_15608)
);

AND2x2_ASAP7_75t_L g15609 ( 
.A(n_15119),
.B(n_14694),
.Y(n_15609)
);

AND2x4_ASAP7_75t_L g15610 ( 
.A(n_15173),
.B(n_14705),
.Y(n_15610)
);

AND2x2_ASAP7_75t_L g15611 ( 
.A(n_14917),
.B(n_14722),
.Y(n_15611)
);

OR2x2_ASAP7_75t_L g15612 ( 
.A(n_14964),
.B(n_14728),
.Y(n_15612)
);

OR2x2_ASAP7_75t_L g15613 ( 
.A(n_15316),
.B(n_14730),
.Y(n_15613)
);

AND2x4_ASAP7_75t_SL g15614 ( 
.A(n_15429),
.B(n_14735),
.Y(n_15614)
);

INVx2_ASAP7_75t_L g15615 ( 
.A(n_15053),
.Y(n_15615)
);

INVx1_ASAP7_75t_L g15616 ( 
.A(n_15117),
.Y(n_15616)
);

NAND2xp5_ASAP7_75t_L g15617 ( 
.A(n_15203),
.B(n_14740),
.Y(n_15617)
);

AND2x2_ASAP7_75t_L g15618 ( 
.A(n_14911),
.B(n_14741),
.Y(n_15618)
);

INVx2_ASAP7_75t_L g15619 ( 
.A(n_15002),
.Y(n_15619)
);

NOR2xp33_ASAP7_75t_L g15620 ( 
.A(n_15379),
.B(n_14742),
.Y(n_15620)
);

HB1xp67_ASAP7_75t_L g15621 ( 
.A(n_15157),
.Y(n_15621)
);

NAND2xp5_ASAP7_75t_L g15622 ( 
.A(n_15211),
.B(n_14743),
.Y(n_15622)
);

NAND2xp5_ASAP7_75t_L g15623 ( 
.A(n_14939),
.B(n_14744),
.Y(n_15623)
);

INVx1_ASAP7_75t_L g15624 ( 
.A(n_15044),
.Y(n_15624)
);

INVx2_ASAP7_75t_L g15625 ( 
.A(n_15059),
.Y(n_15625)
);

AND2x2_ASAP7_75t_L g15626 ( 
.A(n_15147),
.B(n_14762),
.Y(n_15626)
);

NAND2xp5_ASAP7_75t_L g15627 ( 
.A(n_14943),
.B(n_14774),
.Y(n_15627)
);

INVx1_ASAP7_75t_SL g15628 ( 
.A(n_14915),
.Y(n_15628)
);

AND2x2_ASAP7_75t_L g15629 ( 
.A(n_15050),
.B(n_14781),
.Y(n_15629)
);

AND2x2_ASAP7_75t_L g15630 ( 
.A(n_14985),
.B(n_14974),
.Y(n_15630)
);

AND2x2_ASAP7_75t_L g15631 ( 
.A(n_14978),
.B(n_14870),
.Y(n_15631)
);

NAND2xp5_ASAP7_75t_L g15632 ( 
.A(n_14945),
.B(n_14810),
.Y(n_15632)
);

INVx1_ASAP7_75t_L g15633 ( 
.A(n_15047),
.Y(n_15633)
);

AND2x2_ASAP7_75t_L g15634 ( 
.A(n_15290),
.B(n_14887),
.Y(n_15634)
);

NAND2xp5_ASAP7_75t_L g15635 ( 
.A(n_14953),
.B(n_14962),
.Y(n_15635)
);

AND2x2_ASAP7_75t_L g15636 ( 
.A(n_15067),
.B(n_14816),
.Y(n_15636)
);

OR2x2_ASAP7_75t_L g15637 ( 
.A(n_15196),
.B(n_14905),
.Y(n_15637)
);

AND2x2_ASAP7_75t_L g15638 ( 
.A(n_14957),
.B(n_11064),
.Y(n_15638)
);

AND2x4_ASAP7_75t_L g15639 ( 
.A(n_14968),
.B(n_8478),
.Y(n_15639)
);

NAND2x1p5_ASAP7_75t_L g15640 ( 
.A(n_15084),
.B(n_8340),
.Y(n_15640)
);

OR2x2_ASAP7_75t_L g15641 ( 
.A(n_15321),
.B(n_14890),
.Y(n_15641)
);

NAND2xp5_ASAP7_75t_L g15642 ( 
.A(n_15187),
.B(n_11087),
.Y(n_15642)
);

AND2x4_ASAP7_75t_L g15643 ( 
.A(n_15351),
.B(n_8479),
.Y(n_15643)
);

AND2x2_ASAP7_75t_L g15644 ( 
.A(n_14998),
.B(n_11087),
.Y(n_15644)
);

AOI221xp5_ASAP7_75t_L g15645 ( 
.A1(n_14922),
.A2(n_9222),
.B1(n_9237),
.B2(n_9215),
.C(n_9209),
.Y(n_15645)
);

INVx1_ASAP7_75t_L g15646 ( 
.A(n_15051),
.Y(n_15646)
);

INVx1_ASAP7_75t_L g15647 ( 
.A(n_15058),
.Y(n_15647)
);

INVx1_ASAP7_75t_SL g15648 ( 
.A(n_14954),
.Y(n_15648)
);

INVx1_ASAP7_75t_L g15649 ( 
.A(n_15069),
.Y(n_15649)
);

INVx2_ASAP7_75t_L g15650 ( 
.A(n_15009),
.Y(n_15650)
);

AND2x2_ASAP7_75t_L g15651 ( 
.A(n_15018),
.B(n_11090),
.Y(n_15651)
);

BUFx3_ASAP7_75t_L g15652 ( 
.A(n_15029),
.Y(n_15652)
);

AND2x2_ASAP7_75t_L g15653 ( 
.A(n_15026),
.B(n_11090),
.Y(n_15653)
);

INVx1_ASAP7_75t_L g15654 ( 
.A(n_14916),
.Y(n_15654)
);

INVx1_ASAP7_75t_L g15655 ( 
.A(n_15427),
.Y(n_15655)
);

INVx4_ASAP7_75t_L g15656 ( 
.A(n_15289),
.Y(n_15656)
);

INVx2_ASAP7_75t_L g15657 ( 
.A(n_15024),
.Y(n_15657)
);

INVx1_ASAP7_75t_L g15658 ( 
.A(n_15176),
.Y(n_15658)
);

OR2x2_ASAP7_75t_L g15659 ( 
.A(n_15081),
.B(n_11094),
.Y(n_15659)
);

INVx2_ASAP7_75t_L g15660 ( 
.A(n_15078),
.Y(n_15660)
);

AND2x4_ASAP7_75t_L g15661 ( 
.A(n_15177),
.B(n_8479),
.Y(n_15661)
);

INVx1_ASAP7_75t_L g15662 ( 
.A(n_15183),
.Y(n_15662)
);

INVx2_ASAP7_75t_L g15663 ( 
.A(n_15131),
.Y(n_15663)
);

AND2x2_ASAP7_75t_L g15664 ( 
.A(n_15043),
.B(n_11094),
.Y(n_15664)
);

BUFx3_ASAP7_75t_L g15665 ( 
.A(n_14912),
.Y(n_15665)
);

NOR2xp33_ASAP7_75t_L g15666 ( 
.A(n_15379),
.B(n_11100),
.Y(n_15666)
);

OR2x2_ASAP7_75t_L g15667 ( 
.A(n_15151),
.B(n_11100),
.Y(n_15667)
);

INVx1_ASAP7_75t_L g15668 ( 
.A(n_15138),
.Y(n_15668)
);

AND2x4_ASAP7_75t_L g15669 ( 
.A(n_15178),
.B(n_8479),
.Y(n_15669)
);

AND2x2_ASAP7_75t_L g15670 ( 
.A(n_15075),
.B(n_11101),
.Y(n_15670)
);

INVx6_ASAP7_75t_L g15671 ( 
.A(n_15010),
.Y(n_15671)
);

NAND2xp5_ASAP7_75t_L g15672 ( 
.A(n_15189),
.B(n_11101),
.Y(n_15672)
);

NAND2xp5_ASAP7_75t_L g15673 ( 
.A(n_15190),
.B(n_11108),
.Y(n_15673)
);

INVx1_ASAP7_75t_L g15674 ( 
.A(n_15455),
.Y(n_15674)
);

AND2x2_ASAP7_75t_L g15675 ( 
.A(n_15095),
.B(n_11108),
.Y(n_15675)
);

OAI31xp33_ASAP7_75t_L g15676 ( 
.A1(n_15381),
.A2(n_9237),
.A3(n_9256),
.B(n_9222),
.Y(n_15676)
);

INVx1_ASAP7_75t_L g15677 ( 
.A(n_14926),
.Y(n_15677)
);

AND2x2_ASAP7_75t_L g15678 ( 
.A(n_14975),
.B(n_11109),
.Y(n_15678)
);

NAND2xp5_ASAP7_75t_L g15679 ( 
.A(n_14979),
.B(n_11109),
.Y(n_15679)
);

AND2x2_ASAP7_75t_L g15680 ( 
.A(n_15184),
.B(n_11119),
.Y(n_15680)
);

INVx2_ASAP7_75t_L g15681 ( 
.A(n_15071),
.Y(n_15681)
);

AND2x2_ASAP7_75t_L g15682 ( 
.A(n_15200),
.B(n_11119),
.Y(n_15682)
);

INVx1_ASAP7_75t_L g15683 ( 
.A(n_14933),
.Y(n_15683)
);

AND2x2_ASAP7_75t_L g15684 ( 
.A(n_15202),
.B(n_11130),
.Y(n_15684)
);

AND2x2_ASAP7_75t_L g15685 ( 
.A(n_15023),
.B(n_11130),
.Y(n_15685)
);

INVx1_ASAP7_75t_L g15686 ( 
.A(n_14927),
.Y(n_15686)
);

AOI22xp33_ASAP7_75t_L g15687 ( 
.A1(n_15028),
.A2(n_10228),
.B1(n_11227),
.B2(n_11156),
.Y(n_15687)
);

HB1xp67_ASAP7_75t_L g15688 ( 
.A(n_15034),
.Y(n_15688)
);

AND2x4_ASAP7_75t_L g15689 ( 
.A(n_15134),
.B(n_8479),
.Y(n_15689)
);

AND2x2_ASAP7_75t_L g15690 ( 
.A(n_15302),
.B(n_11131),
.Y(n_15690)
);

NAND2x1p5_ASAP7_75t_L g15691 ( 
.A(n_14929),
.B(n_8340),
.Y(n_15691)
);

INVx2_ASAP7_75t_L g15692 ( 
.A(n_15154),
.Y(n_15692)
);

NAND2xp67_ASAP7_75t_L g15693 ( 
.A(n_15255),
.B(n_11131),
.Y(n_15693)
);

INVxp67_ASAP7_75t_L g15694 ( 
.A(n_15260),
.Y(n_15694)
);

AND2x2_ASAP7_75t_L g15695 ( 
.A(n_15040),
.B(n_11133),
.Y(n_15695)
);

INVxp67_ASAP7_75t_L g15696 ( 
.A(n_14993),
.Y(n_15696)
);

AND2x2_ASAP7_75t_L g15697 ( 
.A(n_15020),
.B(n_11133),
.Y(n_15697)
);

AND2x2_ASAP7_75t_L g15698 ( 
.A(n_15413),
.B(n_11137),
.Y(n_15698)
);

AND2x2_ASAP7_75t_L g15699 ( 
.A(n_15402),
.B(n_11137),
.Y(n_15699)
);

OR2x2_ASAP7_75t_L g15700 ( 
.A(n_14981),
.B(n_14914),
.Y(n_15700)
);

NAND2xp5_ASAP7_75t_L g15701 ( 
.A(n_15077),
.B(n_15169),
.Y(n_15701)
);

AND2x2_ASAP7_75t_L g15702 ( 
.A(n_15416),
.B(n_11148),
.Y(n_15702)
);

INVx2_ASAP7_75t_SL g15703 ( 
.A(n_15076),
.Y(n_15703)
);

NAND2xp5_ASAP7_75t_L g15704 ( 
.A(n_15175),
.B(n_11148),
.Y(n_15704)
);

INVx1_ASAP7_75t_L g15705 ( 
.A(n_14977),
.Y(n_15705)
);

INVx1_ASAP7_75t_SL g15706 ( 
.A(n_15052),
.Y(n_15706)
);

INVx2_ASAP7_75t_L g15707 ( 
.A(n_15124),
.Y(n_15707)
);

HB1xp67_ASAP7_75t_L g15708 ( 
.A(n_15126),
.Y(n_15708)
);

BUFx2_ASAP7_75t_L g15709 ( 
.A(n_15148),
.Y(n_15709)
);

OR2x2_ASAP7_75t_L g15710 ( 
.A(n_15035),
.B(n_11149),
.Y(n_15710)
);

AND2x4_ASAP7_75t_L g15711 ( 
.A(n_15377),
.B(n_8479),
.Y(n_15711)
);

AND2x2_ASAP7_75t_L g15712 ( 
.A(n_15308),
.B(n_11149),
.Y(n_15712)
);

INVx2_ASAP7_75t_L g15713 ( 
.A(n_15303),
.Y(n_15713)
);

AND2x2_ASAP7_75t_L g15714 ( 
.A(n_15376),
.B(n_11151),
.Y(n_15714)
);

AND2x2_ASAP7_75t_L g15715 ( 
.A(n_14956),
.B(n_11151),
.Y(n_15715)
);

OR2x2_ASAP7_75t_L g15716 ( 
.A(n_14923),
.B(n_11161),
.Y(n_15716)
);

AOI22xp33_ASAP7_75t_L g15717 ( 
.A1(n_14969),
.A2(n_11267),
.B1(n_9994),
.B2(n_9753),
.Y(n_15717)
);

OR2x2_ASAP7_75t_L g15718 ( 
.A(n_15021),
.B(n_11161),
.Y(n_15718)
);

INVx1_ASAP7_75t_L g15719 ( 
.A(n_15005),
.Y(n_15719)
);

AND2x4_ASAP7_75t_L g15720 ( 
.A(n_15391),
.B(n_8528),
.Y(n_15720)
);

AND2x2_ASAP7_75t_L g15721 ( 
.A(n_15314),
.B(n_11164),
.Y(n_15721)
);

INVx2_ASAP7_75t_SL g15722 ( 
.A(n_15022),
.Y(n_15722)
);

OR2x2_ASAP7_75t_L g15723 ( 
.A(n_15342),
.B(n_11164),
.Y(n_15723)
);

INVx1_ASAP7_75t_L g15724 ( 
.A(n_15001),
.Y(n_15724)
);

OAI22xp5_ASAP7_75t_L g15725 ( 
.A1(n_15073),
.A2(n_10517),
.B1(n_11365),
.B2(n_7870),
.Y(n_15725)
);

NOR2x1_ASAP7_75t_L g15726 ( 
.A(n_15011),
.B(n_15106),
.Y(n_15726)
);

INVx1_ASAP7_75t_L g15727 ( 
.A(n_15127),
.Y(n_15727)
);

NAND2xp5_ASAP7_75t_L g15728 ( 
.A(n_15079),
.B(n_11167),
.Y(n_15728)
);

NAND2xp5_ASAP7_75t_L g15729 ( 
.A(n_15292),
.B(n_11167),
.Y(n_15729)
);

INVx1_ASAP7_75t_L g15730 ( 
.A(n_15165),
.Y(n_15730)
);

NAND2xp5_ASAP7_75t_L g15731 ( 
.A(n_15295),
.B(n_11168),
.Y(n_15731)
);

OR2x6_ASAP7_75t_L g15732 ( 
.A(n_14972),
.B(n_15210),
.Y(n_15732)
);

HB1xp67_ASAP7_75t_L g15733 ( 
.A(n_15329),
.Y(n_15733)
);

INVx2_ASAP7_75t_SL g15734 ( 
.A(n_14994),
.Y(n_15734)
);

INVx2_ASAP7_75t_L g15735 ( 
.A(n_15208),
.Y(n_15735)
);

INVx1_ASAP7_75t_L g15736 ( 
.A(n_14996),
.Y(n_15736)
);

NAND2xp33_ASAP7_75t_R g15737 ( 
.A(n_15000),
.B(n_7182),
.Y(n_15737)
);

AND2x2_ASAP7_75t_L g15738 ( 
.A(n_15459),
.B(n_11168),
.Y(n_15738)
);

AND2x2_ASAP7_75t_L g15739 ( 
.A(n_15037),
.B(n_11171),
.Y(n_15739)
);

AND2x2_ASAP7_75t_L g15740 ( 
.A(n_15418),
.B(n_11171),
.Y(n_15740)
);

AND2x4_ASAP7_75t_L g15741 ( 
.A(n_15226),
.B(n_8528),
.Y(n_15741)
);

INVx1_ASAP7_75t_L g15742 ( 
.A(n_15115),
.Y(n_15742)
);

INVxp67_ASAP7_75t_SL g15743 ( 
.A(n_15068),
.Y(n_15743)
);

INVx2_ASAP7_75t_L g15744 ( 
.A(n_15215),
.Y(n_15744)
);

AND2x2_ASAP7_75t_L g15745 ( 
.A(n_15054),
.B(n_11180),
.Y(n_15745)
);

AND2x2_ASAP7_75t_L g15746 ( 
.A(n_15424),
.B(n_15341),
.Y(n_15746)
);

AND2x2_ASAP7_75t_L g15747 ( 
.A(n_15228),
.B(n_11180),
.Y(n_15747)
);

NOR2xp33_ASAP7_75t_L g15748 ( 
.A(n_15363),
.B(n_15258),
.Y(n_15748)
);

INVx1_ASAP7_75t_L g15749 ( 
.A(n_15091),
.Y(n_15749)
);

INVx1_ASAP7_75t_L g15750 ( 
.A(n_15105),
.Y(n_15750)
);

AND2x2_ASAP7_75t_L g15751 ( 
.A(n_15315),
.B(n_11181),
.Y(n_15751)
);

AND2x2_ASAP7_75t_L g15752 ( 
.A(n_15004),
.B(n_11181),
.Y(n_15752)
);

NAND2xp5_ASAP7_75t_L g15753 ( 
.A(n_15140),
.B(n_11188),
.Y(n_15753)
);

INVx1_ASAP7_75t_L g15754 ( 
.A(n_15142),
.Y(n_15754)
);

AND2x2_ASAP7_75t_L g15755 ( 
.A(n_15013),
.B(n_11188),
.Y(n_15755)
);

BUFx2_ASAP7_75t_SL g15756 ( 
.A(n_15336),
.Y(n_15756)
);

INVx1_ASAP7_75t_SL g15757 ( 
.A(n_15055),
.Y(n_15757)
);

NOR2x1p5_ASAP7_75t_L g15758 ( 
.A(n_15436),
.B(n_15454),
.Y(n_15758)
);

NAND2xp5_ASAP7_75t_L g15759 ( 
.A(n_15205),
.B(n_15213),
.Y(n_15759)
);

INVx2_ASAP7_75t_SL g15760 ( 
.A(n_15031),
.Y(n_15760)
);

OR2x2_ASAP7_75t_L g15761 ( 
.A(n_14918),
.B(n_11189),
.Y(n_15761)
);

INVx1_ASAP7_75t_L g15762 ( 
.A(n_14983),
.Y(n_15762)
);

HB1xp67_ASAP7_75t_L g15763 ( 
.A(n_15313),
.Y(n_15763)
);

AND2x2_ASAP7_75t_L g15764 ( 
.A(n_15484),
.B(n_11189),
.Y(n_15764)
);

NAND4xp25_ASAP7_75t_L g15765 ( 
.A(n_15270),
.B(n_10458),
.C(n_10460),
.D(n_10457),
.Y(n_15765)
);

OR2x2_ASAP7_75t_L g15766 ( 
.A(n_15049),
.B(n_14932),
.Y(n_15766)
);

HB1xp67_ASAP7_75t_L g15767 ( 
.A(n_15339),
.Y(n_15767)
);

NAND2xp5_ASAP7_75t_L g15768 ( 
.A(n_15192),
.B(n_11198),
.Y(n_15768)
);

NAND2xp5_ASAP7_75t_L g15769 ( 
.A(n_15019),
.B(n_11198),
.Y(n_15769)
);

AND2x2_ASAP7_75t_L g15770 ( 
.A(n_15249),
.B(n_15372),
.Y(n_15770)
);

INVx1_ASAP7_75t_L g15771 ( 
.A(n_14992),
.Y(n_15771)
);

INVx1_ASAP7_75t_L g15772 ( 
.A(n_15017),
.Y(n_15772)
);

NAND2xp5_ASAP7_75t_L g15773 ( 
.A(n_15125),
.B(n_11216),
.Y(n_15773)
);

INVx1_ASAP7_75t_SL g15774 ( 
.A(n_14940),
.Y(n_15774)
);

AND2x2_ASAP7_75t_L g15775 ( 
.A(n_15443),
.B(n_11216),
.Y(n_15775)
);

INVx2_ASAP7_75t_L g15776 ( 
.A(n_15216),
.Y(n_15776)
);

AND2x4_ASAP7_75t_L g15777 ( 
.A(n_15248),
.B(n_8528),
.Y(n_15777)
);

HB1xp67_ASAP7_75t_L g15778 ( 
.A(n_15123),
.Y(n_15778)
);

INVx1_ASAP7_75t_L g15779 ( 
.A(n_15128),
.Y(n_15779)
);

AND2x2_ASAP7_75t_L g15780 ( 
.A(n_15497),
.B(n_11219),
.Y(n_15780)
);

INVx1_ASAP7_75t_L g15781 ( 
.A(n_15030),
.Y(n_15781)
);

NAND2xp5_ASAP7_75t_L g15782 ( 
.A(n_15332),
.B(n_11219),
.Y(n_15782)
);

INVx1_ASAP7_75t_L g15783 ( 
.A(n_15036),
.Y(n_15783)
);

BUFx2_ASAP7_75t_L g15784 ( 
.A(n_15406),
.Y(n_15784)
);

OAI22xp5_ASAP7_75t_L g15785 ( 
.A1(n_15070),
.A2(n_11365),
.B1(n_7870),
.B2(n_7711),
.Y(n_15785)
);

NAND2xp5_ASAP7_75t_L g15786 ( 
.A(n_15311),
.B(n_15269),
.Y(n_15786)
);

INVx1_ASAP7_75t_L g15787 ( 
.A(n_15194),
.Y(n_15787)
);

OR2x2_ASAP7_75t_L g15788 ( 
.A(n_14952),
.B(n_11224),
.Y(n_15788)
);

AND2x2_ASAP7_75t_L g15789 ( 
.A(n_15499),
.B(n_15509),
.Y(n_15789)
);

OR2x2_ASAP7_75t_L g15790 ( 
.A(n_15223),
.B(n_11224),
.Y(n_15790)
);

INVx1_ASAP7_75t_L g15791 ( 
.A(n_15274),
.Y(n_15791)
);

INVx1_ASAP7_75t_L g15792 ( 
.A(n_15275),
.Y(n_15792)
);

HB1xp67_ASAP7_75t_L g15793 ( 
.A(n_15179),
.Y(n_15793)
);

INVx2_ASAP7_75t_L g15794 ( 
.A(n_15220),
.Y(n_15794)
);

BUFx2_ASAP7_75t_L g15795 ( 
.A(n_14976),
.Y(n_15795)
);

NAND2xp5_ASAP7_75t_L g15796 ( 
.A(n_15277),
.B(n_11225),
.Y(n_15796)
);

AND2x4_ASAP7_75t_L g15797 ( 
.A(n_15518),
.B(n_8528),
.Y(n_15797)
);

AND2x4_ASAP7_75t_L g15798 ( 
.A(n_14997),
.B(n_8528),
.Y(n_15798)
);

NAND2xp5_ASAP7_75t_L g15799 ( 
.A(n_15224),
.B(n_11225),
.Y(n_15799)
);

OR2x2_ASAP7_75t_L g15800 ( 
.A(n_15242),
.B(n_11233),
.Y(n_15800)
);

NAND2xp5_ASAP7_75t_L g15801 ( 
.A(n_14982),
.B(n_11233),
.Y(n_15801)
);

AND2x2_ASAP7_75t_L g15802 ( 
.A(n_15433),
.B(n_11250),
.Y(n_15802)
);

AND2x2_ASAP7_75t_L g15803 ( 
.A(n_15414),
.B(n_11250),
.Y(n_15803)
);

OR2x2_ASAP7_75t_L g15804 ( 
.A(n_14963),
.B(n_11252),
.Y(n_15804)
);

INVx1_ASAP7_75t_L g15805 ( 
.A(n_15006),
.Y(n_15805)
);

AND2x2_ASAP7_75t_L g15806 ( 
.A(n_15421),
.B(n_11252),
.Y(n_15806)
);

NAND2xp5_ASAP7_75t_L g15807 ( 
.A(n_14988),
.B(n_11254),
.Y(n_15807)
);

INVx2_ASAP7_75t_L g15808 ( 
.A(n_15394),
.Y(n_15808)
);

NAND2x1p5_ASAP7_75t_L g15809 ( 
.A(n_15496),
.B(n_15510),
.Y(n_15809)
);

HB1xp67_ASAP7_75t_L g15810 ( 
.A(n_15085),
.Y(n_15810)
);

AND2x2_ASAP7_75t_L g15811 ( 
.A(n_15130),
.B(n_11254),
.Y(n_15811)
);

AND2x2_ASAP7_75t_L g15812 ( 
.A(n_15382),
.B(n_11266),
.Y(n_15812)
);

HB1xp67_ASAP7_75t_L g15813 ( 
.A(n_15272),
.Y(n_15813)
);

INVx2_ASAP7_75t_L g15814 ( 
.A(n_15281),
.Y(n_15814)
);

AND2x4_ASAP7_75t_SL g15815 ( 
.A(n_14999),
.B(n_6907),
.Y(n_15815)
);

INVx1_ASAP7_75t_SL g15816 ( 
.A(n_14958),
.Y(n_15816)
);

INVx1_ASAP7_75t_L g15817 ( 
.A(n_15014),
.Y(n_15817)
);

INVx2_ASAP7_75t_L g15818 ( 
.A(n_15025),
.Y(n_15818)
);

NOR2xp33_ASAP7_75t_L g15819 ( 
.A(n_15463),
.B(n_11266),
.Y(n_15819)
);

AND2x2_ASAP7_75t_L g15820 ( 
.A(n_15027),
.B(n_11268),
.Y(n_15820)
);

INVx1_ASAP7_75t_L g15821 ( 
.A(n_15032),
.Y(n_15821)
);

INVx2_ASAP7_75t_SL g15822 ( 
.A(n_15137),
.Y(n_15822)
);

INVx1_ASAP7_75t_SL g15823 ( 
.A(n_15086),
.Y(n_15823)
);

AND2x2_ASAP7_75t_L g15824 ( 
.A(n_15033),
.B(n_15423),
.Y(n_15824)
);

INVx1_ASAP7_75t_L g15825 ( 
.A(n_15143),
.Y(n_15825)
);

HB1xp67_ASAP7_75t_L g15826 ( 
.A(n_15286),
.Y(n_15826)
);

INVx1_ASAP7_75t_L g15827 ( 
.A(n_15204),
.Y(n_15827)
);

AND2x2_ASAP7_75t_L g15828 ( 
.A(n_15417),
.B(n_11268),
.Y(n_15828)
);

AND2x4_ASAP7_75t_SL g15829 ( 
.A(n_15456),
.B(n_7042),
.Y(n_15829)
);

AOI221xp5_ASAP7_75t_L g15830 ( 
.A1(n_15380),
.A2(n_9257),
.B1(n_9264),
.B2(n_9256),
.C(n_9237),
.Y(n_15830)
);

NAND2xp5_ASAP7_75t_L g15831 ( 
.A(n_14990),
.B(n_11274),
.Y(n_15831)
);

AND2x2_ASAP7_75t_L g15832 ( 
.A(n_15349),
.B(n_11274),
.Y(n_15832)
);

NAND2xp5_ASAP7_75t_L g15833 ( 
.A(n_15007),
.B(n_11284),
.Y(n_15833)
);

INVx2_ASAP7_75t_L g15834 ( 
.A(n_15392),
.Y(n_15834)
);

INVx1_ASAP7_75t_L g15835 ( 
.A(n_15217),
.Y(n_15835)
);

AND2x2_ASAP7_75t_L g15836 ( 
.A(n_15294),
.B(n_11284),
.Y(n_15836)
);

INVx1_ASAP7_75t_L g15837 ( 
.A(n_14931),
.Y(n_15837)
);

OR2x2_ASAP7_75t_L g15838 ( 
.A(n_14944),
.B(n_11285),
.Y(n_15838)
);

AND2x2_ASAP7_75t_L g15839 ( 
.A(n_15348),
.B(n_11285),
.Y(n_15839)
);

AND2x4_ASAP7_75t_L g15840 ( 
.A(n_15355),
.B(n_8560),
.Y(n_15840)
);

INVx2_ASAP7_75t_L g15841 ( 
.A(n_15251),
.Y(n_15841)
);

INVx1_ASAP7_75t_L g15842 ( 
.A(n_15015),
.Y(n_15842)
);

INVx2_ASAP7_75t_L g15843 ( 
.A(n_15153),
.Y(n_15843)
);

INVx2_ASAP7_75t_L g15844 ( 
.A(n_15252),
.Y(n_15844)
);

INVx1_ASAP7_75t_L g15845 ( 
.A(n_14971),
.Y(n_15845)
);

AND2x2_ASAP7_75t_L g15846 ( 
.A(n_14920),
.B(n_11286),
.Y(n_15846)
);

AND2x2_ASAP7_75t_L g15847 ( 
.A(n_14955),
.B(n_11286),
.Y(n_15847)
);

AND2x2_ASAP7_75t_L g15848 ( 
.A(n_15016),
.B(n_11294),
.Y(n_15848)
);

NAND2xp5_ASAP7_75t_L g15849 ( 
.A(n_15082),
.B(n_11294),
.Y(n_15849)
);

OR2x2_ASAP7_75t_L g15850 ( 
.A(n_15041),
.B(n_11295),
.Y(n_15850)
);

AND2x2_ASAP7_75t_L g15851 ( 
.A(n_15146),
.B(n_11295),
.Y(n_15851)
);

INVxp67_ASAP7_75t_SL g15852 ( 
.A(n_14942),
.Y(n_15852)
);

OR2x2_ASAP7_75t_L g15853 ( 
.A(n_15300),
.B(n_11303),
.Y(n_15853)
);

NAND2xp5_ASAP7_75t_L g15854 ( 
.A(n_15083),
.B(n_11303),
.Y(n_15854)
);

INVx2_ASAP7_75t_L g15855 ( 
.A(n_15475),
.Y(n_15855)
);

NAND2xp5_ASAP7_75t_L g15856 ( 
.A(n_15283),
.B(n_11306),
.Y(n_15856)
);

INVx1_ASAP7_75t_L g15857 ( 
.A(n_15389),
.Y(n_15857)
);

AND2x2_ASAP7_75t_L g15858 ( 
.A(n_15473),
.B(n_11306),
.Y(n_15858)
);

INVx2_ASAP7_75t_L g15859 ( 
.A(n_15129),
.Y(n_15859)
);

AOI22xp33_ASAP7_75t_SL g15860 ( 
.A1(n_14949),
.A2(n_9753),
.B1(n_9994),
.B2(n_10383),
.Y(n_15860)
);

AND2x4_ASAP7_75t_L g15861 ( 
.A(n_15478),
.B(n_8560),
.Y(n_15861)
);

AND2x2_ASAP7_75t_L g15862 ( 
.A(n_15366),
.B(n_11309),
.Y(n_15862)
);

AND2x2_ASAP7_75t_L g15863 ( 
.A(n_15370),
.B(n_11309),
.Y(n_15863)
);

INVx2_ASAP7_75t_L g15864 ( 
.A(n_15422),
.Y(n_15864)
);

NOR2xp33_ASAP7_75t_L g15865 ( 
.A(n_15218),
.B(n_11312),
.Y(n_15865)
);

INVx2_ASAP7_75t_L g15866 ( 
.A(n_15492),
.Y(n_15866)
);

AND2x2_ASAP7_75t_L g15867 ( 
.A(n_15522),
.B(n_11312),
.Y(n_15867)
);

NAND2xp5_ASAP7_75t_L g15868 ( 
.A(n_15291),
.B(n_11313),
.Y(n_15868)
);

AND2x2_ASAP7_75t_L g15869 ( 
.A(n_15268),
.B(n_11313),
.Y(n_15869)
);

INVx1_ASAP7_75t_L g15870 ( 
.A(n_15107),
.Y(n_15870)
);

OR2x2_ASAP7_75t_L g15871 ( 
.A(n_15358),
.B(n_11322),
.Y(n_15871)
);

INVx1_ASAP7_75t_L g15872 ( 
.A(n_15345),
.Y(n_15872)
);

AOI211xp5_ASAP7_75t_L g15873 ( 
.A1(n_15149),
.A2(n_10393),
.B(n_10405),
.C(n_7383),
.Y(n_15873)
);

AND2x2_ASAP7_75t_L g15874 ( 
.A(n_15320),
.B(n_11322),
.Y(n_15874)
);

INVx1_ASAP7_75t_L g15875 ( 
.A(n_15352),
.Y(n_15875)
);

AND2x2_ASAP7_75t_L g15876 ( 
.A(n_15304),
.B(n_11323),
.Y(n_15876)
);

OR2x2_ASAP7_75t_L g15877 ( 
.A(n_15457),
.B(n_11323),
.Y(n_15877)
);

HB1xp67_ASAP7_75t_L g15878 ( 
.A(n_15286),
.Y(n_15878)
);

AND2x2_ASAP7_75t_L g15879 ( 
.A(n_14925),
.B(n_11327),
.Y(n_15879)
);

AND2x2_ASAP7_75t_L g15880 ( 
.A(n_15354),
.B(n_11327),
.Y(n_15880)
);

INVx1_ASAP7_75t_L g15881 ( 
.A(n_15265),
.Y(n_15881)
);

AND2x2_ASAP7_75t_L g15882 ( 
.A(n_15375),
.B(n_11330),
.Y(n_15882)
);

INVx2_ASAP7_75t_L g15883 ( 
.A(n_15097),
.Y(n_15883)
);

AND2x2_ASAP7_75t_L g15884 ( 
.A(n_15353),
.B(n_15474),
.Y(n_15884)
);

AND2x2_ASAP7_75t_L g15885 ( 
.A(n_15219),
.B(n_11330),
.Y(n_15885)
);

NAND2xp5_ASAP7_75t_L g15886 ( 
.A(n_15235),
.B(n_15236),
.Y(n_15886)
);

NOR2xp33_ASAP7_75t_L g15887 ( 
.A(n_15237),
.B(n_11331),
.Y(n_15887)
);

AND2x4_ASAP7_75t_L g15888 ( 
.A(n_15240),
.B(n_8560),
.Y(n_15888)
);

AND2x2_ASAP7_75t_L g15889 ( 
.A(n_15212),
.B(n_11331),
.Y(n_15889)
);

INVx2_ASAP7_75t_L g15890 ( 
.A(n_15139),
.Y(n_15890)
);

INVx2_ASAP7_75t_L g15891 ( 
.A(n_15155),
.Y(n_15891)
);

NAND2xp5_ASAP7_75t_L g15892 ( 
.A(n_15362),
.B(n_11332),
.Y(n_15892)
);

INVx1_ASAP7_75t_L g15893 ( 
.A(n_15253),
.Y(n_15893)
);

NAND2xp5_ASAP7_75t_L g15894 ( 
.A(n_15365),
.B(n_11332),
.Y(n_15894)
);

OR2x2_ASAP7_75t_L g15895 ( 
.A(n_15168),
.B(n_11339),
.Y(n_15895)
);

INVx2_ASAP7_75t_L g15896 ( 
.A(n_15451),
.Y(n_15896)
);

AND2x2_ASAP7_75t_L g15897 ( 
.A(n_15214),
.B(n_15225),
.Y(n_15897)
);

INVx1_ASAP7_75t_L g15898 ( 
.A(n_15133),
.Y(n_15898)
);

HB1xp67_ASAP7_75t_L g15899 ( 
.A(n_15087),
.Y(n_15899)
);

NAND2xp5_ASAP7_75t_L g15900 ( 
.A(n_15385),
.B(n_11339),
.Y(n_15900)
);

INVx2_ASAP7_75t_L g15901 ( 
.A(n_15257),
.Y(n_15901)
);

INVx1_ASAP7_75t_L g15902 ( 
.A(n_15333),
.Y(n_15902)
);

NAND2xp5_ASAP7_75t_L g15903 ( 
.A(n_15199),
.B(n_11342),
.Y(n_15903)
);

AOI22xp33_ASAP7_75t_L g15904 ( 
.A1(n_15039),
.A2(n_15368),
.B1(n_15065),
.B2(n_15412),
.Y(n_15904)
);

INVx2_ASAP7_75t_L g15905 ( 
.A(n_15102),
.Y(n_15905)
);

AND2x2_ASAP7_75t_L g15906 ( 
.A(n_15331),
.B(n_11342),
.Y(n_15906)
);

INVx1_ASAP7_75t_L g15907 ( 
.A(n_15195),
.Y(n_15907)
);

AND2x2_ASAP7_75t_L g15908 ( 
.A(n_15462),
.B(n_11352),
.Y(n_15908)
);

NAND2xp5_ASAP7_75t_L g15909 ( 
.A(n_15334),
.B(n_11352),
.Y(n_15909)
);

INVx2_ASAP7_75t_L g15910 ( 
.A(n_15114),
.Y(n_15910)
);

AND2x4_ASAP7_75t_L g15911 ( 
.A(n_15337),
.B(n_8560),
.Y(n_15911)
);

AND2x4_ASAP7_75t_SL g15912 ( 
.A(n_15430),
.B(n_7042),
.Y(n_15912)
);

HB1xp67_ASAP7_75t_L g15913 ( 
.A(n_15296),
.Y(n_15913)
);

INVx2_ASAP7_75t_L g15914 ( 
.A(n_15094),
.Y(n_15914)
);

AND2x2_ASAP7_75t_L g15915 ( 
.A(n_15476),
.B(n_11353),
.Y(n_15915)
);

NAND2xp5_ASAP7_75t_L g15916 ( 
.A(n_15344),
.B(n_11353),
.Y(n_15916)
);

NAND2xp5_ASAP7_75t_L g15917 ( 
.A(n_15346),
.B(n_11355),
.Y(n_15917)
);

INVx2_ASAP7_75t_L g15918 ( 
.A(n_15324),
.Y(n_15918)
);

INVx1_ASAP7_75t_L g15919 ( 
.A(n_15111),
.Y(n_15919)
);

INVx1_ASAP7_75t_L g15920 ( 
.A(n_15104),
.Y(n_15920)
);

INVx1_ASAP7_75t_L g15921 ( 
.A(n_15159),
.Y(n_15921)
);

AND2x4_ASAP7_75t_L g15922 ( 
.A(n_15232),
.B(n_8560),
.Y(n_15922)
);

OR2x2_ASAP7_75t_L g15923 ( 
.A(n_15387),
.B(n_11355),
.Y(n_15923)
);

AND2x2_ASAP7_75t_L g15924 ( 
.A(n_15166),
.B(n_11360),
.Y(n_15924)
);

INVx1_ASAP7_75t_L g15925 ( 
.A(n_15170),
.Y(n_15925)
);

AND2x2_ASAP7_75t_L g15926 ( 
.A(n_15171),
.B(n_11360),
.Y(n_15926)
);

AND2x2_ASAP7_75t_L g15927 ( 
.A(n_15141),
.B(n_11372),
.Y(n_15927)
);

INVx2_ASAP7_75t_L g15928 ( 
.A(n_15193),
.Y(n_15928)
);

AND2x2_ASAP7_75t_L g15929 ( 
.A(n_15160),
.B(n_11372),
.Y(n_15929)
);

HB1xp67_ASAP7_75t_L g15930 ( 
.A(n_15296),
.Y(n_15930)
);

NAND2xp5_ASAP7_75t_L g15931 ( 
.A(n_15180),
.B(n_11378),
.Y(n_15931)
);

INVx3_ASAP7_75t_L g15932 ( 
.A(n_15328),
.Y(n_15932)
);

AND2x4_ASAP7_75t_L g15933 ( 
.A(n_15477),
.B(n_11208),
.Y(n_15933)
);

NAND2xp5_ASAP7_75t_L g15934 ( 
.A(n_15181),
.B(n_11378),
.Y(n_15934)
);

INVx1_ASAP7_75t_L g15935 ( 
.A(n_15256),
.Y(n_15935)
);

INVx1_ASAP7_75t_L g15936 ( 
.A(n_15109),
.Y(n_15936)
);

INVx2_ASAP7_75t_L g15937 ( 
.A(n_15276),
.Y(n_15937)
);

NAND2xp5_ASAP7_75t_L g15938 ( 
.A(n_15227),
.B(n_11381),
.Y(n_15938)
);

NAND2xp5_ASAP7_75t_L g15939 ( 
.A(n_15230),
.B(n_11381),
.Y(n_15939)
);

AND2x2_ASAP7_75t_L g15940 ( 
.A(n_15234),
.B(n_11399),
.Y(n_15940)
);

AND2x2_ASAP7_75t_L g15941 ( 
.A(n_15371),
.B(n_11399),
.Y(n_15941)
);

NAND2xp5_ASAP7_75t_L g15942 ( 
.A(n_15441),
.B(n_11403),
.Y(n_15942)
);

BUFx2_ASAP7_75t_L g15943 ( 
.A(n_15477),
.Y(n_15943)
);

INVx1_ASAP7_75t_L g15944 ( 
.A(n_15323),
.Y(n_15944)
);

HB1xp67_ASAP7_75t_L g15945 ( 
.A(n_15512),
.Y(n_15945)
);

NAND4xp25_ASAP7_75t_L g15946 ( 
.A(n_15116),
.B(n_10458),
.C(n_10460),
.D(n_10457),
.Y(n_15946)
);

OR2x2_ASAP7_75t_L g15947 ( 
.A(n_15088),
.B(n_11403),
.Y(n_15947)
);

INVx2_ASAP7_75t_L g15948 ( 
.A(n_15440),
.Y(n_15948)
);

INVxp67_ASAP7_75t_L g15949 ( 
.A(n_15056),
.Y(n_15949)
);

INVx1_ASAP7_75t_L g15950 ( 
.A(n_15093),
.Y(n_15950)
);

AND2x2_ASAP7_75t_L g15951 ( 
.A(n_15384),
.B(n_15264),
.Y(n_15951)
);

INVx2_ASAP7_75t_L g15952 ( 
.A(n_15467),
.Y(n_15952)
);

AND2x2_ASAP7_75t_L g15953 ( 
.A(n_15266),
.B(n_11405),
.Y(n_15953)
);

NAND2xp5_ASAP7_75t_L g15954 ( 
.A(n_15172),
.B(n_11405),
.Y(n_15954)
);

NAND2xp5_ASAP7_75t_L g15955 ( 
.A(n_15206),
.B(n_11406),
.Y(n_15955)
);

NAND2x1p5_ASAP7_75t_L g15956 ( 
.A(n_15132),
.B(n_15512),
.Y(n_15956)
);

AND2x2_ASAP7_75t_L g15957 ( 
.A(n_15279),
.B(n_11406),
.Y(n_15957)
);

AND2x4_ASAP7_75t_L g15958 ( 
.A(n_15489),
.B(n_15390),
.Y(n_15958)
);

OR2x2_ASAP7_75t_L g15959 ( 
.A(n_15407),
.B(n_11419),
.Y(n_15959)
);

CKINVDCx5p33_ASAP7_75t_R g15960 ( 
.A(n_15393),
.Y(n_15960)
);

NAND2xp5_ASAP7_75t_L g15961 ( 
.A(n_15479),
.B(n_11419),
.Y(n_15961)
);

AND2x4_ASAP7_75t_L g15962 ( 
.A(n_15399),
.B(n_8592),
.Y(n_15962)
);

NAND2xp5_ASAP7_75t_L g15963 ( 
.A(n_15409),
.B(n_15415),
.Y(n_15963)
);

OR2x2_ASAP7_75t_L g15964 ( 
.A(n_15061),
.B(n_11424),
.Y(n_15964)
);

AND2x4_ASAP7_75t_L g15965 ( 
.A(n_15448),
.B(n_8592),
.Y(n_15965)
);

INVx1_ASAP7_75t_SL g15966 ( 
.A(n_15259),
.Y(n_15966)
);

INVx2_ASAP7_75t_L g15967 ( 
.A(n_15469),
.Y(n_15967)
);

INVx1_ASAP7_75t_L g15968 ( 
.A(n_15096),
.Y(n_15968)
);

AND2x2_ASAP7_75t_L g15969 ( 
.A(n_15245),
.B(n_11424),
.Y(n_15969)
);

AND2x2_ASAP7_75t_L g15970 ( 
.A(n_15254),
.B(n_11425),
.Y(n_15970)
);

INVx4_ASAP7_75t_L g15971 ( 
.A(n_15450),
.Y(n_15971)
);

INVx1_ASAP7_75t_SL g15972 ( 
.A(n_15357),
.Y(n_15972)
);

INVx1_ASAP7_75t_L g15973 ( 
.A(n_15186),
.Y(n_15973)
);

NAND2xp5_ASAP7_75t_L g15974 ( 
.A(n_15305),
.B(n_11425),
.Y(n_15974)
);

NOR2xp33_ASAP7_75t_L g15975 ( 
.A(n_15405),
.B(n_11429),
.Y(n_15975)
);

INVxp67_ASAP7_75t_L g15976 ( 
.A(n_15060),
.Y(n_15976)
);

NAND3xp33_ASAP7_75t_L g15977 ( 
.A(n_15066),
.B(n_11267),
.C(n_9753),
.Y(n_15977)
);

INVx2_ASAP7_75t_L g15978 ( 
.A(n_15470),
.Y(n_15978)
);

NAND2xp5_ASAP7_75t_L g15979 ( 
.A(n_15516),
.B(n_11429),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15118),
.Y(n_15980)
);

NAND2xp5_ASAP7_75t_L g15981 ( 
.A(n_15340),
.B(n_11438),
.Y(n_15981)
);

AND2x2_ASAP7_75t_L g15982 ( 
.A(n_15261),
.B(n_11438),
.Y(n_15982)
);

NAND2xp5_ASAP7_75t_L g15983 ( 
.A(n_15263),
.B(n_11439),
.Y(n_15983)
);

INVx1_ASAP7_75t_L g15984 ( 
.A(n_15144),
.Y(n_15984)
);

AND2x2_ASAP7_75t_SL g15985 ( 
.A(n_15062),
.B(n_8923),
.Y(n_15985)
);

NOR2xp33_ASAP7_75t_L g15986 ( 
.A(n_15293),
.B(n_11439),
.Y(n_15986)
);

NAND2xp5_ASAP7_75t_SL g15987 ( 
.A(n_15410),
.B(n_8340),
.Y(n_15987)
);

OR2x2_ASAP7_75t_L g15988 ( 
.A(n_15307),
.B(n_11441),
.Y(n_15988)
);

INVx2_ASAP7_75t_L g15989 ( 
.A(n_15100),
.Y(n_15989)
);

NAND2xp5_ASAP7_75t_L g15990 ( 
.A(n_15120),
.B(n_11441),
.Y(n_15990)
);

INVx1_ASAP7_75t_L g15991 ( 
.A(n_15161),
.Y(n_15991)
);

AND2x2_ASAP7_75t_L g15992 ( 
.A(n_15103),
.B(n_11445),
.Y(n_15992)
);

INVx1_ASAP7_75t_L g15993 ( 
.A(n_15167),
.Y(n_15993)
);

INVx1_ASAP7_75t_L g15994 ( 
.A(n_15174),
.Y(n_15994)
);

AND2x2_ASAP7_75t_L g15995 ( 
.A(n_15285),
.B(n_11445),
.Y(n_15995)
);

INVx2_ASAP7_75t_SL g15996 ( 
.A(n_15373),
.Y(n_15996)
);

NAND3xp33_ASAP7_75t_L g15997 ( 
.A(n_15063),
.B(n_11267),
.C(n_11458),
.Y(n_15997)
);

AND2x2_ASAP7_75t_L g15998 ( 
.A(n_15503),
.B(n_11458),
.Y(n_15998)
);

NAND2xp5_ASAP7_75t_L g15999 ( 
.A(n_15317),
.B(n_11469),
.Y(n_15999)
);

INVx2_ASAP7_75t_SL g16000 ( 
.A(n_15396),
.Y(n_16000)
);

AND2x4_ASAP7_75t_SL g16001 ( 
.A(n_15356),
.B(n_7042),
.Y(n_16001)
);

INVx1_ASAP7_75t_L g16002 ( 
.A(n_15182),
.Y(n_16002)
);

OR2x2_ASAP7_75t_L g16003 ( 
.A(n_15310),
.B(n_15444),
.Y(n_16003)
);

AND2x2_ASAP7_75t_L g16004 ( 
.A(n_15327),
.B(n_11469),
.Y(n_16004)
);

AND2x2_ASAP7_75t_L g16005 ( 
.A(n_15322),
.B(n_11471),
.Y(n_16005)
);

INVx1_ASAP7_75t_L g16006 ( 
.A(n_15188),
.Y(n_16006)
);

INVx4_ASAP7_75t_L g16007 ( 
.A(n_15517),
.Y(n_16007)
);

HB1xp67_ASAP7_75t_L g16008 ( 
.A(n_15233),
.Y(n_16008)
);

INVx1_ASAP7_75t_L g16009 ( 
.A(n_15191),
.Y(n_16009)
);

AND2x2_ASAP7_75t_L g16010 ( 
.A(n_15325),
.B(n_11471),
.Y(n_16010)
);

AND2x2_ASAP7_75t_L g16011 ( 
.A(n_15330),
.B(n_11474),
.Y(n_16011)
);

NOR2xp67_ASAP7_75t_L g16012 ( 
.A(n_15439),
.B(n_11474),
.Y(n_16012)
);

AND2x2_ASAP7_75t_L g16013 ( 
.A(n_15335),
.B(n_11477),
.Y(n_16013)
);

INVx1_ASAP7_75t_L g16014 ( 
.A(n_15150),
.Y(n_16014)
);

INVx2_ASAP7_75t_L g16015 ( 
.A(n_15359),
.Y(n_16015)
);

INVx1_ASAP7_75t_L g16016 ( 
.A(n_15158),
.Y(n_16016)
);

BUFx2_ASAP7_75t_L g16017 ( 
.A(n_15428),
.Y(n_16017)
);

NAND2xp5_ASAP7_75t_L g16018 ( 
.A(n_15319),
.B(n_11477),
.Y(n_16018)
);

OR2x2_ASAP7_75t_L g16019 ( 
.A(n_15464),
.B(n_11485),
.Y(n_16019)
);

INVx1_ASAP7_75t_L g16020 ( 
.A(n_15231),
.Y(n_16020)
);

INVx1_ASAP7_75t_SL g16021 ( 
.A(n_15419),
.Y(n_16021)
);

INVx1_ASAP7_75t_L g16022 ( 
.A(n_15241),
.Y(n_16022)
);

AND2x2_ASAP7_75t_L g16023 ( 
.A(n_15343),
.B(n_11485),
.Y(n_16023)
);

AND2x2_ASAP7_75t_L g16024 ( 
.A(n_15361),
.B(n_11498),
.Y(n_16024)
);

OR2x2_ASAP7_75t_L g16025 ( 
.A(n_15287),
.B(n_11498),
.Y(n_16025)
);

OR2x2_ASAP7_75t_L g16026 ( 
.A(n_15401),
.B(n_11508),
.Y(n_16026)
);

INVx1_ASAP7_75t_L g16027 ( 
.A(n_15113),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15122),
.Y(n_16028)
);

INVx1_ASAP7_75t_L g16029 ( 
.A(n_15309),
.Y(n_16029)
);

OR2x2_ASAP7_75t_L g16030 ( 
.A(n_15207),
.B(n_11508),
.Y(n_16030)
);

NAND2xp5_ASAP7_75t_L g16031 ( 
.A(n_15374),
.B(n_11510),
.Y(n_16031)
);

INVx1_ASAP7_75t_L g16032 ( 
.A(n_15152),
.Y(n_16032)
);

OR2x2_ASAP7_75t_L g16033 ( 
.A(n_15221),
.B(n_11510),
.Y(n_16033)
);

OR2x2_ASAP7_75t_L g16034 ( 
.A(n_15326),
.B(n_11515),
.Y(n_16034)
);

CKINVDCx20_ASAP7_75t_R g16035 ( 
.A(n_15519),
.Y(n_16035)
);

NAND2xp5_ASAP7_75t_L g16036 ( 
.A(n_15383),
.B(n_11515),
.Y(n_16036)
);

INVx1_ASAP7_75t_L g16037 ( 
.A(n_15156),
.Y(n_16037)
);

INVx3_ASAP7_75t_L g16038 ( 
.A(n_15367),
.Y(n_16038)
);

INVx1_ASAP7_75t_SL g16039 ( 
.A(n_15404),
.Y(n_16039)
);

INVx1_ASAP7_75t_L g16040 ( 
.A(n_15239),
.Y(n_16040)
);

AND2x2_ASAP7_75t_L g16041 ( 
.A(n_15388),
.B(n_15395),
.Y(n_16041)
);

INVx1_ASAP7_75t_SL g16042 ( 
.A(n_15438),
.Y(n_16042)
);

AND2x2_ASAP7_75t_L g16043 ( 
.A(n_15397),
.B(n_11524),
.Y(n_16043)
);

INVx1_ASAP7_75t_L g16044 ( 
.A(n_15250),
.Y(n_16044)
);

OAI22xp5_ASAP7_75t_L g16045 ( 
.A1(n_15386),
.A2(n_11365),
.B1(n_7870),
.B2(n_7711),
.Y(n_16045)
);

NAND2xp5_ASAP7_75t_L g16046 ( 
.A(n_15398),
.B(n_11524),
.Y(n_16046)
);

INVx3_ASAP7_75t_L g16047 ( 
.A(n_15520),
.Y(n_16047)
);

AND2x2_ASAP7_75t_L g16048 ( 
.A(n_15400),
.B(n_11530),
.Y(n_16048)
);

OR2x2_ASAP7_75t_L g16049 ( 
.A(n_15338),
.B(n_11530),
.Y(n_16049)
);

INVx1_ASAP7_75t_L g16050 ( 
.A(n_15297),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15403),
.B(n_11541),
.Y(n_16051)
);

AND2x4_ASAP7_75t_L g16052 ( 
.A(n_15521),
.B(n_15431),
.Y(n_16052)
);

NAND2xp5_ASAP7_75t_L g16053 ( 
.A(n_15411),
.B(n_11541),
.Y(n_16053)
);

AND2x2_ASAP7_75t_L g16054 ( 
.A(n_15481),
.B(n_11218),
.Y(n_16054)
);

INVx1_ASAP7_75t_L g16055 ( 
.A(n_15299),
.Y(n_16055)
);

INVx1_ASAP7_75t_SL g16056 ( 
.A(n_15360),
.Y(n_16056)
);

OR2x2_ASAP7_75t_L g16057 ( 
.A(n_15135),
.B(n_15288),
.Y(n_16057)
);

BUFx2_ASAP7_75t_L g16058 ( 
.A(n_15432),
.Y(n_16058)
);

OR2x2_ASAP7_75t_L g16059 ( 
.A(n_15943),
.B(n_15298),
.Y(n_16059)
);

INVx1_ASAP7_75t_L g16060 ( 
.A(n_15943),
.Y(n_16060)
);

NOR2xp67_ASAP7_75t_L g16061 ( 
.A(n_15945),
.B(n_15465),
.Y(n_16061)
);

AND2x2_ASAP7_75t_L g16062 ( 
.A(n_15585),
.B(n_15435),
.Y(n_16062)
);

INVx2_ASAP7_75t_L g16063 ( 
.A(n_15665),
.Y(n_16063)
);

AND2x2_ASAP7_75t_L g16064 ( 
.A(n_15536),
.B(n_15445),
.Y(n_16064)
);

NAND2x1_ASAP7_75t_SL g16065 ( 
.A(n_15778),
.B(n_15442),
.Y(n_16065)
);

BUFx3_ASAP7_75t_L g16066 ( 
.A(n_15595),
.Y(n_16066)
);

AND2x2_ASAP7_75t_L g16067 ( 
.A(n_15559),
.B(n_15447),
.Y(n_16067)
);

NAND4xp25_ASAP7_75t_L g16068 ( 
.A(n_15537),
.B(n_15425),
.C(n_15466),
.D(n_15437),
.Y(n_16068)
);

AND2x2_ASAP7_75t_L g16069 ( 
.A(n_15524),
.B(n_15458),
.Y(n_16069)
);

BUFx2_ASAP7_75t_SL g16070 ( 
.A(n_15652),
.Y(n_16070)
);

INVx2_ASAP7_75t_L g16071 ( 
.A(n_15671),
.Y(n_16071)
);

INVxp33_ASAP7_75t_L g16072 ( 
.A(n_15809),
.Y(n_16072)
);

INVx1_ASAP7_75t_L g16073 ( 
.A(n_15599),
.Y(n_16073)
);

INVx1_ASAP7_75t_L g16074 ( 
.A(n_15599),
.Y(n_16074)
);

NAND2xp5_ASAP7_75t_L g16075 ( 
.A(n_15722),
.B(n_15461),
.Y(n_16075)
);

INVxp67_ASAP7_75t_L g16076 ( 
.A(n_15756),
.Y(n_16076)
);

AND2x2_ASAP7_75t_L g16077 ( 
.A(n_15630),
.B(n_15590),
.Y(n_16077)
);

NAND3xp33_ASAP7_75t_L g16078 ( 
.A(n_15589),
.B(n_15472),
.C(n_15471),
.Y(n_16078)
);

NAND2xp5_ASAP7_75t_L g16079 ( 
.A(n_15743),
.B(n_15480),
.Y(n_16079)
);

INVx1_ASAP7_75t_L g16080 ( 
.A(n_15709),
.Y(n_16080)
);

AND2x2_ASAP7_75t_L g16081 ( 
.A(n_15528),
.B(n_15482),
.Y(n_16081)
);

INVx1_ASAP7_75t_L g16082 ( 
.A(n_15709),
.Y(n_16082)
);

NAND2xp5_ASAP7_75t_SL g16083 ( 
.A(n_15615),
.B(n_15306),
.Y(n_16083)
);

HB1xp67_ASAP7_75t_L g16084 ( 
.A(n_15576),
.Y(n_16084)
);

NAND2xp5_ASAP7_75t_L g16085 ( 
.A(n_15703),
.B(n_15485),
.Y(n_16085)
);

INVx1_ASAP7_75t_L g16086 ( 
.A(n_15533),
.Y(n_16086)
);

INVx2_ASAP7_75t_L g16087 ( 
.A(n_15671),
.Y(n_16087)
);

AND2x2_ASAP7_75t_L g16088 ( 
.A(n_15535),
.B(n_15490),
.Y(n_16088)
);

AND2x2_ASAP7_75t_L g16089 ( 
.A(n_15631),
.B(n_15582),
.Y(n_16089)
);

AND2x2_ASAP7_75t_L g16090 ( 
.A(n_15629),
.B(n_15495),
.Y(n_16090)
);

INVx1_ASAP7_75t_L g16091 ( 
.A(n_15767),
.Y(n_16091)
);

INVx1_ASAP7_75t_L g16092 ( 
.A(n_15793),
.Y(n_16092)
);

AND2x2_ASAP7_75t_L g16093 ( 
.A(n_15760),
.B(n_15505),
.Y(n_16093)
);

OAI21x1_ASAP7_75t_L g16094 ( 
.A1(n_15554),
.A2(n_15726),
.B(n_15553),
.Y(n_16094)
);

AND2x2_ASAP7_75t_L g16095 ( 
.A(n_15566),
.B(n_15506),
.Y(n_16095)
);

OAI221xp5_ASAP7_75t_L g16096 ( 
.A1(n_15904),
.A2(n_15696),
.B1(n_15687),
.B2(n_15551),
.C(n_15694),
.Y(n_16096)
);

INVx3_ASAP7_75t_L g16097 ( 
.A(n_15549),
.Y(n_16097)
);

AND2x2_ASAP7_75t_L g16098 ( 
.A(n_15824),
.B(n_15508),
.Y(n_16098)
);

INVx2_ASAP7_75t_L g16099 ( 
.A(n_15554),
.Y(n_16099)
);

AND2x2_ASAP7_75t_L g16100 ( 
.A(n_15634),
.B(n_15513),
.Y(n_16100)
);

NOR2xp33_ASAP7_75t_L g16101 ( 
.A(n_15571),
.B(n_15460),
.Y(n_16101)
);

INVx4_ASAP7_75t_L g16102 ( 
.A(n_15656),
.Y(n_16102)
);

NOR2x1_ASAP7_75t_L g16103 ( 
.A(n_15579),
.B(n_15446),
.Y(n_16103)
);

AOI322xp5_ASAP7_75t_L g16104 ( 
.A1(n_15543),
.A2(n_15364),
.A3(n_15280),
.B1(n_15434),
.B2(n_15092),
.C1(n_15453),
.C2(n_15468),
.Y(n_16104)
);

INVx4_ASAP7_75t_L g16105 ( 
.A(n_15610),
.Y(n_16105)
);

INVx2_ASAP7_75t_SL g16106 ( 
.A(n_15574),
.Y(n_16106)
);

NAND2xp5_ASAP7_75t_L g16107 ( 
.A(n_15621),
.B(n_15487),
.Y(n_16107)
);

AND2x2_ASAP7_75t_L g16108 ( 
.A(n_15628),
.B(n_15511),
.Y(n_16108)
);

OR2x2_ASAP7_75t_L g16109 ( 
.A(n_15757),
.B(n_15284),
.Y(n_16109)
);

INVx1_ASAP7_75t_L g16110 ( 
.A(n_15708),
.Y(n_16110)
);

NAND3xp33_ASAP7_75t_L g16111 ( 
.A(n_15763),
.B(n_15121),
.C(n_15488),
.Y(n_16111)
);

AOI21xp5_ASAP7_75t_L g16112 ( 
.A1(n_15784),
.A2(n_15494),
.B(n_15491),
.Y(n_16112)
);

NOR2xp33_ASAP7_75t_L g16113 ( 
.A(n_15541),
.B(n_15449),
.Y(n_16113)
);

INVx1_ASAP7_75t_L g16114 ( 
.A(n_15552),
.Y(n_16114)
);

AND2x4_ASAP7_75t_L g16115 ( 
.A(n_15734),
.B(n_15504),
.Y(n_16115)
);

AND2x2_ASAP7_75t_L g16116 ( 
.A(n_15746),
.B(n_15681),
.Y(n_16116)
);

BUFx2_ASAP7_75t_L g16117 ( 
.A(n_15577),
.Y(n_16117)
);

INVx2_ASAP7_75t_L g16118 ( 
.A(n_16017),
.Y(n_16118)
);

AND2x2_ASAP7_75t_L g16119 ( 
.A(n_15660),
.B(n_15514),
.Y(n_16119)
);

INVx1_ASAP7_75t_L g16120 ( 
.A(n_16017),
.Y(n_16120)
);

AND2x2_ASAP7_75t_L g16121 ( 
.A(n_15546),
.B(n_15493),
.Y(n_16121)
);

AND2x4_ASAP7_75t_SL g16122 ( 
.A(n_15770),
.B(n_15498),
.Y(n_16122)
);

OR2x2_ASAP7_75t_L g16123 ( 
.A(n_15648),
.B(n_15486),
.Y(n_16123)
);

INVx1_ASAP7_75t_L g16124 ( 
.A(n_15784),
.Y(n_16124)
);

AND2x2_ASAP7_75t_L g16125 ( 
.A(n_15572),
.B(n_15500),
.Y(n_16125)
);

INVx1_ASAP7_75t_L g16126 ( 
.A(n_15733),
.Y(n_16126)
);

INVx1_ASAP7_75t_L g16127 ( 
.A(n_15523),
.Y(n_16127)
);

AND2x2_ASAP7_75t_L g16128 ( 
.A(n_15560),
.B(n_15501),
.Y(n_16128)
);

NAND2x1_ASAP7_75t_L g16129 ( 
.A(n_16058),
.B(n_15864),
.Y(n_16129)
);

INVx1_ASAP7_75t_SL g16130 ( 
.A(n_15525),
.Y(n_16130)
);

AND2x2_ASAP7_75t_L g16131 ( 
.A(n_15548),
.B(n_15502),
.Y(n_16131)
);

AND2x4_ASAP7_75t_L g16132 ( 
.A(n_15758),
.B(n_15507),
.Y(n_16132)
);

NAND4xp25_ASAP7_75t_L g16133 ( 
.A(n_15557),
.B(n_15515),
.C(n_15306),
.D(n_15244),
.Y(n_16133)
);

AND2x2_ASAP7_75t_L g16134 ( 
.A(n_15555),
.B(n_15426),
.Y(n_16134)
);

INVx1_ASAP7_75t_L g16135 ( 
.A(n_15527),
.Y(n_16135)
);

AND2x2_ASAP7_75t_L g16136 ( 
.A(n_15706),
.B(n_15244),
.Y(n_16136)
);

INVx1_ASAP7_75t_SL g16137 ( 
.A(n_15774),
.Y(n_16137)
);

NAND3x1_ASAP7_75t_L g16138 ( 
.A(n_15569),
.B(n_10280),
.C(n_10189),
.Y(n_16138)
);

AND2x4_ASAP7_75t_SL g16139 ( 
.A(n_15542),
.B(n_15163),
.Y(n_16139)
);

AND2x2_ASAP7_75t_L g16140 ( 
.A(n_15562),
.B(n_15163),
.Y(n_16140)
);

BUFx3_ASAP7_75t_L g16141 ( 
.A(n_15614),
.Y(n_16141)
);

HB1xp67_ASAP7_75t_L g16142 ( 
.A(n_15866),
.Y(n_16142)
);

NOR2xp33_ASAP7_75t_L g16143 ( 
.A(n_15823),
.B(n_16042),
.Y(n_16143)
);

INVx1_ASAP7_75t_L g16144 ( 
.A(n_15600),
.Y(n_16144)
);

NAND2xp33_ASAP7_75t_SL g16145 ( 
.A(n_16035),
.B(n_15198),
.Y(n_16145)
);

HB1xp67_ASAP7_75t_L g16146 ( 
.A(n_15956),
.Y(n_16146)
);

OR2x2_ASAP7_75t_L g16147 ( 
.A(n_15538),
.B(n_15198),
.Y(n_16147)
);

NOR2xp33_ASAP7_75t_L g16148 ( 
.A(n_16021),
.B(n_15201),
.Y(n_16148)
);

INVx1_ASAP7_75t_SL g16149 ( 
.A(n_15526),
.Y(n_16149)
);

AOI22xp33_ASAP7_75t_L g16150 ( 
.A1(n_15795),
.A2(n_15201),
.B1(n_11505),
.B2(n_11385),
.Y(n_16150)
);

HB1xp67_ASAP7_75t_L g16151 ( 
.A(n_15561),
.Y(n_16151)
);

AND2x2_ASAP7_75t_L g16152 ( 
.A(n_15732),
.B(n_11218),
.Y(n_16152)
);

INVx1_ASAP7_75t_L g16153 ( 
.A(n_15606),
.Y(n_16153)
);

INVx1_ASAP7_75t_L g16154 ( 
.A(n_15540),
.Y(n_16154)
);

INVx1_ASAP7_75t_L g16155 ( 
.A(n_15547),
.Y(n_16155)
);

HB1xp67_ASAP7_75t_L g16156 ( 
.A(n_16058),
.Y(n_16156)
);

INVx1_ASAP7_75t_L g16157 ( 
.A(n_15688),
.Y(n_16157)
);

HB1xp67_ASAP7_75t_L g16158 ( 
.A(n_15570),
.Y(n_16158)
);

AND2x2_ASAP7_75t_L g16159 ( 
.A(n_15732),
.B(n_10462),
.Y(n_16159)
);

INVx1_ASAP7_75t_L g16160 ( 
.A(n_15556),
.Y(n_16160)
);

INVxp67_ASAP7_75t_L g16161 ( 
.A(n_15795),
.Y(n_16161)
);

OR2x2_ASAP7_75t_L g16162 ( 
.A(n_15564),
.B(n_10462),
.Y(n_16162)
);

INVx1_ASAP7_75t_L g16163 ( 
.A(n_15578),
.Y(n_16163)
);

AND2x2_ASAP7_75t_L g16164 ( 
.A(n_15834),
.B(n_10465),
.Y(n_16164)
);

HB1xp67_ASAP7_75t_L g16165 ( 
.A(n_15693),
.Y(n_16165)
);

INVx1_ASAP7_75t_L g16166 ( 
.A(n_15616),
.Y(n_16166)
);

AND2x4_ASAP7_75t_L g16167 ( 
.A(n_15567),
.B(n_8592),
.Y(n_16167)
);

AND2x2_ASAP7_75t_L g16168 ( 
.A(n_15897),
.B(n_10465),
.Y(n_16168)
);

NAND2xp5_ASAP7_75t_L g16169 ( 
.A(n_15619),
.B(n_9810),
.Y(n_16169)
);

HB1xp67_ASAP7_75t_L g16170 ( 
.A(n_15727),
.Y(n_16170)
);

AND2x2_ASAP7_75t_L g16171 ( 
.A(n_15822),
.B(n_15545),
.Y(n_16171)
);

INVx1_ASAP7_75t_L g16172 ( 
.A(n_15558),
.Y(n_16172)
);

INVx1_ASAP7_75t_L g16173 ( 
.A(n_15580),
.Y(n_16173)
);

NAND2xp5_ASAP7_75t_L g16174 ( 
.A(n_15724),
.B(n_15534),
.Y(n_16174)
);

NAND2xp5_ASAP7_75t_L g16175 ( 
.A(n_15573),
.B(n_15736),
.Y(n_16175)
);

INVx2_ASAP7_75t_L g16176 ( 
.A(n_15594),
.Y(n_16176)
);

INVx2_ASAP7_75t_L g16177 ( 
.A(n_15603),
.Y(n_16177)
);

NAND4xp25_ASAP7_75t_L g16178 ( 
.A(n_15748),
.B(n_10471),
.C(n_10472),
.D(n_10469),
.Y(n_16178)
);

INVx2_ASAP7_75t_SL g16179 ( 
.A(n_15598),
.Y(n_16179)
);

NOR3xp33_ASAP7_75t_L g16180 ( 
.A(n_15531),
.B(n_10583),
.C(n_10585),
.Y(n_16180)
);

INVx1_ASAP7_75t_L g16181 ( 
.A(n_15813),
.Y(n_16181)
);

INVx2_ASAP7_75t_L g16182 ( 
.A(n_15932),
.Y(n_16182)
);

INVx3_ASAP7_75t_SL g16183 ( 
.A(n_15960),
.Y(n_16183)
);

INVx1_ASAP7_75t_L g16184 ( 
.A(n_15529),
.Y(n_16184)
);

NAND2xp5_ASAP7_75t_L g16185 ( 
.A(n_15677),
.B(n_9815),
.Y(n_16185)
);

AND2x2_ASAP7_75t_L g16186 ( 
.A(n_15683),
.B(n_10469),
.Y(n_16186)
);

OR2x2_ASAP7_75t_L g16187 ( 
.A(n_15766),
.B(n_10471),
.Y(n_16187)
);

AND4x1_ASAP7_75t_L g16188 ( 
.A(n_15620),
.B(n_7572),
.C(n_7589),
.D(n_7471),
.Y(n_16188)
);

AND2x2_ASAP7_75t_L g16189 ( 
.A(n_15686),
.B(n_10472),
.Y(n_16189)
);

AND2x2_ASAP7_75t_L g16190 ( 
.A(n_15789),
.B(n_10485),
.Y(n_16190)
);

INVx1_ASAP7_75t_L g16191 ( 
.A(n_15532),
.Y(n_16191)
);

AND2x2_ASAP7_75t_L g16192 ( 
.A(n_15611),
.B(n_15884),
.Y(n_16192)
);

AND2x2_ASAP7_75t_L g16193 ( 
.A(n_15539),
.B(n_10485),
.Y(n_16193)
);

AND2x4_ASAP7_75t_L g16194 ( 
.A(n_15989),
.B(n_8592),
.Y(n_16194)
);

NAND2xp5_ASAP7_75t_L g16195 ( 
.A(n_15650),
.B(n_9815),
.Y(n_16195)
);

BUFx2_ASAP7_75t_L g16196 ( 
.A(n_15674),
.Y(n_16196)
);

OR2x2_ASAP7_75t_L g16197 ( 
.A(n_15700),
.B(n_10487),
.Y(n_16197)
);

AND3x1_ASAP7_75t_L g16198 ( 
.A(n_15843),
.B(n_10488),
.C(n_10487),
.Y(n_16198)
);

INVx2_ASAP7_75t_L g16199 ( 
.A(n_16038),
.Y(n_16199)
);

CKINVDCx5p33_ASAP7_75t_R g16200 ( 
.A(n_15810),
.Y(n_16200)
);

OR2x2_ASAP7_75t_L g16201 ( 
.A(n_15588),
.B(n_10488),
.Y(n_16201)
);

AOI21xp33_ASAP7_75t_L g16202 ( 
.A1(n_15816),
.A2(n_10493),
.B(n_10491),
.Y(n_16202)
);

AND2x2_ASAP7_75t_L g16203 ( 
.A(n_15565),
.B(n_10491),
.Y(n_16203)
);

NAND2xp33_ASAP7_75t_L g16204 ( 
.A(n_16000),
.B(n_8340),
.Y(n_16204)
);

INVx1_ASAP7_75t_L g16205 ( 
.A(n_15899),
.Y(n_16205)
);

NAND2xp5_ASAP7_75t_L g16206 ( 
.A(n_15657),
.B(n_9817),
.Y(n_16206)
);

OR2x6_ASAP7_75t_L g16207 ( 
.A(n_15818),
.B(n_6188),
.Y(n_16207)
);

BUFx2_ASAP7_75t_L g16208 ( 
.A(n_15730),
.Y(n_16208)
);

INVx2_ASAP7_75t_L g16209 ( 
.A(n_15691),
.Y(n_16209)
);

OR2x2_ASAP7_75t_L g16210 ( 
.A(n_15592),
.B(n_10493),
.Y(n_16210)
);

INVx1_ASAP7_75t_L g16211 ( 
.A(n_15635),
.Y(n_16211)
);

NAND2xp5_ASAP7_75t_L g16212 ( 
.A(n_15602),
.B(n_15705),
.Y(n_16212)
);

AND2x2_ASAP7_75t_L g16213 ( 
.A(n_15568),
.B(n_10498),
.Y(n_16213)
);

INVx2_ASAP7_75t_L g16214 ( 
.A(n_15640),
.Y(n_16214)
);

INVx1_ASAP7_75t_SL g16215 ( 
.A(n_16039),
.Y(n_16215)
);

AND2x2_ASAP7_75t_L g16216 ( 
.A(n_15841),
.B(n_10498),
.Y(n_16216)
);

AND2x2_ASAP7_75t_SL g16217 ( 
.A(n_15596),
.B(n_8923),
.Y(n_16217)
);

INVx2_ASAP7_75t_L g16218 ( 
.A(n_15575),
.Y(n_16218)
);

AOI22xp5_ASAP7_75t_L g16219 ( 
.A1(n_15737),
.A2(n_8483),
.B1(n_8494),
.B2(n_8340),
.Y(n_16219)
);

BUFx2_ASAP7_75t_L g16220 ( 
.A(n_15719),
.Y(n_16220)
);

NAND2xp5_ASAP7_75t_L g16221 ( 
.A(n_15581),
.B(n_9817),
.Y(n_16221)
);

OR2x2_ASAP7_75t_L g16222 ( 
.A(n_15883),
.B(n_10504),
.Y(n_16222)
);

NAND2xp5_ASAP7_75t_L g16223 ( 
.A(n_15584),
.B(n_9826),
.Y(n_16223)
);

INVx1_ASAP7_75t_L g16224 ( 
.A(n_16041),
.Y(n_16224)
);

AOI22xp33_ASAP7_75t_L g16225 ( 
.A1(n_15661),
.A2(n_11505),
.B1(n_11385),
.B2(n_10505),
.Y(n_16225)
);

INVx1_ASAP7_75t_L g16226 ( 
.A(n_15658),
.Y(n_16226)
);

AND2x2_ASAP7_75t_L g16227 ( 
.A(n_15859),
.B(n_10504),
.Y(n_16227)
);

AND2x2_ASAP7_75t_L g16228 ( 
.A(n_15890),
.B(n_10505),
.Y(n_16228)
);

OR2x2_ASAP7_75t_L g16229 ( 
.A(n_15891),
.B(n_8198),
.Y(n_16229)
);

INVx1_ASAP7_75t_L g16230 ( 
.A(n_15662),
.Y(n_16230)
);

NAND2xp5_ASAP7_75t_L g16231 ( 
.A(n_15586),
.B(n_9826),
.Y(n_16231)
);

OR2x2_ASAP7_75t_L g16232 ( 
.A(n_15905),
.B(n_8198),
.Y(n_16232)
);

HB1xp67_ASAP7_75t_L g16233 ( 
.A(n_16008),
.Y(n_16233)
);

INVx2_ASAP7_75t_L g16234 ( 
.A(n_15910),
.Y(n_16234)
);

AND2x2_ASAP7_75t_L g16235 ( 
.A(n_15844),
.B(n_11079),
.Y(n_16235)
);

AND2x2_ASAP7_75t_L g16236 ( 
.A(n_15901),
.B(n_16015),
.Y(n_16236)
);

NAND4xp25_ASAP7_75t_L g16237 ( 
.A(n_15976),
.B(n_7823),
.C(n_7903),
.D(n_7749),
.Y(n_16237)
);

NAND2xp5_ASAP7_75t_L g16238 ( 
.A(n_15593),
.B(n_9832),
.Y(n_16238)
);

OR2x2_ASAP7_75t_L g16239 ( 
.A(n_15896),
.B(n_8901),
.Y(n_16239)
);

OR2x2_ASAP7_75t_L g16240 ( 
.A(n_15625),
.B(n_8901),
.Y(n_16240)
);

OR2x2_ASAP7_75t_L g16241 ( 
.A(n_15914),
.B(n_15928),
.Y(n_16241)
);

OAI31xp33_ASAP7_75t_L g16242 ( 
.A1(n_15785),
.A2(n_9257),
.A3(n_9264),
.B(n_9256),
.Y(n_16242)
);

INVx1_ASAP7_75t_L g16243 ( 
.A(n_15530),
.Y(n_16243)
);

INVx1_ASAP7_75t_SL g16244 ( 
.A(n_15738),
.Y(n_16244)
);

INVx2_ASAP7_75t_L g16245 ( 
.A(n_15937),
.Y(n_16245)
);

NAND2xp5_ASAP7_75t_L g16246 ( 
.A(n_15624),
.B(n_9832),
.Y(n_16246)
);

AND2x2_ASAP7_75t_L g16247 ( 
.A(n_15618),
.B(n_11079),
.Y(n_16247)
);

INVx2_ASAP7_75t_L g16248 ( 
.A(n_15663),
.Y(n_16248)
);

BUFx2_ASAP7_75t_L g16249 ( 
.A(n_15713),
.Y(n_16249)
);

AND2x4_ASAP7_75t_L g16250 ( 
.A(n_15654),
.B(n_15948),
.Y(n_16250)
);

OR2x2_ASAP7_75t_L g16251 ( 
.A(n_15601),
.B(n_8695),
.Y(n_16251)
);

OAI21xp33_ASAP7_75t_L g16252 ( 
.A1(n_15949),
.A2(n_10583),
.B(n_10889),
.Y(n_16252)
);

AND2x2_ASAP7_75t_L g16253 ( 
.A(n_15857),
.B(n_11110),
.Y(n_16253)
);

INVx2_ASAP7_75t_L g16254 ( 
.A(n_15855),
.Y(n_16254)
);

INVx1_ASAP7_75t_L g16255 ( 
.A(n_15604),
.Y(n_16255)
);

NAND2xp5_ASAP7_75t_L g16256 ( 
.A(n_15633),
.B(n_9833),
.Y(n_16256)
);

NAND2xp5_ASAP7_75t_L g16257 ( 
.A(n_15646),
.B(n_9833),
.Y(n_16257)
);

NAND2xp5_ASAP7_75t_L g16258 ( 
.A(n_15647),
.B(n_9838),
.Y(n_16258)
);

INVx1_ASAP7_75t_SL g16259 ( 
.A(n_16056),
.Y(n_16259)
);

OR2x2_ASAP7_75t_L g16260 ( 
.A(n_15870),
.B(n_8695),
.Y(n_16260)
);

NAND2xp5_ASAP7_75t_L g16261 ( 
.A(n_15649),
.B(n_9838),
.Y(n_16261)
);

NAND2xp5_ASAP7_75t_L g16262 ( 
.A(n_15608),
.B(n_9842),
.Y(n_16262)
);

OR2x2_ASAP7_75t_L g16263 ( 
.A(n_15632),
.B(n_8710),
.Y(n_16263)
);

NOR2x1_ASAP7_75t_L g16264 ( 
.A(n_15971),
.B(n_11385),
.Y(n_16264)
);

NAND3xp33_ASAP7_75t_L g16265 ( 
.A(n_15826),
.B(n_11505),
.C(n_8161),
.Y(n_16265)
);

INVx4_ASAP7_75t_L g16266 ( 
.A(n_16052),
.Y(n_16266)
);

INVx1_ASAP7_75t_L g16267 ( 
.A(n_15617),
.Y(n_16267)
);

INVxp67_ASAP7_75t_L g16268 ( 
.A(n_15913),
.Y(n_16268)
);

AND2x2_ASAP7_75t_L g16269 ( 
.A(n_15951),
.B(n_11110),
.Y(n_16269)
);

NAND2xp33_ASAP7_75t_SL g16270 ( 
.A(n_15805),
.B(n_7182),
.Y(n_16270)
);

OR2x6_ASAP7_75t_L g16271 ( 
.A(n_15825),
.B(n_8802),
.Y(n_16271)
);

NAND2xp5_ASAP7_75t_L g16272 ( 
.A(n_15762),
.B(n_15668),
.Y(n_16272)
);

NAND2xp5_ASAP7_75t_L g16273 ( 
.A(n_15583),
.B(n_9842),
.Y(n_16273)
);

INVxp67_ASAP7_75t_SL g16274 ( 
.A(n_15622),
.Y(n_16274)
);

INVxp67_ASAP7_75t_L g16275 ( 
.A(n_15930),
.Y(n_16275)
);

NOR2x1_ASAP7_75t_L g16276 ( 
.A(n_16007),
.B(n_9134),
.Y(n_16276)
);

OAI21xp5_ASAP7_75t_L g16277 ( 
.A1(n_15701),
.A2(n_10587),
.B(n_10585),
.Y(n_16277)
);

OAI21xp33_ASAP7_75t_L g16278 ( 
.A1(n_15966),
.A2(n_10909),
.B(n_10889),
.Y(n_16278)
);

INVx2_ASAP7_75t_L g16279 ( 
.A(n_15639),
.Y(n_16279)
);

OR2x2_ASAP7_75t_L g16280 ( 
.A(n_15550),
.B(n_8710),
.Y(n_16280)
);

NAND2xp5_ASAP7_75t_L g16281 ( 
.A(n_15952),
.B(n_9843),
.Y(n_16281)
);

AND2x2_ASAP7_75t_L g16282 ( 
.A(n_15846),
.B(n_9964),
.Y(n_16282)
);

INVx1_ASAP7_75t_L g16283 ( 
.A(n_15587),
.Y(n_16283)
);

NAND4xp25_ASAP7_75t_L g16284 ( 
.A(n_15972),
.B(n_7903),
.C(n_7933),
.D(n_7823),
.Y(n_16284)
);

AND2x2_ASAP7_75t_L g16285 ( 
.A(n_15967),
.B(n_9975),
.Y(n_16285)
);

NAND2xp5_ASAP7_75t_L g16286 ( 
.A(n_15978),
.B(n_15817),
.Y(n_16286)
);

NOR2xp33_ASAP7_75t_L g16287 ( 
.A(n_15944),
.B(n_9975),
.Y(n_16287)
);

NAND2xp5_ASAP7_75t_L g16288 ( 
.A(n_15821),
.B(n_9843),
.Y(n_16288)
);

NAND2xp5_ASAP7_75t_L g16289 ( 
.A(n_15664),
.B(n_9852),
.Y(n_16289)
);

AND2x2_ASAP7_75t_L g16290 ( 
.A(n_15591),
.B(n_9975),
.Y(n_16290)
);

NAND2xp5_ASAP7_75t_L g16291 ( 
.A(n_15881),
.B(n_9852),
.Y(n_16291)
);

NAND2x1_ASAP7_75t_L g16292 ( 
.A(n_15958),
.B(n_8431),
.Y(n_16292)
);

NAND2xp5_ASAP7_75t_L g16293 ( 
.A(n_15742),
.B(n_9855),
.Y(n_16293)
);

INVx2_ASAP7_75t_L g16294 ( 
.A(n_15745),
.Y(n_16294)
);

AND2x2_ASAP7_75t_L g16295 ( 
.A(n_15597),
.B(n_9982),
.Y(n_16295)
);

NAND2xp5_ASAP7_75t_L g16296 ( 
.A(n_15898),
.B(n_9855),
.Y(n_16296)
);

INVx1_ASAP7_75t_L g16297 ( 
.A(n_15607),
.Y(n_16297)
);

AND2x4_ASAP7_75t_L g16298 ( 
.A(n_15609),
.B(n_8592),
.Y(n_16298)
);

NAND2xp5_ASAP7_75t_L g16299 ( 
.A(n_15918),
.B(n_9857),
.Y(n_16299)
);

NAND2xp5_ASAP7_75t_L g16300 ( 
.A(n_15973),
.B(n_9857),
.Y(n_16300)
);

INVx3_ASAP7_75t_L g16301 ( 
.A(n_15861),
.Y(n_16301)
);

INVx1_ASAP7_75t_L g16302 ( 
.A(n_15626),
.Y(n_16302)
);

OR2x2_ASAP7_75t_L g16303 ( 
.A(n_15759),
.B(n_8714),
.Y(n_16303)
);

AO21x2_ASAP7_75t_L g16304 ( 
.A1(n_15563),
.A2(n_10594),
.B(n_10587),
.Y(n_16304)
);

INVx2_ASAP7_75t_L g16305 ( 
.A(n_15669),
.Y(n_16305)
);

INVx2_ASAP7_75t_L g16306 ( 
.A(n_15641),
.Y(n_16306)
);

OR2x2_ASAP7_75t_L g16307 ( 
.A(n_15786),
.B(n_8714),
.Y(n_16307)
);

INVx2_ASAP7_75t_L g16308 ( 
.A(n_15689),
.Y(n_16308)
);

HB1xp67_ASAP7_75t_L g16309 ( 
.A(n_15878),
.Y(n_16309)
);

INVx1_ASAP7_75t_L g16310 ( 
.A(n_15613),
.Y(n_16310)
);

NAND2xp5_ASAP7_75t_L g16311 ( 
.A(n_15695),
.B(n_9861),
.Y(n_16311)
);

AND2x2_ASAP7_75t_L g16312 ( 
.A(n_16047),
.B(n_9982),
.Y(n_16312)
);

INVx1_ASAP7_75t_L g16313 ( 
.A(n_15605),
.Y(n_16313)
);

HB1xp67_ASAP7_75t_L g16314 ( 
.A(n_15980),
.Y(n_16314)
);

AND2x2_ASAP7_75t_L g16315 ( 
.A(n_15996),
.B(n_9982),
.Y(n_16315)
);

NAND2xp5_ASAP7_75t_L g16316 ( 
.A(n_15984),
.B(n_9861),
.Y(n_16316)
);

INVx2_ASAP7_75t_L g16317 ( 
.A(n_15798),
.Y(n_16317)
);

INVx1_ASAP7_75t_L g16318 ( 
.A(n_15847),
.Y(n_16318)
);

OR2x2_ASAP7_75t_L g16319 ( 
.A(n_15612),
.B(n_8727),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_15764),
.B(n_9988),
.Y(n_16320)
);

AND2x2_ASAP7_75t_L g16321 ( 
.A(n_15852),
.B(n_9988),
.Y(n_16321)
);

OR2x2_ASAP7_75t_L g16322 ( 
.A(n_15749),
.B(n_8727),
.Y(n_16322)
);

INVx1_ASAP7_75t_L g16323 ( 
.A(n_15690),
.Y(n_16323)
);

INVx2_ASAP7_75t_L g16324 ( 
.A(n_15643),
.Y(n_16324)
);

INVx1_ASAP7_75t_L g16325 ( 
.A(n_15712),
.Y(n_16325)
);

AND2x2_ASAP7_75t_L g16326 ( 
.A(n_15636),
.B(n_15771),
.Y(n_16326)
);

AND2x2_ASAP7_75t_L g16327 ( 
.A(n_15772),
.B(n_15698),
.Y(n_16327)
);

INVx2_ASAP7_75t_L g16328 ( 
.A(n_15814),
.Y(n_16328)
);

NAND2xp5_ASAP7_75t_L g16329 ( 
.A(n_15919),
.B(n_9865),
.Y(n_16329)
);

AND2x2_ASAP7_75t_L g16330 ( 
.A(n_15840),
.B(n_9988),
.Y(n_16330)
);

INVx1_ASAP7_75t_L g16331 ( 
.A(n_15714),
.Y(n_16331)
);

AOI22xp33_ASAP7_75t_SL g16332 ( 
.A1(n_15985),
.A2(n_8483),
.B1(n_8494),
.B2(n_8340),
.Y(n_16332)
);

CKINVDCx5p33_ASAP7_75t_R g16333 ( 
.A(n_15845),
.Y(n_16333)
);

INVx1_ASAP7_75t_SL g16334 ( 
.A(n_15740),
.Y(n_16334)
);

AND2x6_ASAP7_75t_L g16335 ( 
.A(n_15750),
.B(n_8483),
.Y(n_16335)
);

INVx1_ASAP7_75t_L g16336 ( 
.A(n_15752),
.Y(n_16336)
);

INVx1_ASAP7_75t_L g16337 ( 
.A(n_15755),
.Y(n_16337)
);

AND2x2_ASAP7_75t_L g16338 ( 
.A(n_15754),
.B(n_15715),
.Y(n_16338)
);

INVx4_ASAP7_75t_L g16339 ( 
.A(n_15735),
.Y(n_16339)
);

INVx1_ASAP7_75t_L g16340 ( 
.A(n_15659),
.Y(n_16340)
);

OR2x2_ASAP7_75t_L g16341 ( 
.A(n_15787),
.B(n_8769),
.Y(n_16341)
);

INVx1_ASAP7_75t_L g16342 ( 
.A(n_15655),
.Y(n_16342)
);

NAND4xp25_ASAP7_75t_SL g16343 ( 
.A(n_15873),
.B(n_9264),
.C(n_9269),
.D(n_9257),
.Y(n_16343)
);

INVx2_ASAP7_75t_L g16344 ( 
.A(n_15741),
.Y(n_16344)
);

AOI22xp5_ASAP7_75t_L g16345 ( 
.A1(n_15711),
.A2(n_8494),
.B1(n_8526),
.B2(n_8483),
.Y(n_16345)
);

NOR2xp33_ASAP7_75t_L g16346 ( 
.A(n_15779),
.B(n_9991),
.Y(n_16346)
);

AND2x2_ASAP7_75t_L g16347 ( 
.A(n_15781),
.B(n_9991),
.Y(n_16347)
);

INVxp67_ASAP7_75t_SL g16348 ( 
.A(n_15666),
.Y(n_16348)
);

NAND3xp33_ASAP7_75t_L g16349 ( 
.A(n_15819),
.B(n_8161),
.C(n_8156),
.Y(n_16349)
);

INVx1_ASAP7_75t_L g16350 ( 
.A(n_15638),
.Y(n_16350)
);

NAND2xp5_ASAP7_75t_L g16351 ( 
.A(n_15791),
.B(n_9865),
.Y(n_16351)
);

NOR2xp67_ASAP7_75t_L g16352 ( 
.A(n_15761),
.B(n_9991),
.Y(n_16352)
);

INVx2_ASAP7_75t_L g16353 ( 
.A(n_15777),
.Y(n_16353)
);

AND2x2_ASAP7_75t_L g16354 ( 
.A(n_15783),
.B(n_10002),
.Y(n_16354)
);

INVx1_ASAP7_75t_L g16355 ( 
.A(n_15623),
.Y(n_16355)
);

INVx1_ASAP7_75t_L g16356 ( 
.A(n_15627),
.Y(n_16356)
);

AND2x2_ASAP7_75t_L g16357 ( 
.A(n_15802),
.B(n_10002),
.Y(n_16357)
);

HB1xp67_ASAP7_75t_L g16358 ( 
.A(n_15812),
.Y(n_16358)
);

OAI21xp33_ASAP7_75t_L g16359 ( 
.A1(n_15720),
.A2(n_10909),
.B(n_10594),
.Y(n_16359)
);

INVx3_ASAP7_75t_L g16360 ( 
.A(n_15911),
.Y(n_16360)
);

OR2x2_ASAP7_75t_L g16361 ( 
.A(n_15792),
.B(n_15718),
.Y(n_16361)
);

OR2x2_ASAP7_75t_L g16362 ( 
.A(n_16003),
.B(n_15637),
.Y(n_16362)
);

INVx1_ASAP7_75t_L g16363 ( 
.A(n_15716),
.Y(n_16363)
);

AND2x4_ASAP7_75t_L g16364 ( 
.A(n_15920),
.B(n_8700),
.Y(n_16364)
);

NAND2xp5_ASAP7_75t_SL g16365 ( 
.A(n_15797),
.B(n_8483),
.Y(n_16365)
);

NAND2xp5_ASAP7_75t_L g16366 ( 
.A(n_16029),
.B(n_9867),
.Y(n_16366)
);

OR2x2_ASAP7_75t_L g16367 ( 
.A(n_16057),
.B(n_8769),
.Y(n_16367)
);

INVxp67_ASAP7_75t_L g16368 ( 
.A(n_15803),
.Y(n_16368)
);

BUFx3_ASAP7_75t_L g16369 ( 
.A(n_16032),
.Y(n_16369)
);

INVx1_ASAP7_75t_L g16370 ( 
.A(n_15644),
.Y(n_16370)
);

INVx2_ASAP7_75t_L g16371 ( 
.A(n_15744),
.Y(n_16371)
);

AND2x2_ASAP7_75t_L g16372 ( 
.A(n_15806),
.B(n_15837),
.Y(n_16372)
);

INVx1_ASAP7_75t_L g16373 ( 
.A(n_15678),
.Y(n_16373)
);

NAND2xp5_ASAP7_75t_L g16374 ( 
.A(n_16037),
.B(n_9867),
.Y(n_16374)
);

NAND2xp5_ASAP7_75t_L g16375 ( 
.A(n_16040),
.B(n_9870),
.Y(n_16375)
);

NOR2xp33_ASAP7_75t_L g16376 ( 
.A(n_15544),
.B(n_16044),
.Y(n_16376)
);

NAND2xp5_ASAP7_75t_L g16377 ( 
.A(n_16050),
.B(n_9870),
.Y(n_16377)
);

AND2x2_ASAP7_75t_L g16378 ( 
.A(n_15739),
.B(n_10002),
.Y(n_16378)
);

NAND2xp5_ASAP7_75t_L g16379 ( 
.A(n_16055),
.B(n_9871),
.Y(n_16379)
);

NAND2xp5_ASAP7_75t_L g16380 ( 
.A(n_15915),
.B(n_15839),
.Y(n_16380)
);

AND2x2_ASAP7_75t_SL g16381 ( 
.A(n_15723),
.B(n_15879),
.Y(n_16381)
);

INVx1_ASAP7_75t_L g16382 ( 
.A(n_15697),
.Y(n_16382)
);

CKINVDCx16_ASAP7_75t_R g16383 ( 
.A(n_15925),
.Y(n_16383)
);

HB1xp67_ASAP7_75t_L g16384 ( 
.A(n_15692),
.Y(n_16384)
);

O2A1O1Ixp33_ASAP7_75t_SL g16385 ( 
.A1(n_15886),
.A2(n_7978),
.B(n_8021),
.C(n_7908),
.Y(n_16385)
);

AND2x2_ASAP7_75t_L g16386 ( 
.A(n_15670),
.B(n_10017),
.Y(n_16386)
);

NOR2xp33_ASAP7_75t_L g16387 ( 
.A(n_15893),
.B(n_10017),
.Y(n_16387)
);

NAND2xp5_ASAP7_75t_L g16388 ( 
.A(n_15721),
.B(n_9871),
.Y(n_16388)
);

INVx1_ASAP7_75t_L g16389 ( 
.A(n_15776),
.Y(n_16389)
);

INVx1_ASAP7_75t_L g16390 ( 
.A(n_15794),
.Y(n_16390)
);

OR2x2_ASAP7_75t_L g16391 ( 
.A(n_15947),
.B(n_8775),
.Y(n_16391)
);

INVx2_ASAP7_75t_L g16392 ( 
.A(n_15651),
.Y(n_16392)
);

AND2x4_ASAP7_75t_L g16393 ( 
.A(n_15902),
.B(n_8700),
.Y(n_16393)
);

INVx1_ASAP7_75t_L g16394 ( 
.A(n_15653),
.Y(n_16394)
);

NAND2xp33_ASAP7_75t_SL g16395 ( 
.A(n_15685),
.B(n_8483),
.Y(n_16395)
);

AND2x2_ASAP7_75t_L g16396 ( 
.A(n_15675),
.B(n_10017),
.Y(n_16396)
);

AND2x2_ASAP7_75t_L g16397 ( 
.A(n_15848),
.B(n_10022),
.Y(n_16397)
);

AND2x2_ASAP7_75t_L g16398 ( 
.A(n_15680),
.B(n_10022),
.Y(n_16398)
);

AND2x2_ASAP7_75t_L g16399 ( 
.A(n_15682),
.B(n_10022),
.Y(n_16399)
);

NAND2xp5_ASAP7_75t_L g16400 ( 
.A(n_15751),
.B(n_9872),
.Y(n_16400)
);

INVx1_ASAP7_75t_L g16401 ( 
.A(n_15820),
.Y(n_16401)
);

AOI21xp5_ASAP7_75t_L g16402 ( 
.A1(n_15987),
.A2(n_9280),
.B(n_9269),
.Y(n_16402)
);

AND2x2_ASAP7_75t_L g16403 ( 
.A(n_15684),
.B(n_10025),
.Y(n_16403)
);

AOI221xp5_ASAP7_75t_L g16404 ( 
.A1(n_15725),
.A2(n_9284),
.B1(n_9286),
.B2(n_9280),
.C(n_9269),
.Y(n_16404)
);

OAI211xp5_ASAP7_75t_SL g16405 ( 
.A1(n_15991),
.A2(n_9284),
.B(n_9286),
.C(n_9280),
.Y(n_16405)
);

INVx2_ASAP7_75t_L g16406 ( 
.A(n_15940),
.Y(n_16406)
);

INVx1_ASAP7_75t_L g16407 ( 
.A(n_15811),
.Y(n_16407)
);

AND2x2_ASAP7_75t_L g16408 ( 
.A(n_15888),
.B(n_10025),
.Y(n_16408)
);

AOI21xp33_ASAP7_75t_SL g16409 ( 
.A1(n_15838),
.A2(n_11422),
.B(n_11416),
.Y(n_16409)
);

NAND2xp5_ASAP7_75t_L g16410 ( 
.A(n_15842),
.B(n_15747),
.Y(n_16410)
);

BUFx2_ASAP7_75t_L g16411 ( 
.A(n_15808),
.Y(n_16411)
);

AND2x2_ASAP7_75t_L g16412 ( 
.A(n_15962),
.B(n_10025),
.Y(n_16412)
);

AND2x4_ASAP7_75t_SL g16413 ( 
.A(n_15707),
.B(n_7042),
.Y(n_16413)
);

INVx1_ASAP7_75t_L g16414 ( 
.A(n_15858),
.Y(n_16414)
);

AND2x2_ASAP7_75t_L g16415 ( 
.A(n_15965),
.B(n_10027),
.Y(n_16415)
);

OR2x6_ASAP7_75t_L g16416 ( 
.A(n_15963),
.B(n_15872),
.Y(n_16416)
);

INVx1_ASAP7_75t_L g16417 ( 
.A(n_15867),
.Y(n_16417)
);

NAND2xp5_ASAP7_75t_L g16418 ( 
.A(n_15862),
.B(n_9872),
.Y(n_16418)
);

NAND2xp5_ASAP7_75t_L g16419 ( 
.A(n_15863),
.B(n_9875),
.Y(n_16419)
);

AND2x2_ASAP7_75t_SL g16420 ( 
.A(n_15667),
.B(n_8483),
.Y(n_16420)
);

INVx2_ASAP7_75t_L g16421 ( 
.A(n_15929),
.Y(n_16421)
);

NAND4xp25_ASAP7_75t_L g16422 ( 
.A(n_15642),
.B(n_7933),
.C(n_7961),
.D(n_7903),
.Y(n_16422)
);

INVx1_ASAP7_75t_L g16423 ( 
.A(n_15790),
.Y(n_16423)
);

OR2x2_ASAP7_75t_L g16424 ( 
.A(n_15672),
.B(n_8775),
.Y(n_16424)
);

AND2x2_ASAP7_75t_L g16425 ( 
.A(n_15993),
.B(n_10027),
.Y(n_16425)
);

AND2x2_ASAP7_75t_L g16426 ( 
.A(n_15921),
.B(n_10027),
.Y(n_16426)
);

NAND2x1_ASAP7_75t_L g16427 ( 
.A(n_16012),
.B(n_8431),
.Y(n_16427)
);

INVx2_ASAP7_75t_L g16428 ( 
.A(n_15992),
.Y(n_16428)
);

NAND2xp5_ASAP7_75t_L g16429 ( 
.A(n_15874),
.B(n_9875),
.Y(n_16429)
);

INVx1_ASAP7_75t_L g16430 ( 
.A(n_15710),
.Y(n_16430)
);

OR2x6_ASAP7_75t_L g16431 ( 
.A(n_15875),
.B(n_6965),
.Y(n_16431)
);

NAND2xp5_ASAP7_75t_L g16432 ( 
.A(n_15869),
.B(n_9876),
.Y(n_16432)
);

OR2x2_ASAP7_75t_L g16433 ( 
.A(n_15673),
.B(n_8795),
.Y(n_16433)
);

NAND2xp5_ASAP7_75t_SL g16434 ( 
.A(n_15922),
.B(n_8483),
.Y(n_16434)
);

AND2x2_ASAP7_75t_L g16435 ( 
.A(n_15936),
.B(n_16020),
.Y(n_16435)
);

AND2x2_ASAP7_75t_L g16436 ( 
.A(n_15827),
.B(n_10041),
.Y(n_16436)
);

INVx4_ASAP7_75t_L g16437 ( 
.A(n_15835),
.Y(n_16437)
);

AND2x2_ASAP7_75t_L g16438 ( 
.A(n_16027),
.B(n_10041),
.Y(n_16438)
);

INVx2_ASAP7_75t_L g16439 ( 
.A(n_15851),
.Y(n_16439)
);

INVx1_ASAP7_75t_L g16440 ( 
.A(n_15800),
.Y(n_16440)
);

INVx2_ASAP7_75t_L g16441 ( 
.A(n_15927),
.Y(n_16441)
);

BUFx2_ASAP7_75t_L g16442 ( 
.A(n_15850),
.Y(n_16442)
);

AOI221xp5_ASAP7_75t_L g16443 ( 
.A1(n_15997),
.A2(n_9292),
.B1(n_9298),
.B2(n_9286),
.C(n_9284),
.Y(n_16443)
);

AND2x4_ASAP7_75t_L g16444 ( 
.A(n_16028),
.B(n_8700),
.Y(n_16444)
);

OAI211xp5_ASAP7_75t_SL g16445 ( 
.A1(n_15950),
.A2(n_9298),
.B(n_9300),
.C(n_9292),
.Y(n_16445)
);

INVx2_ASAP7_75t_L g16446 ( 
.A(n_15953),
.Y(n_16446)
);

NAND2xp5_ASAP7_75t_L g16447 ( 
.A(n_15876),
.B(n_9876),
.Y(n_16447)
);

INVx1_ASAP7_75t_L g16448 ( 
.A(n_15885),
.Y(n_16448)
);

AND2x2_ASAP7_75t_L g16449 ( 
.A(n_16022),
.B(n_10041),
.Y(n_16449)
);

AND2x2_ASAP7_75t_L g16450 ( 
.A(n_15907),
.B(n_10049),
.Y(n_16450)
);

BUFx2_ASAP7_75t_L g16451 ( 
.A(n_15877),
.Y(n_16451)
);

NAND2xp5_ASAP7_75t_L g16452 ( 
.A(n_15906),
.B(n_15880),
.Y(n_16452)
);

INVx1_ASAP7_75t_SL g16453 ( 
.A(n_15829),
.Y(n_16453)
);

NAND2xp5_ASAP7_75t_L g16454 ( 
.A(n_15882),
.B(n_15699),
.Y(n_16454)
);

INVx4_ASAP7_75t_L g16455 ( 
.A(n_15935),
.Y(n_16455)
);

OR2x2_ASAP7_75t_L g16456 ( 
.A(n_15964),
.B(n_8795),
.Y(n_16456)
);

INVx4_ASAP7_75t_SL g16457 ( 
.A(n_15968),
.Y(n_16457)
);

AND2x2_ASAP7_75t_L g16458 ( 
.A(n_15994),
.B(n_10049),
.Y(n_16458)
);

INVx1_ASAP7_75t_SL g16459 ( 
.A(n_15815),
.Y(n_16459)
);

INVx2_ASAP7_75t_SL g16460 ( 
.A(n_16001),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_15959),
.Y(n_16461)
);

NAND2xp5_ASAP7_75t_L g16462 ( 
.A(n_15702),
.B(n_9879),
.Y(n_16462)
);

OR2x2_ASAP7_75t_L g16463 ( 
.A(n_15990),
.B(n_8803),
.Y(n_16463)
);

AND2x2_ASAP7_75t_L g16464 ( 
.A(n_16002),
.B(n_10049),
.Y(n_16464)
);

NAND2xp33_ASAP7_75t_SL g16465 ( 
.A(n_15828),
.B(n_8494),
.Y(n_16465)
);

CKINVDCx16_ASAP7_75t_R g16466 ( 
.A(n_16006),
.Y(n_16466)
);

INVx1_ASAP7_75t_L g16467 ( 
.A(n_15753),
.Y(n_16467)
);

INVx1_ASAP7_75t_L g16468 ( 
.A(n_15768),
.Y(n_16468)
);

AOI221xp5_ASAP7_75t_L g16469 ( 
.A1(n_15975),
.A2(n_9300),
.B1(n_9304),
.B2(n_9298),
.C(n_9292),
.Y(n_16469)
);

AND2x2_ASAP7_75t_L g16470 ( 
.A(n_16009),
.B(n_10060),
.Y(n_16470)
);

INVx1_ASAP7_75t_L g16471 ( 
.A(n_15728),
.Y(n_16471)
);

OA21x2_ASAP7_75t_L g16472 ( 
.A1(n_15799),
.A2(n_11422),
.B(n_11416),
.Y(n_16472)
);

HB1xp67_ASAP7_75t_L g16473 ( 
.A(n_15836),
.Y(n_16473)
);

INVx5_ASAP7_75t_L g16474 ( 
.A(n_15941),
.Y(n_16474)
);

INVx1_ASAP7_75t_L g16475 ( 
.A(n_15942),
.Y(n_16475)
);

INVx1_ASAP7_75t_L g16476 ( 
.A(n_15679),
.Y(n_16476)
);

AND2x2_ASAP7_75t_L g16477 ( 
.A(n_16014),
.B(n_10060),
.Y(n_16477)
);

INVx1_ASAP7_75t_L g16478 ( 
.A(n_15769),
.Y(n_16478)
);

AND2x4_ASAP7_75t_L g16479 ( 
.A(n_16016),
.B(n_8700),
.Y(n_16479)
);

OR2x2_ASAP7_75t_L g16480 ( 
.A(n_15871),
.B(n_8803),
.Y(n_16480)
);

AND2x2_ASAP7_75t_L g16481 ( 
.A(n_15775),
.B(n_10060),
.Y(n_16481)
);

AND2x2_ASAP7_75t_L g16482 ( 
.A(n_15780),
.B(n_10073),
.Y(n_16482)
);

INVx2_ASAP7_75t_L g16483 ( 
.A(n_15957),
.Y(n_16483)
);

INVx1_ASAP7_75t_L g16484 ( 
.A(n_15782),
.Y(n_16484)
);

NOR2xp67_ASAP7_75t_L g16485 ( 
.A(n_15765),
.B(n_10073),
.Y(n_16485)
);

AND2x2_ASAP7_75t_L g16486 ( 
.A(n_15908),
.B(n_10073),
.Y(n_16486)
);

NAND2xp5_ASAP7_75t_L g16487 ( 
.A(n_15865),
.B(n_9879),
.Y(n_16487)
);

INVx1_ASAP7_75t_L g16488 ( 
.A(n_15773),
.Y(n_16488)
);

AND2x2_ASAP7_75t_L g16489 ( 
.A(n_15924),
.B(n_10074),
.Y(n_16489)
);

NAND2x1p5_ASAP7_75t_L g16490 ( 
.A(n_15788),
.B(n_15804),
.Y(n_16490)
);

INVx2_ASAP7_75t_L g16491 ( 
.A(n_15969),
.Y(n_16491)
);

INVxp67_ASAP7_75t_SL g16492 ( 
.A(n_15887),
.Y(n_16492)
);

OR2x2_ASAP7_75t_L g16493 ( 
.A(n_15853),
.B(n_8594),
.Y(n_16493)
);

AND2x2_ASAP7_75t_L g16494 ( 
.A(n_15926),
.B(n_15889),
.Y(n_16494)
);

NAND2xp5_ASAP7_75t_L g16495 ( 
.A(n_15986),
.B(n_9881),
.Y(n_16495)
);

INVx1_ASAP7_75t_L g16496 ( 
.A(n_15729),
.Y(n_16496)
);

AND2x2_ASAP7_75t_L g16497 ( 
.A(n_15832),
.B(n_10074),
.Y(n_16497)
);

AND2x2_ASAP7_75t_L g16498 ( 
.A(n_15998),
.B(n_10074),
.Y(n_16498)
);

INVx1_ASAP7_75t_L g16499 ( 
.A(n_15731),
.Y(n_16499)
);

NOR3xp33_ASAP7_75t_SL g16500 ( 
.A(n_15704),
.B(n_8556),
.C(n_8552),
.Y(n_16500)
);

OAI221xp5_ASAP7_75t_L g16501 ( 
.A1(n_15860),
.A2(n_9312),
.B1(n_9319),
.B2(n_9304),
.C(n_9300),
.Y(n_16501)
);

NAND2xp5_ASAP7_75t_L g16502 ( 
.A(n_15796),
.B(n_9881),
.Y(n_16502)
);

AND2x4_ASAP7_75t_L g16503 ( 
.A(n_15801),
.B(n_8700),
.Y(n_16503)
);

NAND2xp5_ASAP7_75t_L g16504 ( 
.A(n_16005),
.B(n_9885),
.Y(n_16504)
);

NOR2xp33_ASAP7_75t_SL g16505 ( 
.A(n_15807),
.B(n_8494),
.Y(n_16505)
);

AND2x2_ASAP7_75t_L g16506 ( 
.A(n_15912),
.B(n_10075),
.Y(n_16506)
);

AND2x2_ASAP7_75t_L g16507 ( 
.A(n_16010),
.B(n_10075),
.Y(n_16507)
);

AND2x2_ASAP7_75t_SL g16508 ( 
.A(n_15831),
.B(n_15833),
.Y(n_16508)
);

NAND2xp5_ASAP7_75t_L g16509 ( 
.A(n_16011),
.B(n_16013),
.Y(n_16509)
);

OR2x2_ASAP7_75t_L g16510 ( 
.A(n_15983),
.B(n_8594),
.Y(n_16510)
);

INVx1_ASAP7_75t_L g16511 ( 
.A(n_15895),
.Y(n_16511)
);

AND2x2_ASAP7_75t_L g16512 ( 
.A(n_16023),
.B(n_10075),
.Y(n_16512)
);

AND2x2_ASAP7_75t_L g16513 ( 
.A(n_16024),
.B(n_10077),
.Y(n_16513)
);

AND2x2_ASAP7_75t_L g16514 ( 
.A(n_16043),
.B(n_10077),
.Y(n_16514)
);

AND2x4_ASAP7_75t_L g16515 ( 
.A(n_15892),
.B(n_8717),
.Y(n_16515)
);

NAND2xp5_ASAP7_75t_SL g16516 ( 
.A(n_15933),
.B(n_16054),
.Y(n_16516)
);

AND2x2_ASAP7_75t_L g16517 ( 
.A(n_16048),
.B(n_10077),
.Y(n_16517)
);

INVx1_ASAP7_75t_L g16518 ( 
.A(n_15894),
.Y(n_16518)
);

INVx1_ASAP7_75t_L g16519 ( 
.A(n_15900),
.Y(n_16519)
);

INVx1_ASAP7_75t_L g16520 ( 
.A(n_15909),
.Y(n_16520)
);

OR2x2_ASAP7_75t_L g16521 ( 
.A(n_15954),
.B(n_15955),
.Y(n_16521)
);

NAND2xp5_ASAP7_75t_SL g16522 ( 
.A(n_15933),
.B(n_8494),
.Y(n_16522)
);

AND2x2_ASAP7_75t_L g16523 ( 
.A(n_16051),
.B(n_10084),
.Y(n_16523)
);

AND2x2_ASAP7_75t_L g16524 ( 
.A(n_15970),
.B(n_10084),
.Y(n_16524)
);

BUFx3_ASAP7_75t_L g16525 ( 
.A(n_15849),
.Y(n_16525)
);

INVx2_ASAP7_75t_L g16526 ( 
.A(n_15982),
.Y(n_16526)
);

AND2x2_ASAP7_75t_L g16527 ( 
.A(n_16004),
.B(n_10084),
.Y(n_16527)
);

INVx1_ASAP7_75t_L g16528 ( 
.A(n_15916),
.Y(n_16528)
);

HB1xp67_ASAP7_75t_L g16529 ( 
.A(n_16034),
.Y(n_16529)
);

NAND2xp5_ASAP7_75t_L g16530 ( 
.A(n_15981),
.B(n_9885),
.Y(n_16530)
);

INVx2_ASAP7_75t_L g16531 ( 
.A(n_16049),
.Y(n_16531)
);

INVx1_ASAP7_75t_L g16532 ( 
.A(n_15917),
.Y(n_16532)
);

OR2x2_ASAP7_75t_L g16533 ( 
.A(n_15931),
.B(n_8845),
.Y(n_16533)
);

AND3x2_ASAP7_75t_L g16534 ( 
.A(n_15995),
.B(n_6906),
.C(n_6852),
.Y(n_16534)
);

INVx1_ASAP7_75t_L g16535 ( 
.A(n_15854),
.Y(n_16535)
);

INVx1_ASAP7_75t_L g16536 ( 
.A(n_15856),
.Y(n_16536)
);

AND2x2_ASAP7_75t_L g16537 ( 
.A(n_15868),
.B(n_10107),
.Y(n_16537)
);

INVx1_ASAP7_75t_L g16538 ( 
.A(n_15903),
.Y(n_16538)
);

OR2x6_ASAP7_75t_L g16539 ( 
.A(n_15934),
.B(n_6965),
.Y(n_16539)
);

INVx1_ASAP7_75t_L g16540 ( 
.A(n_15938),
.Y(n_16540)
);

NOR2x1_ASAP7_75t_R g16541 ( 
.A(n_15939),
.B(n_7139),
.Y(n_16541)
);

INVx1_ASAP7_75t_L g16542 ( 
.A(n_15961),
.Y(n_16542)
);

INVx2_ASAP7_75t_L g16543 ( 
.A(n_16019),
.Y(n_16543)
);

INVx1_ASAP7_75t_L g16544 ( 
.A(n_15979),
.Y(n_16544)
);

NOR2xp33_ASAP7_75t_L g16545 ( 
.A(n_15923),
.B(n_15988),
.Y(n_16545)
);

INVx2_ASAP7_75t_L g16546 ( 
.A(n_16025),
.Y(n_16546)
);

INVx1_ASAP7_75t_L g16547 ( 
.A(n_15974),
.Y(n_16547)
);

AND2x2_ASAP7_75t_L g16548 ( 
.A(n_15999),
.B(n_10107),
.Y(n_16548)
);

AND2x6_ASAP7_75t_SL g16549 ( 
.A(n_16018),
.B(n_8852),
.Y(n_16549)
);

INVx1_ASAP7_75t_L g16550 ( 
.A(n_16031),
.Y(n_16550)
);

AND2x2_ASAP7_75t_L g16551 ( 
.A(n_16036),
.B(n_10107),
.Y(n_16551)
);

OR2x2_ASAP7_75t_L g16552 ( 
.A(n_16046),
.B(n_8845),
.Y(n_16552)
);

AND2x2_ASAP7_75t_L g16553 ( 
.A(n_16053),
.B(n_10115),
.Y(n_16553)
);

NAND3x1_ASAP7_75t_L g16554 ( 
.A(n_15676),
.B(n_10280),
.C(n_10189),
.Y(n_16554)
);

INVx2_ASAP7_75t_L g16555 ( 
.A(n_16030),
.Y(n_16555)
);

NAND4xp25_ASAP7_75t_L g16556 ( 
.A(n_16026),
.B(n_7933),
.C(n_7961),
.D(n_7903),
.Y(n_16556)
);

INVx1_ASAP7_75t_L g16557 ( 
.A(n_16033),
.Y(n_16557)
);

INVx2_ASAP7_75t_L g16558 ( 
.A(n_15977),
.Y(n_16558)
);

NOR2x1_ASAP7_75t_L g16559 ( 
.A(n_15946),
.B(n_9901),
.Y(n_16559)
);

AND2x2_ASAP7_75t_L g16560 ( 
.A(n_16045),
.B(n_10115),
.Y(n_16560)
);

HB1xp67_ASAP7_75t_L g16561 ( 
.A(n_15645),
.Y(n_16561)
);

NAND2xp5_ASAP7_75t_L g16562 ( 
.A(n_16077),
.B(n_15717),
.Y(n_16562)
);

OAI33xp33_ASAP7_75t_L g16563 ( 
.A1(n_16078),
.A2(n_16083),
.A3(n_16060),
.B1(n_16073),
.B2(n_16074),
.B3(n_16124),
.Y(n_16563)
);

INVx1_ASAP7_75t_L g16564 ( 
.A(n_16156),
.Y(n_16564)
);

INVx2_ASAP7_75t_L g16565 ( 
.A(n_16099),
.Y(n_16565)
);

NAND2x1_ASAP7_75t_L g16566 ( 
.A(n_16105),
.B(n_10115),
.Y(n_16566)
);

INVx1_ASAP7_75t_L g16567 ( 
.A(n_16059),
.Y(n_16567)
);

NAND2xp5_ASAP7_75t_L g16568 ( 
.A(n_16097),
.B(n_15830),
.Y(n_16568)
);

INVx1_ASAP7_75t_L g16569 ( 
.A(n_16118),
.Y(n_16569)
);

INVx1_ASAP7_75t_L g16570 ( 
.A(n_16120),
.Y(n_16570)
);

OAI322xp33_ASAP7_75t_L g16571 ( 
.A1(n_16376),
.A2(n_9321),
.A3(n_9312),
.B1(n_9319),
.B2(n_9304),
.C1(n_9179),
.C2(n_9175),
.Y(n_16571)
);

OAI22xp5_ASAP7_75t_L g16572 ( 
.A1(n_16072),
.A2(n_16076),
.B1(n_16137),
.B2(n_16268),
.Y(n_16572)
);

AOI22xp5_ASAP7_75t_L g16573 ( 
.A1(n_16070),
.A2(n_8526),
.B1(n_8530),
.B2(n_8494),
.Y(n_16573)
);

INVx1_ASAP7_75t_L g16574 ( 
.A(n_16061),
.Y(n_16574)
);

INVx2_ASAP7_75t_SL g16575 ( 
.A(n_16139),
.Y(n_16575)
);

AOI21xp5_ASAP7_75t_L g16576 ( 
.A1(n_16094),
.A2(n_9319),
.B(n_9312),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_16084),
.Y(n_16577)
);

NAND2x2_ASAP7_75t_L g16578 ( 
.A(n_16141),
.B(n_16066),
.Y(n_16578)
);

AND2x2_ASAP7_75t_L g16579 ( 
.A(n_16089),
.B(n_11467),
.Y(n_16579)
);

INVx1_ASAP7_75t_L g16580 ( 
.A(n_16309),
.Y(n_16580)
);

INVx1_ASAP7_75t_L g16581 ( 
.A(n_16358),
.Y(n_16581)
);

NAND2xp5_ASAP7_75t_L g16582 ( 
.A(n_16192),
.B(n_9901),
.Y(n_16582)
);

OR2x2_ASAP7_75t_L g16583 ( 
.A(n_16179),
.B(n_8574),
.Y(n_16583)
);

NAND2xp5_ASAP7_75t_L g16584 ( 
.A(n_16071),
.B(n_9910),
.Y(n_16584)
);

NAND2xp5_ASAP7_75t_L g16585 ( 
.A(n_16087),
.B(n_9910),
.Y(n_16585)
);

AOI22xp33_ASAP7_75t_L g16586 ( 
.A1(n_16063),
.A2(n_9321),
.B1(n_8526),
.B2(n_8530),
.Y(n_16586)
);

OR2x2_ASAP7_75t_L g16587 ( 
.A(n_16130),
.B(n_8574),
.Y(n_16587)
);

OR2x2_ASAP7_75t_L g16588 ( 
.A(n_16149),
.B(n_8605),
.Y(n_16588)
);

INVx1_ASAP7_75t_L g16589 ( 
.A(n_16474),
.Y(n_16589)
);

INVx1_ASAP7_75t_L g16590 ( 
.A(n_16474),
.Y(n_16590)
);

OAI31xp33_ASAP7_75t_L g16591 ( 
.A1(n_16096),
.A2(n_9321),
.A3(n_8491),
.B(n_8703),
.Y(n_16591)
);

NAND4xp25_ASAP7_75t_L g16592 ( 
.A(n_16143),
.B(n_7933),
.C(n_7961),
.D(n_7903),
.Y(n_16592)
);

INVx1_ASAP7_75t_L g16593 ( 
.A(n_16474),
.Y(n_16593)
);

AOI22xp5_ASAP7_75t_L g16594 ( 
.A1(n_16200),
.A2(n_8526),
.B1(n_8530),
.B2(n_8494),
.Y(n_16594)
);

NOR2xp67_ASAP7_75t_SL g16595 ( 
.A(n_16266),
.B(n_8526),
.Y(n_16595)
);

INVx1_ASAP7_75t_L g16596 ( 
.A(n_16117),
.Y(n_16596)
);

INVxp67_ASAP7_75t_SL g16597 ( 
.A(n_16065),
.Y(n_16597)
);

INVx1_ASAP7_75t_L g16598 ( 
.A(n_16165),
.Y(n_16598)
);

AOI32xp33_ASAP7_75t_L g16599 ( 
.A1(n_16145),
.A2(n_11021),
.A3(n_11025),
.B1(n_10975),
.B2(n_10925),
.Y(n_16599)
);

OR2x2_ASAP7_75t_L g16600 ( 
.A(n_16215),
.B(n_8605),
.Y(n_16600)
);

INVx1_ASAP7_75t_L g16601 ( 
.A(n_16473),
.Y(n_16601)
);

INVx1_ASAP7_75t_L g16602 ( 
.A(n_16116),
.Y(n_16602)
);

INVx2_ASAP7_75t_L g16603 ( 
.A(n_16129),
.Y(n_16603)
);

AND2x2_ASAP7_75t_L g16604 ( 
.A(n_16121),
.B(n_16125),
.Y(n_16604)
);

INVx1_ASAP7_75t_L g16605 ( 
.A(n_16233),
.Y(n_16605)
);

NOR2xp33_ASAP7_75t_SL g16606 ( 
.A(n_16146),
.B(n_8526),
.Y(n_16606)
);

AND2x2_ASAP7_75t_L g16607 ( 
.A(n_16128),
.B(n_11467),
.Y(n_16607)
);

INVx1_ASAP7_75t_L g16608 ( 
.A(n_16158),
.Y(n_16608)
);

NAND2xp5_ASAP7_75t_L g16609 ( 
.A(n_16115),
.B(n_9920),
.Y(n_16609)
);

AND2x4_ASAP7_75t_L g16610 ( 
.A(n_16161),
.B(n_11494),
.Y(n_16610)
);

NAND2xp5_ASAP7_75t_L g16611 ( 
.A(n_16131),
.B(n_9920),
.Y(n_16611)
);

INVxp67_ASAP7_75t_SL g16612 ( 
.A(n_16103),
.Y(n_16612)
);

INVx1_ASAP7_75t_L g16613 ( 
.A(n_16170),
.Y(n_16613)
);

OR2x2_ASAP7_75t_L g16614 ( 
.A(n_16106),
.B(n_8664),
.Y(n_16614)
);

NAND4xp75_ASAP7_75t_SL g16615 ( 
.A(n_16134),
.B(n_10082),
.C(n_10163),
.D(n_10039),
.Y(n_16615)
);

INVxp67_ASAP7_75t_L g16616 ( 
.A(n_16314),
.Y(n_16616)
);

NAND2x2_ASAP7_75t_L g16617 ( 
.A(n_16369),
.B(n_6657),
.Y(n_16617)
);

INVx1_ASAP7_75t_L g16618 ( 
.A(n_16142),
.Y(n_16618)
);

NAND2xp5_ASAP7_75t_L g16619 ( 
.A(n_16140),
.B(n_9922),
.Y(n_16619)
);

NAND2xp5_ASAP7_75t_L g16620 ( 
.A(n_16171),
.B(n_9922),
.Y(n_16620)
);

NAND2x1p5_ASAP7_75t_L g16621 ( 
.A(n_16259),
.B(n_8526),
.Y(n_16621)
);

BUFx2_ASAP7_75t_SL g16622 ( 
.A(n_16069),
.Y(n_16622)
);

CKINVDCx5p33_ASAP7_75t_R g16623 ( 
.A(n_16183),
.Y(n_16623)
);

AND2x4_ASAP7_75t_L g16624 ( 
.A(n_16108),
.B(n_11494),
.Y(n_16624)
);

NAND2xp5_ASAP7_75t_L g16625 ( 
.A(n_16122),
.B(n_9923),
.Y(n_16625)
);

INVx1_ASAP7_75t_L g16626 ( 
.A(n_16220),
.Y(n_16626)
);

OR2x2_ASAP7_75t_L g16627 ( 
.A(n_16147),
.B(n_8664),
.Y(n_16627)
);

NAND2x1p5_ASAP7_75t_L g16628 ( 
.A(n_16244),
.B(n_8526),
.Y(n_16628)
);

INVx1_ASAP7_75t_L g16629 ( 
.A(n_16151),
.Y(n_16629)
);

AOI22xp5_ASAP7_75t_L g16630 ( 
.A1(n_16270),
.A2(n_16275),
.B1(n_16182),
.B2(n_16199),
.Y(n_16630)
);

INVx1_ASAP7_75t_L g16631 ( 
.A(n_16067),
.Y(n_16631)
);

INVxp67_ASAP7_75t_SL g16632 ( 
.A(n_16148),
.Y(n_16632)
);

AND2x4_ASAP7_75t_SL g16633 ( 
.A(n_16119),
.B(n_7042),
.Y(n_16633)
);

INVx1_ASAP7_75t_L g16634 ( 
.A(n_16064),
.Y(n_16634)
);

AOI22xp33_ASAP7_75t_SL g16635 ( 
.A1(n_16208),
.A2(n_8559),
.B1(n_8568),
.B2(n_8530),
.Y(n_16635)
);

INVx1_ASAP7_75t_L g16636 ( 
.A(n_16062),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_16196),
.Y(n_16637)
);

INVx1_ASAP7_75t_L g16638 ( 
.A(n_16384),
.Y(n_16638)
);

INVx1_ASAP7_75t_L g16639 ( 
.A(n_16136),
.Y(n_16639)
);

OAI31xp33_ASAP7_75t_L g16640 ( 
.A1(n_16561),
.A2(n_8491),
.A3(n_8703),
.B(n_8439),
.Y(n_16640)
);

XOR2xp5_ASAP7_75t_L g16641 ( 
.A(n_16068),
.B(n_7933),
.Y(n_16641)
);

OAI22xp33_ASAP7_75t_L g16642 ( 
.A1(n_16383),
.A2(n_8559),
.B1(n_8568),
.B2(n_8530),
.Y(n_16642)
);

INVx1_ASAP7_75t_SL g16643 ( 
.A(n_16381),
.Y(n_16643)
);

NAND2xp5_ASAP7_75t_L g16644 ( 
.A(n_16181),
.B(n_9923),
.Y(n_16644)
);

AOI22xp33_ASAP7_75t_L g16645 ( 
.A1(n_16306),
.A2(n_8559),
.B1(n_8568),
.B2(n_8530),
.Y(n_16645)
);

INVx1_ASAP7_75t_L g16646 ( 
.A(n_16236),
.Y(n_16646)
);

OR2x6_ASAP7_75t_L g16647 ( 
.A(n_16218),
.B(n_7139),
.Y(n_16647)
);

NAND2xp5_ASAP7_75t_L g16648 ( 
.A(n_16172),
.B(n_16173),
.Y(n_16648)
);

INVx1_ASAP7_75t_L g16649 ( 
.A(n_16411),
.Y(n_16649)
);

NAND4xp25_ASAP7_75t_L g16650 ( 
.A(n_16101),
.B(n_7961),
.C(n_8722),
.D(n_8717),
.Y(n_16650)
);

AND2x2_ASAP7_75t_L g16651 ( 
.A(n_16093),
.B(n_11507),
.Y(n_16651)
);

INVx1_ASAP7_75t_L g16652 ( 
.A(n_16442),
.Y(n_16652)
);

INVx1_ASAP7_75t_L g16653 ( 
.A(n_16249),
.Y(n_16653)
);

AND2x2_ASAP7_75t_L g16654 ( 
.A(n_16081),
.B(n_11507),
.Y(n_16654)
);

INVx1_ASAP7_75t_L g16655 ( 
.A(n_16451),
.Y(n_16655)
);

INVx1_ASAP7_75t_L g16656 ( 
.A(n_16088),
.Y(n_16656)
);

NAND2xp5_ASAP7_75t_L g16657 ( 
.A(n_16334),
.B(n_9924),
.Y(n_16657)
);

HB1xp67_ASAP7_75t_L g16658 ( 
.A(n_16457),
.Y(n_16658)
);

O2A1O1Ixp33_ASAP7_75t_L g16659 ( 
.A1(n_16080),
.A2(n_9146),
.B(n_9152),
.C(n_9148),
.Y(n_16659)
);

OAI22xp5_ASAP7_75t_L g16660 ( 
.A1(n_16126),
.A2(n_16362),
.B1(n_16466),
.B2(n_16160),
.Y(n_16660)
);

NAND2xp5_ASAP7_75t_L g16661 ( 
.A(n_16086),
.B(n_16224),
.Y(n_16661)
);

INVx1_ASAP7_75t_L g16662 ( 
.A(n_16098),
.Y(n_16662)
);

INVx3_ASAP7_75t_L g16663 ( 
.A(n_16339),
.Y(n_16663)
);

INVx1_ASAP7_75t_L g16664 ( 
.A(n_16090),
.Y(n_16664)
);

INVxp67_ASAP7_75t_L g16665 ( 
.A(n_16529),
.Y(n_16665)
);

AND2x2_ASAP7_75t_L g16666 ( 
.A(n_16095),
.B(n_16250),
.Y(n_16666)
);

NAND2xp5_ASAP7_75t_L g16667 ( 
.A(n_16294),
.B(n_9924),
.Y(n_16667)
);

INVx1_ASAP7_75t_SL g16668 ( 
.A(n_16123),
.Y(n_16668)
);

INVx1_ASAP7_75t_L g16669 ( 
.A(n_16241),
.Y(n_16669)
);

INVx1_ASAP7_75t_L g16670 ( 
.A(n_16338),
.Y(n_16670)
);

INVx1_ASAP7_75t_L g16671 ( 
.A(n_16380),
.Y(n_16671)
);

NAND2xp5_ASAP7_75t_L g16672 ( 
.A(n_16110),
.B(n_9929),
.Y(n_16672)
);

INVx1_ASAP7_75t_L g16673 ( 
.A(n_16085),
.Y(n_16673)
);

AND2x4_ASAP7_75t_L g16674 ( 
.A(n_16457),
.B(n_11526),
.Y(n_16674)
);

NAND2xp5_ASAP7_75t_L g16675 ( 
.A(n_16114),
.B(n_9929),
.Y(n_16675)
);

INVx1_ASAP7_75t_L g16676 ( 
.A(n_16082),
.Y(n_16676)
);

AND2x4_ASAP7_75t_L g16677 ( 
.A(n_16360),
.B(n_11526),
.Y(n_16677)
);

OAI22xp33_ASAP7_75t_L g16678 ( 
.A1(n_16219),
.A2(n_8559),
.B1(n_8568),
.B2(n_8530),
.Y(n_16678)
);

AND2x2_ASAP7_75t_L g16679 ( 
.A(n_16301),
.B(n_11536),
.Y(n_16679)
);

NAND2xp5_ASAP7_75t_L g16680 ( 
.A(n_16157),
.B(n_9955),
.Y(n_16680)
);

INVx1_ASAP7_75t_L g16681 ( 
.A(n_16100),
.Y(n_16681)
);

INVx2_ASAP7_75t_L g16682 ( 
.A(n_16534),
.Y(n_16682)
);

NOR2xp33_ASAP7_75t_SL g16683 ( 
.A(n_16102),
.B(n_8530),
.Y(n_16683)
);

NOR3xp33_ASAP7_75t_L g16684 ( 
.A(n_16286),
.B(n_10975),
.C(n_10925),
.Y(n_16684)
);

OR2x2_ASAP7_75t_L g16685 ( 
.A(n_16109),
.B(n_8678),
.Y(n_16685)
);

INVx2_ASAP7_75t_L g16686 ( 
.A(n_16494),
.Y(n_16686)
);

INVxp33_ASAP7_75t_L g16687 ( 
.A(n_16541),
.Y(n_16687)
);

OAI22xp33_ASAP7_75t_L g16688 ( 
.A1(n_16558),
.A2(n_8568),
.B1(n_8595),
.B2(n_8559),
.Y(n_16688)
);

INVxp33_ASAP7_75t_L g16689 ( 
.A(n_16113),
.Y(n_16689)
);

INVx1_ASAP7_75t_L g16690 ( 
.A(n_16159),
.Y(n_16690)
);

OA222x2_ASAP7_75t_L g16691 ( 
.A1(n_16416),
.A2(n_8022),
.B1(n_7768),
.B2(n_8186),
.C1(n_8038),
.C2(n_7917),
.Y(n_16691)
);

AND2x2_ASAP7_75t_L g16692 ( 
.A(n_16305),
.B(n_16254),
.Y(n_16692)
);

AOI22xp5_ASAP7_75t_L g16693 ( 
.A1(n_16333),
.A2(n_8559),
.B1(n_8595),
.B2(n_8568),
.Y(n_16693)
);

NAND2xp33_ASAP7_75t_L g16694 ( 
.A(n_16205),
.B(n_8559),
.Y(n_16694)
);

INVx1_ASAP7_75t_L g16695 ( 
.A(n_16075),
.Y(n_16695)
);

INVx1_ASAP7_75t_L g16696 ( 
.A(n_16175),
.Y(n_16696)
);

NAND2x1p5_ASAP7_75t_L g16697 ( 
.A(n_16437),
.B(n_8559),
.Y(n_16697)
);

AOI21xp5_ASAP7_75t_L g16698 ( 
.A1(n_16516),
.A2(n_10119),
.B(n_10118),
.Y(n_16698)
);

INVx1_ASAP7_75t_SL g16699 ( 
.A(n_16361),
.Y(n_16699)
);

AOI22xp5_ASAP7_75t_L g16700 ( 
.A1(n_16453),
.A2(n_8568),
.B1(n_8606),
.B2(n_8595),
.Y(n_16700)
);

INVx2_ASAP7_75t_L g16701 ( 
.A(n_16392),
.Y(n_16701)
);

A2O1A1Ixp33_ASAP7_75t_L g16702 ( 
.A1(n_16112),
.A2(n_11025),
.B(n_11031),
.C(n_11021),
.Y(n_16702)
);

INVx1_ASAP7_75t_L g16703 ( 
.A(n_16212),
.Y(n_16703)
);

NAND4xp75_ASAP7_75t_SL g16704 ( 
.A(n_16326),
.B(n_10082),
.C(n_10163),
.D(n_10039),
.Y(n_16704)
);

NAND2xp5_ASAP7_75t_L g16705 ( 
.A(n_16336),
.B(n_9955),
.Y(n_16705)
);

OR2x2_ASAP7_75t_L g16706 ( 
.A(n_16177),
.B(n_8678),
.Y(n_16706)
);

INVx1_ASAP7_75t_L g16707 ( 
.A(n_16509),
.Y(n_16707)
);

NAND3xp33_ASAP7_75t_L g16708 ( 
.A(n_16111),
.B(n_9228),
.C(n_9126),
.Y(n_16708)
);

INVx1_ASAP7_75t_L g16709 ( 
.A(n_16174),
.Y(n_16709)
);

INVx2_ASAP7_75t_SL g16710 ( 
.A(n_16162),
.Y(n_16710)
);

INVx2_ASAP7_75t_L g16711 ( 
.A(n_16490),
.Y(n_16711)
);

INVx2_ASAP7_75t_L g16712 ( 
.A(n_16428),
.Y(n_16712)
);

INVx1_ASAP7_75t_L g16713 ( 
.A(n_16337),
.Y(n_16713)
);

INVx1_ASAP7_75t_L g16714 ( 
.A(n_16079),
.Y(n_16714)
);

NOR2x1_ASAP7_75t_L g16715 ( 
.A(n_16091),
.B(n_10118),
.Y(n_16715)
);

OR2x6_ASAP7_75t_L g16716 ( 
.A(n_16416),
.B(n_7139),
.Y(n_16716)
);

HB1xp67_ASAP7_75t_L g16717 ( 
.A(n_16198),
.Y(n_16717)
);

INVx1_ASAP7_75t_L g16718 ( 
.A(n_16350),
.Y(n_16718)
);

NAND2xp33_ASAP7_75t_L g16719 ( 
.A(n_16310),
.B(n_8568),
.Y(n_16719)
);

INVx1_ASAP7_75t_L g16720 ( 
.A(n_16370),
.Y(n_16720)
);

OAI22xp5_ASAP7_75t_L g16721 ( 
.A1(n_16274),
.A2(n_8606),
.B1(n_8674),
.B2(n_8595),
.Y(n_16721)
);

OR2x2_ASAP7_75t_L g16722 ( 
.A(n_16373),
.B(n_10118),
.Y(n_16722)
);

INVx1_ASAP7_75t_L g16723 ( 
.A(n_16382),
.Y(n_16723)
);

O2A1O1Ixp33_ASAP7_75t_SL g16724 ( 
.A1(n_16092),
.A2(n_7978),
.B(n_8021),
.C(n_7908),
.Y(n_16724)
);

INVx2_ASAP7_75t_L g16725 ( 
.A(n_16439),
.Y(n_16725)
);

NAND2xp5_ASAP7_75t_L g16726 ( 
.A(n_16394),
.B(n_16323),
.Y(n_16726)
);

INVx1_ASAP7_75t_L g16727 ( 
.A(n_16325),
.Y(n_16727)
);

AND2x2_ASAP7_75t_L g16728 ( 
.A(n_16324),
.B(n_11536),
.Y(n_16728)
);

INVxp67_ASAP7_75t_L g16729 ( 
.A(n_16216),
.Y(n_16729)
);

NAND2xp5_ASAP7_75t_L g16730 ( 
.A(n_16331),
.B(n_9958),
.Y(n_16730)
);

INVx1_ASAP7_75t_L g16731 ( 
.A(n_16452),
.Y(n_16731)
);

AOI22xp5_ASAP7_75t_L g16732 ( 
.A1(n_16298),
.A2(n_16194),
.B1(n_16459),
.B2(n_16460),
.Y(n_16732)
);

INVx1_ASAP7_75t_L g16733 ( 
.A(n_16327),
.Y(n_16733)
);

INVx1_ASAP7_75t_L g16734 ( 
.A(n_16107),
.Y(n_16734)
);

INVx1_ASAP7_75t_L g16735 ( 
.A(n_16454),
.Y(n_16735)
);

INVx1_ASAP7_75t_L g16736 ( 
.A(n_16401),
.Y(n_16736)
);

NOR4xp25_ASAP7_75t_L g16737 ( 
.A(n_16127),
.B(n_9148),
.C(n_9152),
.D(n_9146),
.Y(n_16737)
);

INVx1_ASAP7_75t_L g16738 ( 
.A(n_16407),
.Y(n_16738)
);

INVx1_ASAP7_75t_L g16739 ( 
.A(n_16283),
.Y(n_16739)
);

NAND4xp75_ASAP7_75t_L g16740 ( 
.A(n_16154),
.B(n_10055),
.C(n_9228),
.D(n_9126),
.Y(n_16740)
);

AND3x1_ASAP7_75t_SL g16741 ( 
.A(n_16297),
.B(n_16302),
.C(n_16166),
.Y(n_16741)
);

OAI322xp33_ASAP7_75t_L g16742 ( 
.A1(n_16155),
.A2(n_9146),
.A3(n_9175),
.B1(n_9148),
.B2(n_9180),
.C1(n_9179),
.C2(n_9152),
.Y(n_16742)
);

INVx1_ASAP7_75t_L g16743 ( 
.A(n_16441),
.Y(n_16743)
);

HB1xp67_ASAP7_75t_L g16744 ( 
.A(n_16207),
.Y(n_16744)
);

INVx1_ASAP7_75t_L g16745 ( 
.A(n_16446),
.Y(n_16745)
);

HB1xp67_ASAP7_75t_L g16746 ( 
.A(n_16207),
.Y(n_16746)
);

AND2x2_ASAP7_75t_L g16747 ( 
.A(n_16279),
.B(n_10119),
.Y(n_16747)
);

AOI22xp33_ASAP7_75t_L g16748 ( 
.A1(n_16317),
.A2(n_8606),
.B1(n_8674),
.B2(n_8595),
.Y(n_16748)
);

OR2x6_ASAP7_75t_L g16749 ( 
.A(n_16234),
.B(n_7139),
.Y(n_16749)
);

OAI32xp33_ASAP7_75t_L g16750 ( 
.A1(n_16163),
.A2(n_9180),
.A3(n_9179),
.B1(n_9175),
.B2(n_7768),
.Y(n_16750)
);

INVx2_ASAP7_75t_L g16751 ( 
.A(n_16483),
.Y(n_16751)
);

INVx1_ASAP7_75t_L g16752 ( 
.A(n_16491),
.Y(n_16752)
);

INVx1_ASAP7_75t_L g16753 ( 
.A(n_16526),
.Y(n_16753)
);

AND2x2_ASAP7_75t_L g16754 ( 
.A(n_16308),
.B(n_10119),
.Y(n_16754)
);

OA222x2_ASAP7_75t_L g16755 ( 
.A1(n_16144),
.A2(n_8022),
.B1(n_7768),
.B2(n_8186),
.C1(n_8038),
.C2(n_7917),
.Y(n_16755)
);

AND2x2_ASAP7_75t_L g16756 ( 
.A(n_16193),
.B(n_10120),
.Y(n_16756)
);

INVx1_ASAP7_75t_L g16757 ( 
.A(n_16421),
.Y(n_16757)
);

INVx1_ASAP7_75t_SL g16758 ( 
.A(n_16187),
.Y(n_16758)
);

AND2x2_ASAP7_75t_L g16759 ( 
.A(n_16245),
.B(n_10120),
.Y(n_16759)
);

NAND2x1_ASAP7_75t_L g16760 ( 
.A(n_16335),
.B(n_10120),
.Y(n_16760)
);

INVx1_ASAP7_75t_SL g16761 ( 
.A(n_16132),
.Y(n_16761)
);

NOR2xp33_ASAP7_75t_SL g16762 ( 
.A(n_16455),
.B(n_8595),
.Y(n_16762)
);

INVx2_ASAP7_75t_L g16763 ( 
.A(n_16328),
.Y(n_16763)
);

INVx1_ASAP7_75t_L g16764 ( 
.A(n_16318),
.Y(n_16764)
);

INVxp67_ASAP7_75t_L g16765 ( 
.A(n_16164),
.Y(n_16765)
);

NAND2xp5_ASAP7_75t_L g16766 ( 
.A(n_16406),
.B(n_9958),
.Y(n_16766)
);

INVxp67_ASAP7_75t_L g16767 ( 
.A(n_16227),
.Y(n_16767)
);

AND4x1_ASAP7_75t_L g16768 ( 
.A(n_16255),
.B(n_7572),
.C(n_7471),
.D(n_8552),
.Y(n_16768)
);

NAND2xp5_ASAP7_75t_L g16769 ( 
.A(n_16176),
.B(n_9961),
.Y(n_16769)
);

O2A1O1Ixp5_ASAP7_75t_R g16770 ( 
.A1(n_16272),
.A2(n_8556),
.B(n_7067),
.C(n_7062),
.Y(n_16770)
);

INVx1_ASAP7_75t_L g16771 ( 
.A(n_16135),
.Y(n_16771)
);

AOI211xp5_ASAP7_75t_L g16772 ( 
.A1(n_16133),
.A2(n_11070),
.B(n_11031),
.C(n_11244),
.Y(n_16772)
);

OR2x2_ASAP7_75t_L g16773 ( 
.A(n_16371),
.B(n_10123),
.Y(n_16773)
);

OAI211xp5_ASAP7_75t_L g16774 ( 
.A1(n_16104),
.A2(n_11070),
.B(n_9126),
.C(n_9228),
.Y(n_16774)
);

INVx6_ASAP7_75t_L g16775 ( 
.A(n_16372),
.Y(n_16775)
);

INVx1_ASAP7_75t_L g16776 ( 
.A(n_16448),
.Y(n_16776)
);

INVx2_ASAP7_75t_L g16777 ( 
.A(n_16167),
.Y(n_16777)
);

INVx1_ASAP7_75t_L g16778 ( 
.A(n_16414),
.Y(n_16778)
);

INVx1_ASAP7_75t_L g16779 ( 
.A(n_16417),
.Y(n_16779)
);

AND2x2_ASAP7_75t_L g16780 ( 
.A(n_16344),
.B(n_10123),
.Y(n_16780)
);

OAI22xp5_ASAP7_75t_L g16781 ( 
.A1(n_16368),
.A2(n_8606),
.B1(n_8674),
.B2(n_8595),
.Y(n_16781)
);

A2O1A1Ixp33_ASAP7_75t_L g16782 ( 
.A1(n_16264),
.A2(n_11245),
.B(n_11280),
.C(n_11244),
.Y(n_16782)
);

INVxp67_ASAP7_75t_L g16783 ( 
.A(n_16228),
.Y(n_16783)
);

OAI22xp5_ASAP7_75t_L g16784 ( 
.A1(n_16229),
.A2(n_8606),
.B1(n_8674),
.B2(n_8595),
.Y(n_16784)
);

AND2x2_ASAP7_75t_L g16785 ( 
.A(n_16353),
.B(n_10123),
.Y(n_16785)
);

INVx2_ASAP7_75t_L g16786 ( 
.A(n_16168),
.Y(n_16786)
);

NOR3xp33_ASAP7_75t_L g16787 ( 
.A(n_16184),
.B(n_11280),
.C(n_11245),
.Y(n_16787)
);

AOI21x1_ASAP7_75t_L g16788 ( 
.A1(n_16423),
.A2(n_9268),
.B(n_9236),
.Y(n_16788)
);

AND2x4_ASAP7_75t_L g16789 ( 
.A(n_16363),
.B(n_11302),
.Y(n_16789)
);

INVx2_ASAP7_75t_L g16790 ( 
.A(n_16304),
.Y(n_16790)
);

OR2x2_ASAP7_75t_L g16791 ( 
.A(n_16248),
.B(n_10127),
.Y(n_16791)
);

AND2x2_ASAP7_75t_L g16792 ( 
.A(n_16431),
.B(n_10127),
.Y(n_16792)
);

A2O1A1Ixp33_ASAP7_75t_L g16793 ( 
.A1(n_16545),
.A2(n_11324),
.B(n_11340),
.C(n_11302),
.Y(n_16793)
);

INVx2_ASAP7_75t_L g16794 ( 
.A(n_16190),
.Y(n_16794)
);

AO22x1_ASAP7_75t_L g16795 ( 
.A1(n_16492),
.A2(n_6757),
.B1(n_6781),
.B2(n_6648),
.Y(n_16795)
);

OR2x2_ASAP7_75t_L g16796 ( 
.A(n_16232),
.B(n_10127),
.Y(n_16796)
);

OAI22xp5_ASAP7_75t_L g16797 ( 
.A1(n_16191),
.A2(n_8674),
.B1(n_8851),
.B2(n_8606),
.Y(n_16797)
);

INVx1_ASAP7_75t_L g16798 ( 
.A(n_16197),
.Y(n_16798)
);

NAND2xp5_ASAP7_75t_L g16799 ( 
.A(n_16340),
.B(n_9961),
.Y(n_16799)
);

O2A1O1Ixp5_ASAP7_75t_R g16800 ( 
.A1(n_16410),
.A2(n_6741),
.B(n_6748),
.C(n_6830),
.Y(n_16800)
);

NAND2xp5_ASAP7_75t_SL g16801 ( 
.A(n_16332),
.B(n_8606),
.Y(n_16801)
);

INVx2_ASAP7_75t_L g16802 ( 
.A(n_16203),
.Y(n_16802)
);

NAND2xp5_ASAP7_75t_L g16803 ( 
.A(n_16213),
.B(n_9967),
.Y(n_16803)
);

INVx1_ASAP7_75t_L g16804 ( 
.A(n_16201),
.Y(n_16804)
);

NAND2xp5_ASAP7_75t_L g16805 ( 
.A(n_16389),
.B(n_9967),
.Y(n_16805)
);

OAI21xp33_ASAP7_75t_L g16806 ( 
.A1(n_16284),
.A2(n_9180),
.B(n_11324),
.Y(n_16806)
);

AOI33xp33_ASAP7_75t_L g16807 ( 
.A1(n_16267),
.A2(n_8085),
.A3(n_7978),
.B1(n_8103),
.B2(n_8021),
.B3(n_7908),
.Y(n_16807)
);

NAND2xp5_ASAP7_75t_L g16808 ( 
.A(n_16390),
.B(n_9970),
.Y(n_16808)
);

A2O1A1Ixp33_ASAP7_75t_L g16809 ( 
.A1(n_16211),
.A2(n_11340),
.B(n_9287),
.C(n_9330),
.Y(n_16809)
);

INVxp33_ASAP7_75t_L g16810 ( 
.A(n_16312),
.Y(n_16810)
);

INVx2_ASAP7_75t_SL g16811 ( 
.A(n_16420),
.Y(n_16811)
);

AOI22xp5_ASAP7_75t_L g16812 ( 
.A1(n_16364),
.A2(n_8606),
.B1(n_8851),
.B2(n_8674),
.Y(n_16812)
);

INVx1_ASAP7_75t_L g16813 ( 
.A(n_16210),
.Y(n_16813)
);

AOI22xp5_ASAP7_75t_L g16814 ( 
.A1(n_16393),
.A2(n_8674),
.B1(n_8867),
.B2(n_8851),
.Y(n_16814)
);

AOI22xp5_ASAP7_75t_L g16815 ( 
.A1(n_16444),
.A2(n_16479),
.B1(n_16243),
.B2(n_16313),
.Y(n_16815)
);

XNOR2xp5_ASAP7_75t_L g16816 ( 
.A(n_16508),
.B(n_8852),
.Y(n_16816)
);

HB1xp67_ASAP7_75t_L g16817 ( 
.A(n_16431),
.Y(n_16817)
);

AND2x2_ASAP7_75t_L g16818 ( 
.A(n_16348),
.B(n_16531),
.Y(n_16818)
);

INVx1_ASAP7_75t_L g16819 ( 
.A(n_16186),
.Y(n_16819)
);

INVx3_ASAP7_75t_L g16820 ( 
.A(n_16539),
.Y(n_16820)
);

A2O1A1Ixp33_ASAP7_75t_L g16821 ( 
.A1(n_16485),
.A2(n_9287),
.B(n_9330),
.C(n_9270),
.Y(n_16821)
);

INVx1_ASAP7_75t_L g16822 ( 
.A(n_16189),
.Y(n_16822)
);

OR2x2_ASAP7_75t_L g16823 ( 
.A(n_16543),
.B(n_16546),
.Y(n_16823)
);

INVx1_ASAP7_75t_L g16824 ( 
.A(n_16153),
.Y(n_16824)
);

NAND2xp5_ASAP7_75t_L g16825 ( 
.A(n_16555),
.B(n_9970),
.Y(n_16825)
);

AOI22xp33_ASAP7_75t_L g16826 ( 
.A1(n_16237),
.A2(n_8851),
.B1(n_8867),
.B2(n_8674),
.Y(n_16826)
);

INVx1_ASAP7_75t_L g16827 ( 
.A(n_16260),
.Y(n_16827)
);

INVxp67_ASAP7_75t_SL g16828 ( 
.A(n_16214),
.Y(n_16828)
);

OAI22xp5_ASAP7_75t_L g16829 ( 
.A1(n_16263),
.A2(n_8867),
.B1(n_8939),
.B2(n_8851),
.Y(n_16829)
);

OAI22xp5_ASAP7_75t_L g16830 ( 
.A1(n_16251),
.A2(n_8867),
.B1(n_8939),
.B2(n_8851),
.Y(n_16830)
);

NOR2xp67_ASAP7_75t_R g16831 ( 
.A(n_16557),
.B(n_8851),
.Y(n_16831)
);

NOR4xp25_ASAP7_75t_L g16832 ( 
.A(n_16226),
.B(n_9974),
.C(n_9981),
.D(n_9972),
.Y(n_16832)
);

INVx1_ASAP7_75t_L g16833 ( 
.A(n_16430),
.Y(n_16833)
);

NAND2x2_ASAP7_75t_L g16834 ( 
.A(n_16525),
.B(n_6657),
.Y(n_16834)
);

OR3x2_ASAP7_75t_L g16835 ( 
.A(n_16521),
.B(n_9268),
.C(n_9236),
.Y(n_16835)
);

OAI322xp33_ASAP7_75t_L g16836 ( 
.A1(n_16355),
.A2(n_8832),
.A3(n_8995),
.B1(n_8778),
.B2(n_7929),
.C1(n_7772),
.C2(n_7872),
.Y(n_16836)
);

INVx2_ASAP7_75t_L g16837 ( 
.A(n_16427),
.Y(n_16837)
);

NAND2xp5_ASAP7_75t_L g16838 ( 
.A(n_16440),
.B(n_16315),
.Y(n_16838)
);

INVx1_ASAP7_75t_L g16839 ( 
.A(n_16341),
.Y(n_16839)
);

NAND2xp5_ASAP7_75t_L g16840 ( 
.A(n_16461),
.B(n_16511),
.Y(n_16840)
);

AND2x2_ASAP7_75t_L g16841 ( 
.A(n_16435),
.B(n_10130),
.Y(n_16841)
);

INVx1_ASAP7_75t_SL g16842 ( 
.A(n_16152),
.Y(n_16842)
);

INVx1_ASAP7_75t_L g16843 ( 
.A(n_16322),
.Y(n_16843)
);

INVx1_ASAP7_75t_L g16844 ( 
.A(n_16240),
.Y(n_16844)
);

INVx1_ASAP7_75t_L g16845 ( 
.A(n_16367),
.Y(n_16845)
);

INVxp33_ASAP7_75t_L g16846 ( 
.A(n_16280),
.Y(n_16846)
);

AND2x4_ASAP7_75t_SL g16847 ( 
.A(n_16539),
.B(n_7042),
.Y(n_16847)
);

INVx1_ASAP7_75t_L g16848 ( 
.A(n_16321),
.Y(n_16848)
);

OR2x2_ASAP7_75t_L g16849 ( 
.A(n_16239),
.B(n_10130),
.Y(n_16849)
);

NAND2xp5_ASAP7_75t_L g16850 ( 
.A(n_16209),
.B(n_16475),
.Y(n_16850)
);

INVx1_ASAP7_75t_L g16851 ( 
.A(n_16319),
.Y(n_16851)
);

AOI22xp5_ASAP7_75t_L g16852 ( 
.A1(n_16503),
.A2(n_8867),
.B1(n_8939),
.B2(n_8851),
.Y(n_16852)
);

INVx1_ASAP7_75t_L g16853 ( 
.A(n_16230),
.Y(n_16853)
);

INVx1_ASAP7_75t_L g16854 ( 
.A(n_16222),
.Y(n_16854)
);

AOI22xp5_ASAP7_75t_L g16855 ( 
.A1(n_16515),
.A2(n_8939),
.B1(n_8948),
.B2(n_8867),
.Y(n_16855)
);

NAND2xp5_ASAP7_75t_L g16856 ( 
.A(n_16347),
.B(n_9972),
.Y(n_16856)
);

INVx1_ASAP7_75t_L g16857 ( 
.A(n_16303),
.Y(n_16857)
);

A2O1A1Ixp33_ASAP7_75t_L g16858 ( 
.A1(n_16287),
.A2(n_9465),
.B(n_9504),
.C(n_9270),
.Y(n_16858)
);

INVx1_ASAP7_75t_L g16859 ( 
.A(n_16307),
.Y(n_16859)
);

AOI22xp5_ASAP7_75t_L g16860 ( 
.A1(n_16343),
.A2(n_8939),
.B1(n_8948),
.B2(n_8867),
.Y(n_16860)
);

O2A1O1Ixp5_ASAP7_75t_R g16861 ( 
.A1(n_16262),
.A2(n_6741),
.B(n_6748),
.C(n_6830),
.Y(n_16861)
);

INVx1_ASAP7_75t_L g16862 ( 
.A(n_16195),
.Y(n_16862)
);

AOI32xp33_ASAP7_75t_L g16863 ( 
.A1(n_16356),
.A2(n_9653),
.A3(n_9905),
.B1(n_9651),
.B2(n_9419),
.Y(n_16863)
);

INVx1_ASAP7_75t_L g16864 ( 
.A(n_16206),
.Y(n_16864)
);

NAND4xp75_ASAP7_75t_L g16865 ( 
.A(n_16467),
.B(n_10055),
.C(n_9228),
.D(n_9126),
.Y(n_16865)
);

NAND4xp25_ASAP7_75t_L g16866 ( 
.A(n_16542),
.B(n_7961),
.C(n_8722),
.D(n_8717),
.Y(n_16866)
);

INVx4_ASAP7_75t_L g16867 ( 
.A(n_16342),
.Y(n_16867)
);

INVxp67_ASAP7_75t_SL g16868 ( 
.A(n_16204),
.Y(n_16868)
);

OR2x2_ASAP7_75t_L g16869 ( 
.A(n_16391),
.B(n_10130),
.Y(n_16869)
);

OR2x2_ASAP7_75t_L g16870 ( 
.A(n_16456),
.B(n_10132),
.Y(n_16870)
);

AND2x2_ASAP7_75t_L g16871 ( 
.A(n_16544),
.B(n_16540),
.Y(n_16871)
);

INVx1_ASAP7_75t_L g16872 ( 
.A(n_16273),
.Y(n_16872)
);

AOI22xp5_ASAP7_75t_L g16873 ( 
.A1(n_16235),
.A2(n_8939),
.B1(n_8948),
.B2(n_8867),
.Y(n_16873)
);

INVxp67_ASAP7_75t_L g16874 ( 
.A(n_16346),
.Y(n_16874)
);

INVx2_ASAP7_75t_L g16875 ( 
.A(n_16378),
.Y(n_16875)
);

INVx1_ASAP7_75t_L g16876 ( 
.A(n_16169),
.Y(n_16876)
);

INVx2_ASAP7_75t_L g16877 ( 
.A(n_16320),
.Y(n_16877)
);

AOI32xp33_ASAP7_75t_L g16878 ( 
.A1(n_16413),
.A2(n_9653),
.A3(n_9905),
.B1(n_9651),
.B2(n_9419),
.Y(n_16878)
);

OR2x2_ASAP7_75t_L g16879 ( 
.A(n_16493),
.B(n_10132),
.Y(n_16879)
);

INVx1_ASAP7_75t_SL g16880 ( 
.A(n_16290),
.Y(n_16880)
);

OR2x2_ASAP7_75t_L g16881 ( 
.A(n_16480),
.B(n_10132),
.Y(n_16881)
);

INVx1_ASAP7_75t_L g16882 ( 
.A(n_16299),
.Y(n_16882)
);

A2O1A1Ixp33_ASAP7_75t_L g16883 ( 
.A1(n_16202),
.A2(n_9504),
.B(n_9641),
.C(n_9465),
.Y(n_16883)
);

OAI21xp5_ASAP7_75t_L g16884 ( 
.A1(n_16547),
.A2(n_9663),
.B(n_9641),
.Y(n_16884)
);

INVx1_ASAP7_75t_L g16885 ( 
.A(n_16296),
.Y(n_16885)
);

AND2x4_ASAP7_75t_L g16886 ( 
.A(n_16468),
.B(n_10142),
.Y(n_16886)
);

AND2x4_ASAP7_75t_L g16887 ( 
.A(n_16471),
.B(n_10142),
.Y(n_16887)
);

AOI33xp33_ASAP7_75t_L g16888 ( 
.A1(n_16550),
.A2(n_8274),
.A3(n_8103),
.B1(n_8311),
.B2(n_8228),
.B3(n_8085),
.Y(n_16888)
);

OR2x2_ASAP7_75t_L g16889 ( 
.A(n_16424),
.B(n_10142),
.Y(n_16889)
);

NAND2xp5_ASAP7_75t_L g16890 ( 
.A(n_16354),
.B(n_9974),
.Y(n_16890)
);

AOI211xp5_ASAP7_75t_L g16891 ( 
.A1(n_16476),
.A2(n_6757),
.B(n_6781),
.C(n_6648),
.Y(n_16891)
);

INVx1_ASAP7_75t_SL g16892 ( 
.A(n_16295),
.Y(n_16892)
);

INVx2_ASAP7_75t_L g16893 ( 
.A(n_16386),
.Y(n_16893)
);

NAND2xp5_ASAP7_75t_L g16894 ( 
.A(n_16478),
.B(n_9981),
.Y(n_16894)
);

INVx1_ASAP7_75t_SL g16895 ( 
.A(n_16253),
.Y(n_16895)
);

NAND2x1_ASAP7_75t_L g16896 ( 
.A(n_16335),
.B(n_10145),
.Y(n_16896)
);

OAI211xp5_ASAP7_75t_L g16897 ( 
.A1(n_16488),
.A2(n_9275),
.B(n_10055),
.C(n_10314),
.Y(n_16897)
);

INVxp67_ASAP7_75t_L g16898 ( 
.A(n_16387),
.Y(n_16898)
);

AOI22xp5_ASAP7_75t_L g16899 ( 
.A1(n_16505),
.A2(n_8948),
.B1(n_9008),
.B2(n_8939),
.Y(n_16899)
);

NAND4xp75_ASAP7_75t_L g16900 ( 
.A(n_16484),
.B(n_10055),
.C(n_8405),
.D(n_8359),
.Y(n_16900)
);

INVx2_ASAP7_75t_L g16901 ( 
.A(n_16396),
.Y(n_16901)
);

XOR2x2_ASAP7_75t_L g16902 ( 
.A(n_16496),
.B(n_16499),
.Y(n_16902)
);

OR2x2_ASAP7_75t_L g16903 ( 
.A(n_16433),
.B(n_10145),
.Y(n_16903)
);

INVx2_ASAP7_75t_SL g16904 ( 
.A(n_16271),
.Y(n_16904)
);

INVx1_ASAP7_75t_SL g16905 ( 
.A(n_16549),
.Y(n_16905)
);

INVx1_ASAP7_75t_L g16906 ( 
.A(n_16300),
.Y(n_16906)
);

OAI32xp33_ASAP7_75t_L g16907 ( 
.A1(n_16533),
.A2(n_7768),
.A3(n_8038),
.B1(n_8022),
.B2(n_7917),
.Y(n_16907)
);

OAI22xp5_ASAP7_75t_L g16908 ( 
.A1(n_16510),
.A2(n_8948),
.B1(n_9008),
.B2(n_8939),
.Y(n_16908)
);

INVxp67_ASAP7_75t_SL g16909 ( 
.A(n_16352),
.Y(n_16909)
);

INVx1_ASAP7_75t_L g16910 ( 
.A(n_16329),
.Y(n_16910)
);

NOR2xp33_ASAP7_75t_L g16911 ( 
.A(n_16518),
.B(n_10145),
.Y(n_16911)
);

OR2x2_ASAP7_75t_L g16912 ( 
.A(n_16552),
.B(n_10156),
.Y(n_16912)
);

INVx1_ASAP7_75t_L g16913 ( 
.A(n_16281),
.Y(n_16913)
);

INVx1_ASAP7_75t_L g16914 ( 
.A(n_16291),
.Y(n_16914)
);

NOR3xp33_ASAP7_75t_L g16915 ( 
.A(n_16519),
.B(n_9275),
.C(n_9663),
.Y(n_16915)
);

INVx2_ASAP7_75t_L g16916 ( 
.A(n_16398),
.Y(n_16916)
);

OAI221xp5_ASAP7_75t_SL g16917 ( 
.A1(n_16278),
.A2(n_8832),
.B1(n_8995),
.B2(n_8778),
.C(n_8440),
.Y(n_16917)
);

O2A1O1Ixp5_ASAP7_75t_R g16918 ( 
.A1(n_16288),
.A2(n_6830),
.B(n_6990),
.C(n_6970),
.Y(n_16918)
);

OAI322xp33_ASAP7_75t_L g16919 ( 
.A1(n_16185),
.A2(n_16535),
.A3(n_16528),
.B1(n_16536),
.B2(n_16538),
.C1(n_16532),
.C2(n_16520),
.Y(n_16919)
);

INVx1_ASAP7_75t_L g16920 ( 
.A(n_16366),
.Y(n_16920)
);

NOR2xp33_ASAP7_75t_L g16921 ( 
.A(n_16374),
.B(n_10156),
.Y(n_16921)
);

NAND2xp5_ASAP7_75t_L g16922 ( 
.A(n_16426),
.B(n_9998),
.Y(n_16922)
);

OAI22xp5_ASAP7_75t_L g16923 ( 
.A1(n_16500),
.A2(n_9008),
.B1(n_8948),
.B2(n_10156),
.Y(n_16923)
);

INVx1_ASAP7_75t_L g16924 ( 
.A(n_16375),
.Y(n_16924)
);

A2O1A1Ixp33_ASAP7_75t_L g16925 ( 
.A1(n_16276),
.A2(n_9724),
.B(n_9728),
.C(n_9691),
.Y(n_16925)
);

INVx1_ASAP7_75t_SL g16926 ( 
.A(n_16285),
.Y(n_16926)
);

INVx1_ASAP7_75t_SL g16927 ( 
.A(n_16282),
.Y(n_16927)
);

OAI22xp5_ASAP7_75t_L g16928 ( 
.A1(n_16150),
.A2(n_16463),
.B1(n_16271),
.B2(n_16345),
.Y(n_16928)
);

NAND2xp5_ASAP7_75t_L g16929 ( 
.A(n_16450),
.B(n_9998),
.Y(n_16929)
);

HB1xp67_ASAP7_75t_L g16930 ( 
.A(n_16335),
.Y(n_16930)
);

AND2x2_ASAP7_75t_L g16931 ( 
.A(n_16436),
.B(n_10171),
.Y(n_16931)
);

NAND2xp5_ASAP7_75t_L g16932 ( 
.A(n_16438),
.B(n_10004),
.Y(n_16932)
);

INVx1_ASAP7_75t_L g16933 ( 
.A(n_16377),
.Y(n_16933)
);

A2O1A1Ixp33_ASAP7_75t_L g16934 ( 
.A1(n_16292),
.A2(n_16252),
.B(n_16559),
.C(n_16180),
.Y(n_16934)
);

AOI22xp5_ASAP7_75t_L g16935 ( 
.A1(n_16422),
.A2(n_9008),
.B1(n_8948),
.B2(n_8722),
.Y(n_16935)
);

INVx1_ASAP7_75t_L g16936 ( 
.A(n_16379),
.Y(n_16936)
);

INVx1_ASAP7_75t_L g16937 ( 
.A(n_16316),
.Y(n_16937)
);

INVx2_ASAP7_75t_L g16938 ( 
.A(n_16399),
.Y(n_16938)
);

AND2x4_ASAP7_75t_L g16939 ( 
.A(n_16221),
.B(n_8717),
.Y(n_16939)
);

INVx1_ASAP7_75t_L g16940 ( 
.A(n_16223),
.Y(n_16940)
);

INVx2_ASAP7_75t_SL g16941 ( 
.A(n_16247),
.Y(n_16941)
);

OR2x2_ASAP7_75t_L g16942 ( 
.A(n_16289),
.B(n_10171),
.Y(n_16942)
);

AND2x2_ASAP7_75t_L g16943 ( 
.A(n_16269),
.B(n_10171),
.Y(n_16943)
);

NOR4xp25_ASAP7_75t_SL g16944 ( 
.A(n_16395),
.B(n_10010),
.C(n_10012),
.D(n_10004),
.Y(n_16944)
);

INVxp67_ASAP7_75t_SL g16945 ( 
.A(n_16231),
.Y(n_16945)
);

OR2x2_ASAP7_75t_L g16946 ( 
.A(n_16311),
.B(n_10173),
.Y(n_16946)
);

INVx2_ASAP7_75t_L g16947 ( 
.A(n_16403),
.Y(n_16947)
);

NAND3xp33_ASAP7_75t_L g16948 ( 
.A(n_16465),
.B(n_8161),
.C(n_8156),
.Y(n_16948)
);

INVx2_ASAP7_75t_L g16949 ( 
.A(n_16357),
.Y(n_16949)
);

HB1xp67_ASAP7_75t_L g16950 ( 
.A(n_16449),
.Y(n_16950)
);

BUFx2_ASAP7_75t_L g16951 ( 
.A(n_16425),
.Y(n_16951)
);

NAND2xp5_ASAP7_75t_L g16952 ( 
.A(n_16458),
.B(n_10010),
.Y(n_16952)
);

INVx2_ASAP7_75t_L g16953 ( 
.A(n_16524),
.Y(n_16953)
);

OR2x2_ASAP7_75t_L g16954 ( 
.A(n_16388),
.B(n_10173),
.Y(n_16954)
);

INVx1_ASAP7_75t_L g16955 ( 
.A(n_16238),
.Y(n_16955)
);

INVx1_ASAP7_75t_L g16956 ( 
.A(n_16246),
.Y(n_16956)
);

INVx1_ASAP7_75t_L g16957 ( 
.A(n_16256),
.Y(n_16957)
);

NAND2xp5_ASAP7_75t_L g16958 ( 
.A(n_16464),
.B(n_16470),
.Y(n_16958)
);

OR2x6_ASAP7_75t_L g16959 ( 
.A(n_16257),
.B(n_7139),
.Y(n_16959)
);

INVx1_ASAP7_75t_L g16960 ( 
.A(n_16258),
.Y(n_16960)
);

O2A1O1Ixp33_ASAP7_75t_L g16961 ( 
.A1(n_16261),
.A2(n_8161),
.B(n_8156),
.C(n_8098),
.Y(n_16961)
);

NOR2x1p5_ASAP7_75t_L g16962 ( 
.A(n_16293),
.B(n_8948),
.Y(n_16962)
);

INVx1_ASAP7_75t_L g16963 ( 
.A(n_16351),
.Y(n_16963)
);

OR2x6_ASAP7_75t_L g16964 ( 
.A(n_16477),
.B(n_7376),
.Y(n_16964)
);

OR2x2_ASAP7_75t_L g16965 ( 
.A(n_16400),
.B(n_10173),
.Y(n_16965)
);

AND2x2_ASAP7_75t_L g16966 ( 
.A(n_16188),
.B(n_10186),
.Y(n_16966)
);

OR2x2_ASAP7_75t_L g16967 ( 
.A(n_16504),
.B(n_10186),
.Y(n_16967)
);

AOI22xp33_ASAP7_75t_L g16968 ( 
.A1(n_16556),
.A2(n_9008),
.B1(n_8536),
.B2(n_8501),
.Y(n_16968)
);

NOR2xp33_ASAP7_75t_L g16969 ( 
.A(n_16563),
.B(n_16495),
.Y(n_16969)
);

NOR2xp67_ASAP7_75t_SL g16970 ( 
.A(n_16622),
.B(n_16663),
.Y(n_16970)
);

NAND2xp5_ASAP7_75t_L g16971 ( 
.A(n_16604),
.B(n_16537),
.Y(n_16971)
);

NAND3xp33_ASAP7_75t_L g16972 ( 
.A(n_16612),
.B(n_16178),
.C(n_16434),
.Y(n_16972)
);

HB1xp67_ASAP7_75t_L g16973 ( 
.A(n_16658),
.Y(n_16973)
);

INVx1_ASAP7_75t_L g16974 ( 
.A(n_16589),
.Y(n_16974)
);

AND2x2_ASAP7_75t_L g16975 ( 
.A(n_16666),
.B(n_16330),
.Y(n_16975)
);

AND2x4_ASAP7_75t_L g16976 ( 
.A(n_16575),
.B(n_16497),
.Y(n_16976)
);

NAND2xp5_ASAP7_75t_SL g16977 ( 
.A(n_16643),
.B(n_16277),
.Y(n_16977)
);

INVx1_ASAP7_75t_L g16978 ( 
.A(n_16590),
.Y(n_16978)
);

INVxp67_ASAP7_75t_L g16979 ( 
.A(n_16597),
.Y(n_16979)
);

AND2x2_ASAP7_75t_L g16980 ( 
.A(n_16686),
.B(n_16527),
.Y(n_16980)
);

AND2x2_ASAP7_75t_L g16981 ( 
.A(n_16692),
.B(n_16548),
.Y(n_16981)
);

AND2x2_ASAP7_75t_L g16982 ( 
.A(n_16649),
.B(n_16551),
.Y(n_16982)
);

NAND2xp5_ASAP7_75t_L g16983 ( 
.A(n_16574),
.B(n_16603),
.Y(n_16983)
);

INVx2_ASAP7_75t_L g16984 ( 
.A(n_16775),
.Y(n_16984)
);

INVx1_ASAP7_75t_SL g16985 ( 
.A(n_16775),
.Y(n_16985)
);

INVx1_ASAP7_75t_L g16986 ( 
.A(n_16593),
.Y(n_16986)
);

NAND2xp5_ASAP7_75t_SL g16987 ( 
.A(n_16626),
.B(n_16660),
.Y(n_16987)
);

INVx1_ASAP7_75t_L g16988 ( 
.A(n_16717),
.Y(n_16988)
);

NAND2xp5_ASAP7_75t_L g16989 ( 
.A(n_16567),
.B(n_16487),
.Y(n_16989)
);

AOI22xp5_ASAP7_75t_L g16990 ( 
.A1(n_16572),
.A2(n_16365),
.B1(n_16522),
.B2(n_16397),
.Y(n_16990)
);

INVx1_ASAP7_75t_L g16991 ( 
.A(n_16653),
.Y(n_16991)
);

AND2x2_ASAP7_75t_L g16992 ( 
.A(n_16596),
.B(n_16553),
.Y(n_16992)
);

INVx1_ASAP7_75t_L g16993 ( 
.A(n_16580),
.Y(n_16993)
);

AND2x2_ASAP7_75t_L g16994 ( 
.A(n_16639),
.B(n_16646),
.Y(n_16994)
);

INVx1_ASAP7_75t_L g16995 ( 
.A(n_16565),
.Y(n_16995)
);

NOR2x1_ASAP7_75t_L g16996 ( 
.A(n_16790),
.B(n_16418),
.Y(n_16996)
);

AOI221xp5_ASAP7_75t_L g16997 ( 
.A1(n_16616),
.A2(n_16530),
.B1(n_16502),
.B2(n_16462),
.C(n_16432),
.Y(n_16997)
);

NAND2xp5_ASAP7_75t_L g16998 ( 
.A(n_16652),
.B(n_16419),
.Y(n_16998)
);

OAI221xp5_ASAP7_75t_L g16999 ( 
.A1(n_16591),
.A2(n_16447),
.B1(n_16429),
.B2(n_16242),
.C(n_16359),
.Y(n_16999)
);

AND2x2_ASAP7_75t_L g17000 ( 
.A(n_16631),
.B(n_16408),
.Y(n_17000)
);

AND2x2_ASAP7_75t_L g17001 ( 
.A(n_16634),
.B(n_16412),
.Y(n_17001)
);

NAND4xp25_ASAP7_75t_L g17002 ( 
.A(n_16630),
.B(n_16506),
.C(n_16415),
.D(n_16482),
.Y(n_17002)
);

NAND2xp5_ASAP7_75t_SL g17003 ( 
.A(n_16668),
.B(n_16409),
.Y(n_17003)
);

NOR4xp25_ASAP7_75t_SL g17004 ( 
.A(n_16623),
.B(n_16385),
.C(n_16445),
.D(n_16405),
.Y(n_17004)
);

INVx1_ASAP7_75t_L g17005 ( 
.A(n_16564),
.Y(n_17005)
);

INVx1_ASAP7_75t_L g17006 ( 
.A(n_16655),
.Y(n_17006)
);

INVx1_ASAP7_75t_L g17007 ( 
.A(n_16823),
.Y(n_17007)
);

INVx3_ASAP7_75t_SL g17008 ( 
.A(n_16699),
.Y(n_17008)
);

NAND5xp2_ASAP7_75t_SL g17009 ( 
.A(n_16732),
.B(n_16481),
.C(n_16486),
.D(n_16498),
.E(n_16507),
.Y(n_17009)
);

AND2x2_ASAP7_75t_L g17010 ( 
.A(n_16636),
.B(n_16489),
.Y(n_17010)
);

INVx1_ASAP7_75t_L g17011 ( 
.A(n_16637),
.Y(n_17011)
);

NAND2xp5_ASAP7_75t_L g17012 ( 
.A(n_16761),
.B(n_16512),
.Y(n_17012)
);

AND2x2_ASAP7_75t_L g17013 ( 
.A(n_16662),
.B(n_16513),
.Y(n_17013)
);

INVx1_ASAP7_75t_L g17014 ( 
.A(n_16930),
.Y(n_17014)
);

NOR2xp33_ASAP7_75t_R g17015 ( 
.A(n_16605),
.B(n_16514),
.Y(n_17015)
);

OR2x2_ASAP7_75t_L g17016 ( 
.A(n_16638),
.B(n_16517),
.Y(n_17016)
);

OR2x2_ASAP7_75t_L g17017 ( 
.A(n_16601),
.B(n_16523),
.Y(n_17017)
);

NAND2xp33_ASAP7_75t_SL g17018 ( 
.A(n_16689),
.B(n_16560),
.Y(n_17018)
);

AND2x2_ASAP7_75t_L g17019 ( 
.A(n_16656),
.B(n_16217),
.Y(n_17019)
);

AND2x2_ASAP7_75t_L g17020 ( 
.A(n_16818),
.B(n_16472),
.Y(n_17020)
);

INVx1_ASAP7_75t_L g17021 ( 
.A(n_16950),
.Y(n_17021)
);

NAND2xp5_ASAP7_75t_L g17022 ( 
.A(n_16602),
.B(n_16225),
.Y(n_17022)
);

XNOR2x1_ASAP7_75t_L g17023 ( 
.A(n_16902),
.B(n_16265),
.Y(n_17023)
);

INVx1_ASAP7_75t_L g17024 ( 
.A(n_16577),
.Y(n_17024)
);

AND2x2_ASAP7_75t_L g17025 ( 
.A(n_16681),
.B(n_16349),
.Y(n_17025)
);

OAI31xp33_ASAP7_75t_L g17026 ( 
.A1(n_16613),
.A2(n_16501),
.A3(n_16402),
.B(n_16554),
.Y(n_17026)
);

NAND2xp5_ASAP7_75t_L g17027 ( 
.A(n_16618),
.B(n_16138),
.Y(n_17027)
);

NOR4xp25_ASAP7_75t_SL g17028 ( 
.A(n_16951),
.B(n_16443),
.C(n_16404),
.D(n_16469),
.Y(n_17028)
);

OR2x2_ASAP7_75t_L g17029 ( 
.A(n_16711),
.B(n_10012),
.Y(n_17029)
);

INVx2_ASAP7_75t_L g17030 ( 
.A(n_16628),
.Y(n_17030)
);

NAND2xp5_ASAP7_75t_L g17031 ( 
.A(n_16670),
.B(n_10186),
.Y(n_17031)
);

INVx4_ASAP7_75t_L g17032 ( 
.A(n_16867),
.Y(n_17032)
);

AND2x2_ASAP7_75t_L g17033 ( 
.A(n_16733),
.B(n_10187),
.Y(n_17033)
);

NAND2xp5_ASAP7_75t_L g17034 ( 
.A(n_16608),
.B(n_10187),
.Y(n_17034)
);

NAND2xp5_ASAP7_75t_L g17035 ( 
.A(n_16664),
.B(n_10187),
.Y(n_17035)
);

INVx1_ASAP7_75t_L g17036 ( 
.A(n_16909),
.Y(n_17036)
);

AND2x2_ASAP7_75t_L g17037 ( 
.A(n_16632),
.B(n_10191),
.Y(n_17037)
);

NOR2xp33_ASAP7_75t_L g17038 ( 
.A(n_16810),
.B(n_10191),
.Y(n_17038)
);

NAND2xp5_ASAP7_75t_SL g17039 ( 
.A(n_16665),
.B(n_16682),
.Y(n_17039)
);

INVxp67_ASAP7_75t_SL g17040 ( 
.A(n_16566),
.Y(n_17040)
);

OR2x2_ASAP7_75t_L g17041 ( 
.A(n_16880),
.B(n_10013),
.Y(n_17041)
);

NAND2xp33_ASAP7_75t_R g17042 ( 
.A(n_16669),
.B(n_8359),
.Y(n_17042)
);

INVx2_ASAP7_75t_L g17043 ( 
.A(n_16621),
.Y(n_17043)
);

NAND3xp33_ASAP7_75t_L g17044 ( 
.A(n_16581),
.B(n_9008),
.C(n_7870),
.Y(n_17044)
);

INVx2_ASAP7_75t_L g17045 ( 
.A(n_16697),
.Y(n_17045)
);

INVx1_ASAP7_75t_L g17046 ( 
.A(n_16744),
.Y(n_17046)
);

NOR2xp33_ASAP7_75t_L g17047 ( 
.A(n_16892),
.B(n_10191),
.Y(n_17047)
);

OR2x2_ASAP7_75t_L g17048 ( 
.A(n_16569),
.B(n_10013),
.Y(n_17048)
);

NOR3xp33_ASAP7_75t_SL g17049 ( 
.A(n_16919),
.B(n_7108),
.C(n_6990),
.Y(n_17049)
);

HB1xp67_ASAP7_75t_L g17050 ( 
.A(n_16716),
.Y(n_17050)
);

NAND2xp5_ASAP7_75t_L g17051 ( 
.A(n_16828),
.B(n_10197),
.Y(n_17051)
);

AND2x2_ASAP7_75t_L g17052 ( 
.A(n_16701),
.B(n_10197),
.Y(n_17052)
);

INVx1_ASAP7_75t_L g17053 ( 
.A(n_16746),
.Y(n_17053)
);

NAND2xp5_ASAP7_75t_L g17054 ( 
.A(n_16629),
.B(n_10197),
.Y(n_17054)
);

HB1xp67_ASAP7_75t_L g17055 ( 
.A(n_16716),
.Y(n_17055)
);

AND2x2_ASAP7_75t_L g17056 ( 
.A(n_16712),
.B(n_10205),
.Y(n_17056)
);

BUFx2_ASAP7_75t_L g17057 ( 
.A(n_16647),
.Y(n_17057)
);

INVx1_ASAP7_75t_L g17058 ( 
.A(n_16661),
.Y(n_17058)
);

AND2x2_ASAP7_75t_L g17059 ( 
.A(n_16725),
.B(n_10205),
.Y(n_17059)
);

NOR2x1_ASAP7_75t_L g17060 ( 
.A(n_16598),
.B(n_10205),
.Y(n_17060)
);

INVx1_ASAP7_75t_L g17061 ( 
.A(n_16726),
.Y(n_17061)
);

NOR3xp33_ASAP7_75t_SL g17062 ( 
.A(n_16568),
.B(n_7108),
.C(n_6959),
.Y(n_17062)
);

AND2x2_ASAP7_75t_L g17063 ( 
.A(n_16751),
.B(n_10212),
.Y(n_17063)
);

BUFx2_ASAP7_75t_L g17064 ( 
.A(n_16647),
.Y(n_17064)
);

OR2x2_ASAP7_75t_L g17065 ( 
.A(n_16786),
.B(n_10015),
.Y(n_17065)
);

INVx2_ASAP7_75t_L g17066 ( 
.A(n_16794),
.Y(n_17066)
);

OR2x2_ASAP7_75t_L g17067 ( 
.A(n_16927),
.B(n_10015),
.Y(n_17067)
);

NOR2xp33_ASAP7_75t_L g17068 ( 
.A(n_16846),
.B(n_10212),
.Y(n_17068)
);

OAI21xp33_ASAP7_75t_L g17069 ( 
.A1(n_16687),
.A2(n_8722),
.B(n_8717),
.Y(n_17069)
);

NAND2x1_ASAP7_75t_SL g17070 ( 
.A(n_16837),
.B(n_10314),
.Y(n_17070)
);

INVx1_ASAP7_75t_L g17071 ( 
.A(n_16838),
.Y(n_17071)
);

OAI211xp5_ASAP7_75t_SL g17072 ( 
.A1(n_16815),
.A2(n_7768),
.B(n_8022),
.C(n_7917),
.Y(n_17072)
);

INVx1_ASAP7_75t_L g17073 ( 
.A(n_16570),
.Y(n_17073)
);

OR2x2_ASAP7_75t_L g17074 ( 
.A(n_16758),
.B(n_10016),
.Y(n_17074)
);

NOR2xp67_ASAP7_75t_L g17075 ( 
.A(n_16710),
.B(n_16811),
.Y(n_17075)
);

INVx1_ASAP7_75t_L g17076 ( 
.A(n_16690),
.Y(n_17076)
);

INVx1_ASAP7_75t_SL g17077 ( 
.A(n_16926),
.Y(n_17077)
);

OAI211xp5_ASAP7_75t_L g17078 ( 
.A1(n_16562),
.A2(n_9691),
.B(n_9728),
.C(n_9724),
.Y(n_17078)
);

NAND2xp5_ASAP7_75t_L g17079 ( 
.A(n_16941),
.B(n_10212),
.Y(n_17079)
);

INVx2_ASAP7_75t_L g17080 ( 
.A(n_16802),
.Y(n_17080)
);

OAI22xp5_ASAP7_75t_L g17081 ( 
.A1(n_16578),
.A2(n_10218),
.B1(n_10230),
.B2(n_10226),
.Y(n_17081)
);

INVx1_ASAP7_75t_L g17082 ( 
.A(n_16848),
.Y(n_17082)
);

NAND2xp5_ASAP7_75t_L g17083 ( 
.A(n_16895),
.B(n_10218),
.Y(n_17083)
);

INVx1_ASAP7_75t_L g17084 ( 
.A(n_16648),
.Y(n_17084)
);

INVx1_ASAP7_75t_L g17085 ( 
.A(n_16676),
.Y(n_17085)
);

INVx2_ASAP7_75t_SL g17086 ( 
.A(n_16847),
.Y(n_17086)
);

INVx1_ASAP7_75t_L g17087 ( 
.A(n_16743),
.Y(n_17087)
);

OR2x4_ASAP7_75t_L g17088 ( 
.A(n_16745),
.B(n_9008),
.Y(n_17088)
);

NAND2xp5_ASAP7_75t_L g17089 ( 
.A(n_16752),
.B(n_10218),
.Y(n_17089)
);

NOR2xp33_ASAP7_75t_L g17090 ( 
.A(n_16729),
.B(n_10226),
.Y(n_17090)
);

BUFx4f_ASAP7_75t_SL g17091 ( 
.A(n_16763),
.Y(n_17091)
);

NAND2xp5_ASAP7_75t_SL g17092 ( 
.A(n_16635),
.B(n_9008),
.Y(n_17092)
);

NAND2xp5_ASAP7_75t_L g17093 ( 
.A(n_16753),
.B(n_10226),
.Y(n_17093)
);

OR2x2_ASAP7_75t_L g17094 ( 
.A(n_16757),
.B(n_10016),
.Y(n_17094)
);

NAND2x1p5_ASAP7_75t_L g17095 ( 
.A(n_16845),
.B(n_9781),
.Y(n_17095)
);

NAND3xp33_ASAP7_75t_L g17096 ( 
.A(n_16606),
.B(n_7870),
.C(n_7711),
.Y(n_17096)
);

HB1xp67_ASAP7_75t_L g17097 ( 
.A(n_16749),
.Y(n_17097)
);

NOR2x1_ASAP7_75t_L g17098 ( 
.A(n_16798),
.B(n_10230),
.Y(n_17098)
);

INVx1_ASAP7_75t_L g17099 ( 
.A(n_16600),
.Y(n_17099)
);

NAND2xp5_ASAP7_75t_SL g17100 ( 
.A(n_16640),
.B(n_7711),
.Y(n_17100)
);

INVx5_ASAP7_75t_L g17101 ( 
.A(n_16871),
.Y(n_17101)
);

NAND2xp33_ASAP7_75t_SL g17102 ( 
.A(n_16595),
.B(n_6648),
.Y(n_17102)
);

INVx1_ASAP7_75t_L g17103 ( 
.A(n_16819),
.Y(n_17103)
);

NOR4xp25_ASAP7_75t_SL g17104 ( 
.A(n_16868),
.B(n_10019),
.C(n_10020),
.D(n_10018),
.Y(n_17104)
);

HB1xp67_ASAP7_75t_L g17105 ( 
.A(n_16749),
.Y(n_17105)
);

AND2x4_ASAP7_75t_SL g17106 ( 
.A(n_16817),
.B(n_7272),
.Y(n_17106)
);

INVx1_ASAP7_75t_L g17107 ( 
.A(n_16822),
.Y(n_17107)
);

HB1xp67_ASAP7_75t_L g17108 ( 
.A(n_16959),
.Y(n_17108)
);

AOI21xp5_ASAP7_75t_L g17109 ( 
.A1(n_16840),
.A2(n_10242),
.B(n_10230),
.Y(n_17109)
);

AOI33xp33_ASAP7_75t_L g17110 ( 
.A1(n_16905),
.A2(n_8274),
.A3(n_8103),
.B1(n_8311),
.B2(n_8228),
.B3(n_8085),
.Y(n_17110)
);

NOR2xp33_ASAP7_75t_SL g17111 ( 
.A(n_16851),
.B(n_8228),
.Y(n_17111)
);

INVx2_ASAP7_75t_L g17112 ( 
.A(n_16875),
.Y(n_17112)
);

INVx1_ASAP7_75t_L g17113 ( 
.A(n_16713),
.Y(n_17113)
);

INVx1_ASAP7_75t_L g17114 ( 
.A(n_16718),
.Y(n_17114)
);

OAI211xp5_ASAP7_75t_SL g17115 ( 
.A1(n_16707),
.A2(n_7917),
.B(n_8038),
.C(n_8022),
.Y(n_17115)
);

INVx1_ASAP7_75t_SL g17116 ( 
.A(n_16588),
.Y(n_17116)
);

OR2x2_ASAP7_75t_L g17117 ( 
.A(n_16720),
.B(n_10018),
.Y(n_17117)
);

INVx1_ASAP7_75t_L g17118 ( 
.A(n_16723),
.Y(n_17118)
);

OR2x2_ASAP7_75t_L g17119 ( 
.A(n_16727),
.B(n_10019),
.Y(n_17119)
);

INVx1_ASAP7_75t_SL g17120 ( 
.A(n_16842),
.Y(n_17120)
);

AND2x4_ASAP7_75t_SL g17121 ( 
.A(n_16777),
.B(n_7272),
.Y(n_17121)
);

INVx1_ASAP7_75t_L g17122 ( 
.A(n_16736),
.Y(n_17122)
);

INVx1_ASAP7_75t_L g17123 ( 
.A(n_16614),
.Y(n_17123)
);

NAND2xp5_ASAP7_75t_L g17124 ( 
.A(n_16877),
.B(n_16953),
.Y(n_17124)
);

INVx1_ASAP7_75t_L g17125 ( 
.A(n_16958),
.Y(n_17125)
);

NAND2xp33_ASAP7_75t_R g17126 ( 
.A(n_16820),
.B(n_8359),
.Y(n_17126)
);

INVx1_ASAP7_75t_SL g17127 ( 
.A(n_16839),
.Y(n_17127)
);

INVx2_ASAP7_75t_L g17128 ( 
.A(n_16760),
.Y(n_17128)
);

INVx1_ASAP7_75t_L g17129 ( 
.A(n_16583),
.Y(n_17129)
);

INVxp67_ASAP7_75t_SL g17130 ( 
.A(n_16715),
.Y(n_17130)
);

INVx2_ASAP7_75t_L g17131 ( 
.A(n_16896),
.Y(n_17131)
);

INVx2_ASAP7_75t_L g17132 ( 
.A(n_16893),
.Y(n_17132)
);

NAND2xp5_ASAP7_75t_L g17133 ( 
.A(n_16764),
.B(n_10242),
.Y(n_17133)
);

NAND2xp5_ASAP7_75t_L g17134 ( 
.A(n_16901),
.B(n_10242),
.Y(n_17134)
);

AND2x2_ASAP7_75t_L g17135 ( 
.A(n_16671),
.B(n_10244),
.Y(n_17135)
);

INVx2_ASAP7_75t_L g17136 ( 
.A(n_16916),
.Y(n_17136)
);

AND2x2_ASAP7_75t_L g17137 ( 
.A(n_16739),
.B(n_10244),
.Y(n_17137)
);

INVx2_ASAP7_75t_L g17138 ( 
.A(n_16938),
.Y(n_17138)
);

NAND2xp5_ASAP7_75t_L g17139 ( 
.A(n_16947),
.B(n_10244),
.Y(n_17139)
);

OR2x2_ASAP7_75t_L g17140 ( 
.A(n_16949),
.B(n_10020),
.Y(n_17140)
);

AND2x2_ASAP7_75t_L g17141 ( 
.A(n_16731),
.B(n_10247),
.Y(n_17141)
);

AND2x2_ASAP7_75t_L g17142 ( 
.A(n_16765),
.B(n_16767),
.Y(n_17142)
);

AND2x2_ASAP7_75t_L g17143 ( 
.A(n_16783),
.B(n_10247),
.Y(n_17143)
);

AND2x2_ASAP7_75t_L g17144 ( 
.A(n_16735),
.B(n_10247),
.Y(n_17144)
);

INVx2_ASAP7_75t_L g17145 ( 
.A(n_16627),
.Y(n_17145)
);

AND2x2_ASAP7_75t_L g17146 ( 
.A(n_16709),
.B(n_16673),
.Y(n_17146)
);

HB1xp67_ASAP7_75t_L g17147 ( 
.A(n_16959),
.Y(n_17147)
);

INVx1_ASAP7_75t_L g17148 ( 
.A(n_16833),
.Y(n_17148)
);

INVx2_ASAP7_75t_L g17149 ( 
.A(n_16579),
.Y(n_17149)
);

INVx1_ASAP7_75t_L g17150 ( 
.A(n_16738),
.Y(n_17150)
);

NAND2xp33_ASAP7_75t_SL g17151 ( 
.A(n_16843),
.B(n_6648),
.Y(n_17151)
);

AND2x2_ASAP7_75t_L g17152 ( 
.A(n_16695),
.B(n_10249),
.Y(n_17152)
);

INVx2_ASAP7_75t_SL g17153 ( 
.A(n_16962),
.Y(n_17153)
);

INVxp67_ASAP7_75t_L g17154 ( 
.A(n_16683),
.Y(n_17154)
);

AND2x2_ASAP7_75t_L g17155 ( 
.A(n_16776),
.B(n_16778),
.Y(n_17155)
);

INVx1_ASAP7_75t_L g17156 ( 
.A(n_16779),
.Y(n_17156)
);

NAND2xp33_ASAP7_75t_R g17157 ( 
.A(n_16854),
.B(n_8359),
.Y(n_17157)
);

INVx2_ASAP7_75t_L g17158 ( 
.A(n_16756),
.Y(n_17158)
);

NOR2x1_ASAP7_75t_L g17159 ( 
.A(n_16804),
.B(n_10249),
.Y(n_17159)
);

NOR3xp33_ASAP7_75t_L g17160 ( 
.A(n_16850),
.B(n_16734),
.C(n_16714),
.Y(n_17160)
);

NAND2xp5_ASAP7_75t_L g17161 ( 
.A(n_16827),
.B(n_10249),
.Y(n_17161)
);

INVx1_ASAP7_75t_L g17162 ( 
.A(n_16771),
.Y(n_17162)
);

INVx1_ASAP7_75t_L g17163 ( 
.A(n_16625),
.Y(n_17163)
);

INVx2_ASAP7_75t_L g17164 ( 
.A(n_16964),
.Y(n_17164)
);

NOR2x1_ASAP7_75t_L g17165 ( 
.A(n_16813),
.B(n_10258),
.Y(n_17165)
);

HB1xp67_ASAP7_75t_L g17166 ( 
.A(n_16844),
.Y(n_17166)
);

INVx2_ASAP7_75t_L g17167 ( 
.A(n_16964),
.Y(n_17167)
);

INVx1_ASAP7_75t_L g17168 ( 
.A(n_16609),
.Y(n_17168)
);

NAND2xp5_ASAP7_75t_L g17169 ( 
.A(n_16641),
.B(n_10258),
.Y(n_17169)
);

NOR4xp25_ASAP7_75t_SL g17170 ( 
.A(n_16934),
.B(n_10023),
.C(n_10029),
.D(n_10021),
.Y(n_17170)
);

NAND3xp33_ASAP7_75t_SL g17171 ( 
.A(n_16857),
.B(n_8323),
.C(n_8293),
.Y(n_17171)
);

NAND2xp5_ASAP7_75t_L g17172 ( 
.A(n_16904),
.B(n_10258),
.Y(n_17172)
);

OR2x2_ASAP7_75t_L g17173 ( 
.A(n_16587),
.B(n_16685),
.Y(n_17173)
);

AND2x2_ASAP7_75t_L g17174 ( 
.A(n_16703),
.B(n_10262),
.Y(n_17174)
);

AND2x2_ASAP7_75t_L g17175 ( 
.A(n_16696),
.B(n_10262),
.Y(n_17175)
);

HB1xp67_ASAP7_75t_L g17176 ( 
.A(n_16816),
.Y(n_17176)
);

NAND2xp5_ASAP7_75t_L g17177 ( 
.A(n_16841),
.B(n_10262),
.Y(n_17177)
);

NAND2xp5_ASAP7_75t_L g17178 ( 
.A(n_16747),
.B(n_10264),
.Y(n_17178)
);

AND2x2_ASAP7_75t_L g17179 ( 
.A(n_16859),
.B(n_10264),
.Y(n_17179)
);

OR2x2_ASAP7_75t_L g17180 ( 
.A(n_16620),
.B(n_10021),
.Y(n_17180)
);

AND2x2_ASAP7_75t_L g17181 ( 
.A(n_16754),
.B(n_10264),
.Y(n_17181)
);

INVx1_ASAP7_75t_L g17182 ( 
.A(n_16582),
.Y(n_17182)
);

AND2x2_ASAP7_75t_L g17183 ( 
.A(n_16780),
.B(n_10266),
.Y(n_17183)
);

INVx2_ASAP7_75t_L g17184 ( 
.A(n_16869),
.Y(n_17184)
);

NAND2xp5_ASAP7_75t_L g17185 ( 
.A(n_16785),
.B(n_10266),
.Y(n_17185)
);

INVx1_ASAP7_75t_L g17186 ( 
.A(n_16657),
.Y(n_17186)
);

INVx1_ASAP7_75t_L g17187 ( 
.A(n_16611),
.Y(n_17187)
);

NAND3xp33_ASAP7_75t_L g17188 ( 
.A(n_16824),
.B(n_7870),
.C(n_7711),
.Y(n_17188)
);

OR2x2_ASAP7_75t_L g17189 ( 
.A(n_16706),
.B(n_10023),
.Y(n_17189)
);

AND2x2_ASAP7_75t_L g17190 ( 
.A(n_16898),
.B(n_10266),
.Y(n_17190)
);

OR2x2_ASAP7_75t_L g17191 ( 
.A(n_16619),
.B(n_10029),
.Y(n_17191)
);

INVx2_ASAP7_75t_L g17192 ( 
.A(n_16870),
.Y(n_17192)
);

BUFx2_ASAP7_75t_L g17193 ( 
.A(n_16945),
.Y(n_17193)
);

AND2x2_ASAP7_75t_L g17194 ( 
.A(n_16874),
.B(n_10267),
.Y(n_17194)
);

AND2x2_ASAP7_75t_SL g17195 ( 
.A(n_16853),
.B(n_8359),
.Y(n_17195)
);

AND2x2_ASAP7_75t_L g17196 ( 
.A(n_16633),
.B(n_10267),
.Y(n_17196)
);

AND2x2_ASAP7_75t_L g17197 ( 
.A(n_16939),
.B(n_10267),
.Y(n_17197)
);

BUFx2_ASAP7_75t_SL g17198 ( 
.A(n_16882),
.Y(n_17198)
);

INVx2_ASAP7_75t_L g17199 ( 
.A(n_16881),
.Y(n_17199)
);

INVx1_ASAP7_75t_SL g17200 ( 
.A(n_16722),
.Y(n_17200)
);

AND2x2_ASAP7_75t_L g17201 ( 
.A(n_16966),
.B(n_10283),
.Y(n_17201)
);

NAND2xp33_ASAP7_75t_R g17202 ( 
.A(n_16885),
.B(n_8405),
.Y(n_17202)
);

AND2x2_ASAP7_75t_L g17203 ( 
.A(n_16759),
.B(n_10283),
.Y(n_17203)
);

NAND2xp5_ASAP7_75t_L g17204 ( 
.A(n_16862),
.B(n_10283),
.Y(n_17204)
);

INVx1_ASAP7_75t_L g17205 ( 
.A(n_16825),
.Y(n_17205)
);

NAND2xp5_ASAP7_75t_L g17206 ( 
.A(n_16864),
.B(n_16876),
.Y(n_17206)
);

NOR2xp33_ASAP7_75t_L g17207 ( 
.A(n_16928),
.B(n_10287),
.Y(n_17207)
);

OR2x2_ASAP7_75t_L g17208 ( 
.A(n_16584),
.B(n_10032),
.Y(n_17208)
);

NAND3xp33_ASAP7_75t_L g17209 ( 
.A(n_16762),
.B(n_7870),
.C(n_7711),
.Y(n_17209)
);

INVx2_ASAP7_75t_L g17210 ( 
.A(n_16849),
.Y(n_17210)
);

INVx1_ASAP7_75t_L g17211 ( 
.A(n_16667),
.Y(n_17211)
);

NOR2x1_ASAP7_75t_L g17212 ( 
.A(n_16906),
.B(n_10287),
.Y(n_17212)
);

AND2x2_ASAP7_75t_L g17213 ( 
.A(n_16910),
.B(n_10287),
.Y(n_17213)
);

NAND2xp5_ASAP7_75t_L g17214 ( 
.A(n_16913),
.B(n_10291),
.Y(n_17214)
);

NAND2x1p5_ASAP7_75t_L g17215 ( 
.A(n_16914),
.B(n_9781),
.Y(n_17215)
);

INVx2_ASAP7_75t_L g17216 ( 
.A(n_16889),
.Y(n_17216)
);

INVx1_ASAP7_75t_L g17217 ( 
.A(n_16766),
.Y(n_17217)
);

AND2x2_ASAP7_75t_L g17218 ( 
.A(n_16920),
.B(n_10291),
.Y(n_17218)
);

NOR3xp33_ASAP7_75t_L g17219 ( 
.A(n_16872),
.B(n_9811),
.C(n_9793),
.Y(n_17219)
);

INVx1_ASAP7_75t_L g17220 ( 
.A(n_16672),
.Y(n_17220)
);

AND2x2_ASAP7_75t_L g17221 ( 
.A(n_16924),
.B(n_10291),
.Y(n_17221)
);

NAND5xp2_ASAP7_75t_SL g17222 ( 
.A(n_16693),
.B(n_8903),
.C(n_9811),
.D(n_9793),
.E(n_9866),
.Y(n_17222)
);

OAI21xp33_ASAP7_75t_L g17223 ( 
.A1(n_16592),
.A2(n_8731),
.B(n_8722),
.Y(n_17223)
);

INVx1_ASAP7_75t_L g17224 ( 
.A(n_16585),
.Y(n_17224)
);

NAND2xp5_ASAP7_75t_L g17225 ( 
.A(n_16933),
.B(n_10298),
.Y(n_17225)
);

AOI21xp33_ASAP7_75t_SL g17226 ( 
.A1(n_16795),
.A2(n_9943),
.B(n_9866),
.Y(n_17226)
);

NOR2x1_ASAP7_75t_L g17227 ( 
.A(n_16936),
.B(n_10298),
.Y(n_17227)
);

NOR2xp33_ASAP7_75t_L g17228 ( 
.A(n_16937),
.B(n_10298),
.Y(n_17228)
);

OR2x2_ASAP7_75t_L g17229 ( 
.A(n_16866),
.B(n_10032),
.Y(n_17229)
);

NOR3xp33_ASAP7_75t_L g17230 ( 
.A(n_16940),
.B(n_10014),
.C(n_9943),
.Y(n_17230)
);

HB1xp67_ASAP7_75t_L g17231 ( 
.A(n_16617),
.Y(n_17231)
);

NOR3xp33_ASAP7_75t_L g17232 ( 
.A(n_16955),
.B(n_10028),
.C(n_10014),
.Y(n_17232)
);

OR2x2_ASAP7_75t_L g17233 ( 
.A(n_16650),
.B(n_10035),
.Y(n_17233)
);

NAND2xp5_ASAP7_75t_L g17234 ( 
.A(n_16956),
.B(n_10305),
.Y(n_17234)
);

AND2x2_ASAP7_75t_L g17235 ( 
.A(n_16728),
.B(n_10305),
.Y(n_17235)
);

INVx1_ASAP7_75t_L g17236 ( 
.A(n_16799),
.Y(n_17236)
);

AND2x2_ASAP7_75t_L g17237 ( 
.A(n_16957),
.B(n_10305),
.Y(n_17237)
);

INVx1_ASAP7_75t_L g17238 ( 
.A(n_16705),
.Y(n_17238)
);

NAND2xp5_ASAP7_75t_L g17239 ( 
.A(n_16960),
.B(n_10311),
.Y(n_17239)
);

INVx2_ASAP7_75t_SL g17240 ( 
.A(n_16834),
.Y(n_17240)
);

INVx2_ASAP7_75t_L g17241 ( 
.A(n_16903),
.Y(n_17241)
);

NAND2xp5_ASAP7_75t_L g17242 ( 
.A(n_16963),
.B(n_10311),
.Y(n_17242)
);

INVx2_ASAP7_75t_L g17243 ( 
.A(n_16879),
.Y(n_17243)
);

INVx1_ASAP7_75t_L g17244 ( 
.A(n_16730),
.Y(n_17244)
);

INVx1_ASAP7_75t_L g17245 ( 
.A(n_16644),
.Y(n_17245)
);

HB1xp67_ASAP7_75t_L g17246 ( 
.A(n_16792),
.Y(n_17246)
);

AND2x2_ASAP7_75t_L g17247 ( 
.A(n_16651),
.B(n_10311),
.Y(n_17247)
);

INVx1_ASAP7_75t_L g17248 ( 
.A(n_16680),
.Y(n_17248)
);

INVx1_ASAP7_75t_L g17249 ( 
.A(n_16675),
.Y(n_17249)
);

AND2x2_ASAP7_75t_L g17250 ( 
.A(n_16654),
.B(n_10318),
.Y(n_17250)
);

AOI22xp33_ASAP7_75t_L g17251 ( 
.A1(n_16684),
.A2(n_8536),
.B1(n_7870),
.B2(n_7711),
.Y(n_17251)
);

INVx1_ASAP7_75t_L g17252 ( 
.A(n_16769),
.Y(n_17252)
);

NAND2xp33_ASAP7_75t_SL g17253 ( 
.A(n_16944),
.B(n_6757),
.Y(n_17253)
);

AND2x2_ASAP7_75t_L g17254 ( 
.A(n_16679),
.B(n_10318),
.Y(n_17254)
);

OR2x2_ASAP7_75t_L g17255 ( 
.A(n_16917),
.B(n_10035),
.Y(n_17255)
);

OR2x2_ASAP7_75t_L g17256 ( 
.A(n_16791),
.B(n_10042),
.Y(n_17256)
);

NAND2xp5_ASAP7_75t_L g17257 ( 
.A(n_16911),
.B(n_10318),
.Y(n_17257)
);

NAND2xp5_ASAP7_75t_L g17258 ( 
.A(n_16886),
.B(n_10319),
.Y(n_17258)
);

OAI221xp5_ASAP7_75t_L g17259 ( 
.A1(n_16891),
.A2(n_8274),
.B1(n_8334),
.B2(n_8318),
.C(n_8311),
.Y(n_17259)
);

CKINVDCx5p33_ASAP7_75t_R g17260 ( 
.A(n_16741),
.Y(n_17260)
);

NOR2xp33_ASAP7_75t_L g17261 ( 
.A(n_16894),
.B(n_10319),
.Y(n_17261)
);

INVx1_ASAP7_75t_L g17262 ( 
.A(n_16805),
.Y(n_17262)
);

AOI22xp33_ASAP7_75t_L g17263 ( 
.A1(n_16806),
.A2(n_8536),
.B1(n_7711),
.B2(n_8903),
.Y(n_17263)
);

INVx1_ASAP7_75t_L g17264 ( 
.A(n_16808),
.Y(n_17264)
);

INVx1_ASAP7_75t_L g17265 ( 
.A(n_16773),
.Y(n_17265)
);

CKINVDCx16_ASAP7_75t_R g17266 ( 
.A(n_16886),
.Y(n_17266)
);

INVx1_ASAP7_75t_L g17267 ( 
.A(n_16887),
.Y(n_17267)
);

INVx1_ASAP7_75t_L g17268 ( 
.A(n_16887),
.Y(n_17268)
);

OAI31xp33_ASAP7_75t_L g17269 ( 
.A1(n_16688),
.A2(n_8334),
.A3(n_8353),
.B(n_8318),
.Y(n_17269)
);

INVx2_ASAP7_75t_L g17270 ( 
.A(n_16931),
.Y(n_17270)
);

NAND3xp33_ASAP7_75t_L g17271 ( 
.A(n_16694),
.B(n_8405),
.C(n_8550),
.Y(n_17271)
);

AND2x4_ASAP7_75t_L g17272 ( 
.A(n_16607),
.B(n_10028),
.Y(n_17272)
);

INVx1_ASAP7_75t_L g17273 ( 
.A(n_16803),
.Y(n_17273)
);

AND2x2_ASAP7_75t_L g17274 ( 
.A(n_16768),
.B(n_10319),
.Y(n_17274)
);

INVx2_ASAP7_75t_L g17275 ( 
.A(n_16796),
.Y(n_17275)
);

BUFx3_ASAP7_75t_L g17276 ( 
.A(n_16594),
.Y(n_17276)
);

NAND2xp5_ASAP7_75t_L g17277 ( 
.A(n_16921),
.B(n_10320),
.Y(n_17277)
);

NAND2xp5_ASAP7_75t_SL g17278 ( 
.A(n_16573),
.B(n_10056),
.Y(n_17278)
);

AND2x2_ASAP7_75t_L g17279 ( 
.A(n_16645),
.B(n_10320),
.Y(n_17279)
);

INVx1_ASAP7_75t_L g17280 ( 
.A(n_16856),
.Y(n_17280)
);

INVx1_ASAP7_75t_L g17281 ( 
.A(n_16890),
.Y(n_17281)
);

INVxp67_ASAP7_75t_L g17282 ( 
.A(n_16831),
.Y(n_17282)
);

AND2x2_ASAP7_75t_SL g17283 ( 
.A(n_16719),
.B(n_8405),
.Y(n_17283)
);

NAND2xp5_ASAP7_75t_L g17284 ( 
.A(n_16832),
.B(n_10320),
.Y(n_17284)
);

AOI22xp33_ASAP7_75t_L g17285 ( 
.A1(n_16748),
.A2(n_8536),
.B1(n_8903),
.B2(n_8501),
.Y(n_17285)
);

OR2x2_ASAP7_75t_L g17286 ( 
.A(n_16922),
.B(n_10042),
.Y(n_17286)
);

INVx1_ASAP7_75t_L g17287 ( 
.A(n_16929),
.Y(n_17287)
);

OR2x2_ASAP7_75t_L g17288 ( 
.A(n_16932),
.B(n_10047),
.Y(n_17288)
);

AND2x2_ASAP7_75t_L g17289 ( 
.A(n_16935),
.B(n_10322),
.Y(n_17289)
);

AND2x2_ASAP7_75t_SL g17290 ( 
.A(n_16770),
.B(n_16912),
.Y(n_17290)
);

OAI221xp5_ASAP7_75t_L g17291 ( 
.A1(n_16772),
.A2(n_8318),
.B1(n_8357),
.B2(n_8353),
.C(n_8334),
.Y(n_17291)
);

CKINVDCx16_ASAP7_75t_R g17292 ( 
.A(n_16700),
.Y(n_17292)
);

NOR2xp33_ASAP7_75t_L g17293 ( 
.A(n_16836),
.B(n_10322),
.Y(n_17293)
);

NAND2xp5_ASAP7_75t_L g17294 ( 
.A(n_16952),
.B(n_10322),
.Y(n_17294)
);

NAND2xp33_ASAP7_75t_SL g17295 ( 
.A(n_16954),
.B(n_16965),
.Y(n_17295)
);

INVx1_ASAP7_75t_L g17296 ( 
.A(n_16942),
.Y(n_17296)
);

INVx2_ASAP7_75t_SL g17297 ( 
.A(n_16946),
.Y(n_17297)
);

INVx1_ASAP7_75t_L g17298 ( 
.A(n_16967),
.Y(n_17298)
);

INVxp67_ASAP7_75t_L g17299 ( 
.A(n_16801),
.Y(n_17299)
);

NAND2xp5_ASAP7_75t_L g17300 ( 
.A(n_16800),
.B(n_10323),
.Y(n_17300)
);

OR2x2_ASAP7_75t_L g17301 ( 
.A(n_16861),
.B(n_10047),
.Y(n_17301)
);

AND2x2_ASAP7_75t_L g17302 ( 
.A(n_16826),
.B(n_10323),
.Y(n_17302)
);

OAI31xp33_ASAP7_75t_SL g17303 ( 
.A1(n_16774),
.A2(n_10092),
.A3(n_10151),
.B(n_10056),
.Y(n_17303)
);

INVxp33_ASAP7_75t_SL g17304 ( 
.A(n_16721),
.Y(n_17304)
);

AND2x2_ASAP7_75t_L g17305 ( 
.A(n_16943),
.B(n_10323),
.Y(n_17305)
);

INVx1_ASAP7_75t_L g17306 ( 
.A(n_16835),
.Y(n_17306)
);

AND2x2_ASAP7_75t_L g17307 ( 
.A(n_16918),
.B(n_16807),
.Y(n_17307)
);

AND2x4_ASAP7_75t_L g17308 ( 
.A(n_16812),
.B(n_16814),
.Y(n_17308)
);

NAND2xp5_ASAP7_75t_L g17309 ( 
.A(n_16642),
.B(n_10327),
.Y(n_17309)
);

INVx1_ASAP7_75t_L g17310 ( 
.A(n_16788),
.Y(n_17310)
);

NAND2xp5_ASAP7_75t_L g17311 ( 
.A(n_16698),
.B(n_10327),
.Y(n_17311)
);

AND2x2_ASAP7_75t_L g17312 ( 
.A(n_16888),
.B(n_10327),
.Y(n_17312)
);

NAND2x1_ASAP7_75t_L g17313 ( 
.A(n_16674),
.B(n_10332),
.Y(n_17313)
);

NAND2xp5_ASAP7_75t_L g17314 ( 
.A(n_16599),
.B(n_10332),
.Y(n_17314)
);

AOI31xp33_ASAP7_75t_L g17315 ( 
.A1(n_16797),
.A2(n_8323),
.A3(n_8366),
.B(n_8293),
.Y(n_17315)
);

NAND2xp5_ASAP7_75t_L g17316 ( 
.A(n_16678),
.B(n_10332),
.Y(n_17316)
);

OR2x2_ASAP7_75t_L g17317 ( 
.A(n_16923),
.B(n_10053),
.Y(n_17317)
);

AND2x2_ASAP7_75t_L g17318 ( 
.A(n_16852),
.B(n_10349),
.Y(n_17318)
);

AND2x2_ASAP7_75t_L g17319 ( 
.A(n_16855),
.B(n_10349),
.Y(n_17319)
);

INVx2_ASAP7_75t_L g17320 ( 
.A(n_16674),
.Y(n_17320)
);

INVx1_ASAP7_75t_L g17321 ( 
.A(n_16576),
.Y(n_17321)
);

NOR2x1_ASAP7_75t_L g17322 ( 
.A(n_16615),
.B(n_16708),
.Y(n_17322)
);

INVx1_ASAP7_75t_L g17323 ( 
.A(n_16750),
.Y(n_17323)
);

AND2x2_ASAP7_75t_L g17324 ( 
.A(n_16873),
.B(n_10349),
.Y(n_17324)
);

HB1xp67_ASAP7_75t_L g17325 ( 
.A(n_16781),
.Y(n_17325)
);

INVx3_ASAP7_75t_SL g17326 ( 
.A(n_16789),
.Y(n_17326)
);

OR2x2_ASAP7_75t_L g17327 ( 
.A(n_16968),
.B(n_10053),
.Y(n_17327)
);

AND2x2_ASAP7_75t_L g17328 ( 
.A(n_16586),
.B(n_10351),
.Y(n_17328)
);

AND2x2_ASAP7_75t_L g17329 ( 
.A(n_16691),
.B(n_10351),
.Y(n_17329)
);

NAND3xp33_ASAP7_75t_L g17330 ( 
.A(n_16787),
.B(n_8405),
.C(n_8550),
.Y(n_17330)
);

HB1xp67_ASAP7_75t_L g17331 ( 
.A(n_16789),
.Y(n_17331)
);

AND2x2_ASAP7_75t_L g17332 ( 
.A(n_16624),
.B(n_10351),
.Y(n_17332)
);

INVx1_ASAP7_75t_L g17333 ( 
.A(n_16948),
.Y(n_17333)
);

NAND2xp5_ASAP7_75t_L g17334 ( 
.A(n_16610),
.B(n_10357),
.Y(n_17334)
);

INVxp67_ASAP7_75t_L g17335 ( 
.A(n_16830),
.Y(n_17335)
);

OR2x2_ASAP7_75t_L g17336 ( 
.A(n_16737),
.B(n_10059),
.Y(n_17336)
);

INVxp67_ASAP7_75t_L g17337 ( 
.A(n_16829),
.Y(n_17337)
);

NAND2xp5_ASAP7_75t_L g17338 ( 
.A(n_16610),
.B(n_10357),
.Y(n_17338)
);

AND2x2_ASAP7_75t_L g17339 ( 
.A(n_16624),
.B(n_10357),
.Y(n_17339)
);

CKINVDCx16_ASAP7_75t_R g17340 ( 
.A(n_16908),
.Y(n_17340)
);

AND2x4_ASAP7_75t_L g17341 ( 
.A(n_16677),
.B(n_16899),
.Y(n_17341)
);

NAND2xp5_ASAP7_75t_L g17342 ( 
.A(n_16702),
.B(n_10358),
.Y(n_17342)
);

INVx5_ASAP7_75t_L g17343 ( 
.A(n_16677),
.Y(n_17343)
);

NOR2xp33_ASAP7_75t_L g17344 ( 
.A(n_16784),
.B(n_10358),
.Y(n_17344)
);

AND2x2_ASAP7_75t_L g17345 ( 
.A(n_16860),
.B(n_10358),
.Y(n_17345)
);

INVx1_ASAP7_75t_L g17346 ( 
.A(n_16659),
.Y(n_17346)
);

AND2x4_ASAP7_75t_L g17347 ( 
.A(n_16884),
.B(n_10367),
.Y(n_17347)
);

NAND3xp33_ASAP7_75t_SL g17348 ( 
.A(n_16915),
.B(n_16782),
.C(n_16793),
.Y(n_17348)
);

INVxp67_ASAP7_75t_SL g17349 ( 
.A(n_16961),
.Y(n_17349)
);

NAND4xp25_ASAP7_75t_L g17350 ( 
.A(n_16821),
.B(n_8755),
.C(n_8800),
.D(n_8731),
.Y(n_17350)
);

AND2x2_ASAP7_75t_L g17351 ( 
.A(n_16755),
.B(n_10367),
.Y(n_17351)
);

NAND4xp25_ASAP7_75t_L g17352 ( 
.A(n_16883),
.B(n_8755),
.C(n_8800),
.D(n_8731),
.Y(n_17352)
);

NAND2xp5_ASAP7_75t_L g17353 ( 
.A(n_16724),
.B(n_10367),
.Y(n_17353)
);

INVx1_ASAP7_75t_L g17354 ( 
.A(n_16740),
.Y(n_17354)
);

OR2x2_ASAP7_75t_L g17355 ( 
.A(n_16897),
.B(n_10059),
.Y(n_17355)
);

INVx1_ASAP7_75t_L g17356 ( 
.A(n_16571),
.Y(n_17356)
);

INVx1_ASAP7_75t_SL g17357 ( 
.A(n_17008),
.Y(n_17357)
);

AND2x2_ASAP7_75t_L g17358 ( 
.A(n_16975),
.B(n_16925),
.Y(n_17358)
);

AND2x2_ASAP7_75t_L g17359 ( 
.A(n_16976),
.B(n_16809),
.Y(n_17359)
);

INVx2_ASAP7_75t_L g17360 ( 
.A(n_17101),
.Y(n_17360)
);

INVx1_ASAP7_75t_L g17361 ( 
.A(n_16973),
.Y(n_17361)
);

INVx1_ASAP7_75t_L g17362 ( 
.A(n_17343),
.Y(n_17362)
);

AND2x2_ASAP7_75t_L g17363 ( 
.A(n_16985),
.B(n_16858),
.Y(n_17363)
);

BUFx3_ASAP7_75t_L g17364 ( 
.A(n_16984),
.Y(n_17364)
);

AND2x2_ASAP7_75t_L g17365 ( 
.A(n_16994),
.B(n_16865),
.Y(n_17365)
);

NAND2xp5_ASAP7_75t_L g17366 ( 
.A(n_17266),
.B(n_16878),
.Y(n_17366)
);

INVxp67_ASAP7_75t_L g17367 ( 
.A(n_16970),
.Y(n_17367)
);

AND2x2_ASAP7_75t_L g17368 ( 
.A(n_16980),
.B(n_16907),
.Y(n_17368)
);

NAND2xp5_ASAP7_75t_L g17369 ( 
.A(n_17101),
.B(n_16863),
.Y(n_17369)
);

INVx1_ASAP7_75t_L g17370 ( 
.A(n_17343),
.Y(n_17370)
);

BUFx2_ASAP7_75t_L g17371 ( 
.A(n_17101),
.Y(n_17371)
);

INVx2_ASAP7_75t_L g17372 ( 
.A(n_17343),
.Y(n_17372)
);

NAND2xp5_ASAP7_75t_L g17373 ( 
.A(n_17075),
.B(n_16900),
.Y(n_17373)
);

INVx1_ASAP7_75t_L g17374 ( 
.A(n_17331),
.Y(n_17374)
);

NOR2xp33_ASAP7_75t_L g17375 ( 
.A(n_17032),
.B(n_16742),
.Y(n_17375)
);

AND2x2_ASAP7_75t_L g17376 ( 
.A(n_16981),
.B(n_16704),
.Y(n_17376)
);

NAND2xp5_ASAP7_75t_L g17377 ( 
.A(n_17326),
.B(n_10371),
.Y(n_17377)
);

NOR2xp33_ASAP7_75t_L g17378 ( 
.A(n_16979),
.B(n_10371),
.Y(n_17378)
);

NAND2xp5_ASAP7_75t_SL g17379 ( 
.A(n_17260),
.B(n_10371),
.Y(n_17379)
);

OR2x2_ASAP7_75t_L g17380 ( 
.A(n_17012),
.B(n_10068),
.Y(n_17380)
);

NAND2xp5_ASAP7_75t_L g17381 ( 
.A(n_16988),
.B(n_10068),
.Y(n_17381)
);

INVx1_ASAP7_75t_L g17382 ( 
.A(n_17040),
.Y(n_17382)
);

NOR2x1_ASAP7_75t_L g17383 ( 
.A(n_16996),
.B(n_17007),
.Y(n_17383)
);

AND2x2_ASAP7_75t_L g17384 ( 
.A(n_17066),
.B(n_10092),
.Y(n_17384)
);

AND2x4_ASAP7_75t_L g17385 ( 
.A(n_17112),
.B(n_10151),
.Y(n_17385)
);

BUFx3_ASAP7_75t_L g17386 ( 
.A(n_17193),
.Y(n_17386)
);

HB1xp67_ASAP7_75t_L g17387 ( 
.A(n_17166),
.Y(n_17387)
);

AOI22xp33_ASAP7_75t_L g17388 ( 
.A1(n_17091),
.A2(n_8903),
.B1(n_8536),
.B2(n_8550),
.Y(n_17388)
);

INVx1_ASAP7_75t_SL g17389 ( 
.A(n_17173),
.Y(n_17389)
);

AND2x2_ASAP7_75t_L g17390 ( 
.A(n_17080),
.B(n_10188),
.Y(n_17390)
);

INVx3_ASAP7_75t_L g17391 ( 
.A(n_17016),
.Y(n_17391)
);

OR2x2_ASAP7_75t_L g17392 ( 
.A(n_16971),
.B(n_10079),
.Y(n_17392)
);

INVxp67_ASAP7_75t_L g17393 ( 
.A(n_16987),
.Y(n_17393)
);

NAND2xp5_ASAP7_75t_L g17394 ( 
.A(n_17077),
.B(n_10079),
.Y(n_17394)
);

OAI22xp5_ASAP7_75t_L g17395 ( 
.A1(n_17120),
.A2(n_17053),
.B1(n_17046),
.B2(n_17127),
.Y(n_17395)
);

INVx2_ASAP7_75t_L g17396 ( 
.A(n_17351),
.Y(n_17396)
);

INVx1_ASAP7_75t_SL g17397 ( 
.A(n_17116),
.Y(n_17397)
);

INVx1_ASAP7_75t_SL g17398 ( 
.A(n_17015),
.Y(n_17398)
);

OR2x6_ASAP7_75t_L g17399 ( 
.A(n_17198),
.B(n_7376),
.Y(n_17399)
);

BUFx2_ASAP7_75t_L g17400 ( 
.A(n_17088),
.Y(n_17400)
);

INVx1_ASAP7_75t_L g17401 ( 
.A(n_17130),
.Y(n_17401)
);

OR2x2_ASAP7_75t_L g17402 ( 
.A(n_17017),
.B(n_10080),
.Y(n_17402)
);

INVx1_ASAP7_75t_L g17403 ( 
.A(n_17320),
.Y(n_17403)
);

AND2x2_ASAP7_75t_L g17404 ( 
.A(n_17132),
.B(n_10188),
.Y(n_17404)
);

INVxp67_ASAP7_75t_L g17405 ( 
.A(n_16969),
.Y(n_17405)
);

INVx2_ASAP7_75t_SL g17406 ( 
.A(n_17106),
.Y(n_17406)
);

NAND2xp5_ASAP7_75t_L g17407 ( 
.A(n_17021),
.B(n_10080),
.Y(n_17407)
);

AND2x2_ASAP7_75t_L g17408 ( 
.A(n_17136),
.B(n_10297),
.Y(n_17408)
);

NOR2xp33_ASAP7_75t_L g17409 ( 
.A(n_17002),
.B(n_8038),
.Y(n_17409)
);

INVx2_ASAP7_75t_L g17410 ( 
.A(n_17128),
.Y(n_17410)
);

INVx1_ASAP7_75t_SL g17411 ( 
.A(n_17018),
.Y(n_17411)
);

AND2x2_ASAP7_75t_L g17412 ( 
.A(n_17138),
.B(n_10297),
.Y(n_17412)
);

AND2x2_ASAP7_75t_L g17413 ( 
.A(n_16982),
.B(n_10337),
.Y(n_17413)
);

OR2x2_ASAP7_75t_L g17414 ( 
.A(n_16983),
.B(n_10083),
.Y(n_17414)
);

NOR2xp33_ASAP7_75t_L g17415 ( 
.A(n_16995),
.B(n_8186),
.Y(n_17415)
);

INVx1_ASAP7_75t_SL g17416 ( 
.A(n_17057),
.Y(n_17416)
);

HB1xp67_ASAP7_75t_L g17417 ( 
.A(n_17282),
.Y(n_17417)
);

INVx2_ASAP7_75t_L g17418 ( 
.A(n_17131),
.Y(n_17418)
);

INVx1_ASAP7_75t_SL g17419 ( 
.A(n_17064),
.Y(n_17419)
);

INVx1_ASAP7_75t_L g17420 ( 
.A(n_17246),
.Y(n_17420)
);

AND2x4_ASAP7_75t_L g17421 ( 
.A(n_17010),
.B(n_17013),
.Y(n_17421)
);

AND2x2_ASAP7_75t_L g17422 ( 
.A(n_16992),
.B(n_10337),
.Y(n_17422)
);

NOR2xp33_ASAP7_75t_L g17423 ( 
.A(n_16991),
.B(n_8186),
.Y(n_17423)
);

INVx1_ASAP7_75t_L g17424 ( 
.A(n_17124),
.Y(n_17424)
);

AND2x2_ASAP7_75t_L g17425 ( 
.A(n_17000),
.B(n_10348),
.Y(n_17425)
);

AND2x2_ASAP7_75t_L g17426 ( 
.A(n_17001),
.B(n_10348),
.Y(n_17426)
);

INVx1_ASAP7_75t_L g17427 ( 
.A(n_17310),
.Y(n_17427)
);

INVx1_ASAP7_75t_L g17428 ( 
.A(n_17020),
.Y(n_17428)
);

INVx1_ASAP7_75t_L g17429 ( 
.A(n_16974),
.Y(n_17429)
);

AND2x2_ASAP7_75t_L g17430 ( 
.A(n_17142),
.B(n_8731),
.Y(n_17430)
);

INVx1_ASAP7_75t_L g17431 ( 
.A(n_16978),
.Y(n_17431)
);

AOI22xp33_ASAP7_75t_L g17432 ( 
.A1(n_17006),
.A2(n_8536),
.B1(n_8550),
.B2(n_8437),
.Y(n_17432)
);

INVx1_ASAP7_75t_L g17433 ( 
.A(n_16986),
.Y(n_17433)
);

INVx1_ASAP7_75t_SL g17434 ( 
.A(n_17019),
.Y(n_17434)
);

AOI22xp33_ASAP7_75t_L g17435 ( 
.A1(n_17009),
.A2(n_8550),
.B1(n_8437),
.B2(n_7975),
.Y(n_17435)
);

INVx1_ASAP7_75t_L g17436 ( 
.A(n_17267),
.Y(n_17436)
);

NOR2xp33_ASAP7_75t_L g17437 ( 
.A(n_17005),
.B(n_8186),
.Y(n_17437)
);

INVxp67_ASAP7_75t_L g17438 ( 
.A(n_17050),
.Y(n_17438)
);

AOI22xp33_ASAP7_75t_SL g17439 ( 
.A1(n_17111),
.A2(n_8357),
.B1(n_8390),
.B2(n_8353),
.Y(n_17439)
);

NAND2xp5_ASAP7_75t_L g17440 ( 
.A(n_17014),
.B(n_10083),
.Y(n_17440)
);

HB1xp67_ASAP7_75t_L g17441 ( 
.A(n_17313),
.Y(n_17441)
);

INVx1_ASAP7_75t_L g17442 ( 
.A(n_17268),
.Y(n_17442)
);

AND2x2_ASAP7_75t_L g17443 ( 
.A(n_17011),
.B(n_8731),
.Y(n_17443)
);

AND2x2_ASAP7_75t_L g17444 ( 
.A(n_17145),
.B(n_8755),
.Y(n_17444)
);

NAND2xp5_ASAP7_75t_L g17445 ( 
.A(n_17036),
.B(n_10094),
.Y(n_17445)
);

INVx1_ASAP7_75t_L g17446 ( 
.A(n_17155),
.Y(n_17446)
);

NAND2xp5_ASAP7_75t_L g17447 ( 
.A(n_17076),
.B(n_10094),
.Y(n_17447)
);

CKINVDCx16_ASAP7_75t_R g17448 ( 
.A(n_17340),
.Y(n_17448)
);

CKINVDCx16_ASAP7_75t_R g17449 ( 
.A(n_17292),
.Y(n_17449)
);

CKINVDCx5p33_ASAP7_75t_R g17450 ( 
.A(n_17071),
.Y(n_17450)
);

NAND2xp5_ASAP7_75t_L g17451 ( 
.A(n_16993),
.B(n_17024),
.Y(n_17451)
);

INVxp67_ASAP7_75t_L g17452 ( 
.A(n_17055),
.Y(n_17452)
);

INVx1_ASAP7_75t_L g17453 ( 
.A(n_17097),
.Y(n_17453)
);

INVxp67_ASAP7_75t_L g17454 ( 
.A(n_17105),
.Y(n_17454)
);

INVxp67_ASAP7_75t_SL g17455 ( 
.A(n_17060),
.Y(n_17455)
);

AND2x2_ASAP7_75t_L g17456 ( 
.A(n_17099),
.B(n_17129),
.Y(n_17456)
);

OR2x2_ASAP7_75t_L g17457 ( 
.A(n_17158),
.B(n_17149),
.Y(n_17457)
);

AND3x2_ASAP7_75t_L g17458 ( 
.A(n_17160),
.B(n_17147),
.C(n_17108),
.Y(n_17458)
);

INVxp67_ASAP7_75t_L g17459 ( 
.A(n_17207),
.Y(n_17459)
);

NAND2xp5_ASAP7_75t_L g17460 ( 
.A(n_17200),
.B(n_10109),
.Y(n_17460)
);

AND2x4_ASAP7_75t_L g17461 ( 
.A(n_17123),
.B(n_8755),
.Y(n_17461)
);

INVx1_ASAP7_75t_L g17462 ( 
.A(n_17037),
.Y(n_17462)
);

INVx1_ASAP7_75t_L g17463 ( 
.A(n_17325),
.Y(n_17463)
);

INVx2_ASAP7_75t_L g17464 ( 
.A(n_17336),
.Y(n_17464)
);

OR2x2_ASAP7_75t_L g17465 ( 
.A(n_17270),
.B(n_10109),
.Y(n_17465)
);

AND2x2_ASAP7_75t_L g17466 ( 
.A(n_17231),
.B(n_8755),
.Y(n_17466)
);

INVx1_ASAP7_75t_L g17467 ( 
.A(n_17027),
.Y(n_17467)
);

NOR2xp33_ASAP7_75t_L g17468 ( 
.A(n_17039),
.B(n_8205),
.Y(n_17468)
);

NAND2xp5_ASAP7_75t_L g17469 ( 
.A(n_17082),
.B(n_10111),
.Y(n_17469)
);

INVx1_ASAP7_75t_L g17470 ( 
.A(n_17022),
.Y(n_17470)
);

AND2x2_ASAP7_75t_L g17471 ( 
.A(n_17307),
.B(n_8800),
.Y(n_17471)
);

INVx1_ASAP7_75t_L g17472 ( 
.A(n_17103),
.Y(n_17472)
);

AOI22x1_ASAP7_75t_L g17473 ( 
.A1(n_17043),
.A2(n_6781),
.B1(n_6757),
.B2(n_8357),
.Y(n_17473)
);

INVx2_ASAP7_75t_L g17474 ( 
.A(n_17070),
.Y(n_17474)
);

INVx2_ASAP7_75t_L g17475 ( 
.A(n_17341),
.Y(n_17475)
);

INVx3_ASAP7_75t_L g17476 ( 
.A(n_17030),
.Y(n_17476)
);

INVx1_ASAP7_75t_L g17477 ( 
.A(n_17107),
.Y(n_17477)
);

INVxp33_ASAP7_75t_L g17478 ( 
.A(n_17023),
.Y(n_17478)
);

INVx2_ASAP7_75t_SL g17479 ( 
.A(n_17121),
.Y(n_17479)
);

AND3x1_ASAP7_75t_L g17480 ( 
.A(n_17028),
.B(n_8270),
.C(n_8205),
.Y(n_17480)
);

AND2x4_ASAP7_75t_L g17481 ( 
.A(n_17086),
.B(n_8800),
.Y(n_17481)
);

INVx1_ASAP7_75t_SL g17482 ( 
.A(n_17151),
.Y(n_17482)
);

INVxp67_ASAP7_75t_L g17483 ( 
.A(n_17047),
.Y(n_17483)
);

NOR2x1_ASAP7_75t_L g17484 ( 
.A(n_16972),
.B(n_10111),
.Y(n_17484)
);

INVx1_ASAP7_75t_SL g17485 ( 
.A(n_17074),
.Y(n_17485)
);

AND2x2_ASAP7_75t_L g17486 ( 
.A(n_17146),
.B(n_8800),
.Y(n_17486)
);

AND2x2_ASAP7_75t_L g17487 ( 
.A(n_17125),
.B(n_8810),
.Y(n_17487)
);

OR2x2_ASAP7_75t_L g17488 ( 
.A(n_17073),
.B(n_10113),
.Y(n_17488)
);

NAND2xp5_ASAP7_75t_L g17489 ( 
.A(n_17290),
.B(n_17085),
.Y(n_17489)
);

AND2x2_ASAP7_75t_L g17490 ( 
.A(n_17164),
.B(n_8810),
.Y(n_17490)
);

INVx2_ASAP7_75t_L g17491 ( 
.A(n_17041),
.Y(n_17491)
);

OR2x2_ASAP7_75t_L g17492 ( 
.A(n_17087),
.B(n_10113),
.Y(n_17492)
);

INVx1_ASAP7_75t_L g17493 ( 
.A(n_17067),
.Y(n_17493)
);

INVx1_ASAP7_75t_SL g17494 ( 
.A(n_17295),
.Y(n_17494)
);

OR2x2_ASAP7_75t_L g17495 ( 
.A(n_16989),
.B(n_10116),
.Y(n_17495)
);

INVx1_ASAP7_75t_L g17496 ( 
.A(n_17051),
.Y(n_17496)
);

INVx1_ASAP7_75t_L g17497 ( 
.A(n_17148),
.Y(n_17497)
);

INVx1_ASAP7_75t_SL g17498 ( 
.A(n_17102),
.Y(n_17498)
);

OR2x2_ASAP7_75t_L g17499 ( 
.A(n_16998),
.B(n_10116),
.Y(n_17499)
);

AND2x2_ASAP7_75t_L g17500 ( 
.A(n_17167),
.B(n_8810),
.Y(n_17500)
);

AND2x2_ASAP7_75t_L g17501 ( 
.A(n_17240),
.B(n_8810),
.Y(n_17501)
);

INVx1_ASAP7_75t_SL g17502 ( 
.A(n_17003),
.Y(n_17502)
);

AND2x2_ASAP7_75t_L g17503 ( 
.A(n_17176),
.B(n_8810),
.Y(n_17503)
);

INVxp67_ASAP7_75t_L g17504 ( 
.A(n_17090),
.Y(n_17504)
);

OR2x2_ASAP7_75t_L g17505 ( 
.A(n_17275),
.B(n_10124),
.Y(n_17505)
);

NAND2xp5_ASAP7_75t_L g17506 ( 
.A(n_16990),
.B(n_10124),
.Y(n_17506)
);

INVx1_ASAP7_75t_L g17507 ( 
.A(n_17113),
.Y(n_17507)
);

INVx4_ASAP7_75t_L g17508 ( 
.A(n_17216),
.Y(n_17508)
);

NAND2xp5_ASAP7_75t_L g17509 ( 
.A(n_17243),
.B(n_10128),
.Y(n_17509)
);

NAND2xp5_ASAP7_75t_L g17510 ( 
.A(n_17114),
.B(n_10128),
.Y(n_17510)
);

AND2x2_ASAP7_75t_L g17511 ( 
.A(n_17058),
.B(n_8823),
.Y(n_17511)
);

INVx1_ASAP7_75t_SL g17512 ( 
.A(n_17025),
.Y(n_17512)
);

INVx1_ASAP7_75t_L g17513 ( 
.A(n_17118),
.Y(n_17513)
);

AND2x2_ASAP7_75t_L g17514 ( 
.A(n_17061),
.B(n_8823),
.Y(n_17514)
);

AND2x2_ASAP7_75t_L g17515 ( 
.A(n_17084),
.B(n_8823),
.Y(n_17515)
);

NAND2xp5_ASAP7_75t_L g17516 ( 
.A(n_17122),
.B(n_10134),
.Y(n_17516)
);

NAND2xp5_ASAP7_75t_L g17517 ( 
.A(n_17150),
.B(n_17156),
.Y(n_17517)
);

INVx1_ASAP7_75t_L g17518 ( 
.A(n_17321),
.Y(n_17518)
);

INVx1_ASAP7_75t_L g17519 ( 
.A(n_17184),
.Y(n_17519)
);

AND2x2_ASAP7_75t_L g17520 ( 
.A(n_17049),
.B(n_8823),
.Y(n_17520)
);

OR2x2_ASAP7_75t_L g17521 ( 
.A(n_17301),
.B(n_10134),
.Y(n_17521)
);

NAND2xp5_ASAP7_75t_L g17522 ( 
.A(n_17306),
.B(n_10135),
.Y(n_17522)
);

INVxp67_ASAP7_75t_L g17523 ( 
.A(n_16977),
.Y(n_17523)
);

INVx1_ASAP7_75t_L g17524 ( 
.A(n_17192),
.Y(n_17524)
);

INVx1_ASAP7_75t_L g17525 ( 
.A(n_17199),
.Y(n_17525)
);

NOR2xp33_ASAP7_75t_L g17526 ( 
.A(n_17304),
.B(n_8205),
.Y(n_17526)
);

AOI222xp33_ASAP7_75t_L g17527 ( 
.A1(n_17348),
.A2(n_9317),
.B1(n_9305),
.B2(n_9651),
.C1(n_9653),
.C2(n_9419),
.Y(n_17527)
);

HB1xp67_ASAP7_75t_L g17528 ( 
.A(n_17098),
.Y(n_17528)
);

INVx1_ASAP7_75t_L g17529 ( 
.A(n_17210),
.Y(n_17529)
);

INVx1_ASAP7_75t_SL g17530 ( 
.A(n_17253),
.Y(n_17530)
);

AND2x2_ASAP7_75t_L g17531 ( 
.A(n_17276),
.B(n_8823),
.Y(n_17531)
);

OR2x2_ASAP7_75t_L g17532 ( 
.A(n_17241),
.B(n_10135),
.Y(n_17532)
);

NAND2xp5_ASAP7_75t_SL g17533 ( 
.A(n_17026),
.B(n_8205),
.Y(n_17533)
);

OR2x2_ASAP7_75t_L g17534 ( 
.A(n_17255),
.B(n_10138),
.Y(n_17534)
);

OAI21x1_ASAP7_75t_L g17535 ( 
.A1(n_17159),
.A2(n_9905),
.B(n_9317),
.Y(n_17535)
);

AND2x4_ASAP7_75t_L g17536 ( 
.A(n_17154),
.B(n_8835),
.Y(n_17536)
);

INVx2_ASAP7_75t_L g17537 ( 
.A(n_17181),
.Y(n_17537)
);

NOR2xp33_ASAP7_75t_L g17538 ( 
.A(n_17335),
.B(n_8205),
.Y(n_17538)
);

NAND2xp5_ASAP7_75t_L g17539 ( 
.A(n_17356),
.B(n_10138),
.Y(n_17539)
);

INVx2_ASAP7_75t_L g17540 ( 
.A(n_17183),
.Y(n_17540)
);

INVx1_ASAP7_75t_SL g17541 ( 
.A(n_17179),
.Y(n_17541)
);

INVx2_ASAP7_75t_L g17542 ( 
.A(n_17305),
.Y(n_17542)
);

AOI22xp5_ASAP7_75t_L g17543 ( 
.A1(n_17069),
.A2(n_8403),
.B1(n_8408),
.B2(n_8390),
.Y(n_17543)
);

INVx2_ASAP7_75t_L g17544 ( 
.A(n_17203),
.Y(n_17544)
);

NAND2xp5_ASAP7_75t_L g17545 ( 
.A(n_17323),
.B(n_17265),
.Y(n_17545)
);

AND3x1_ASAP7_75t_L g17546 ( 
.A(n_17004),
.B(n_8288),
.C(n_8270),
.Y(n_17546)
);

AND2x2_ASAP7_75t_L g17547 ( 
.A(n_17062),
.B(n_17299),
.Y(n_17547)
);

INVx2_ASAP7_75t_L g17548 ( 
.A(n_17189),
.Y(n_17548)
);

INVx1_ASAP7_75t_SL g17549 ( 
.A(n_17029),
.Y(n_17549)
);

AND2x2_ASAP7_75t_L g17550 ( 
.A(n_17322),
.B(n_8835),
.Y(n_17550)
);

HB1xp67_ASAP7_75t_L g17551 ( 
.A(n_17165),
.Y(n_17551)
);

AND2x2_ASAP7_75t_L g17552 ( 
.A(n_17308),
.B(n_8835),
.Y(n_17552)
);

INVx1_ASAP7_75t_L g17553 ( 
.A(n_17048),
.Y(n_17553)
);

INVx2_ASAP7_75t_L g17554 ( 
.A(n_17355),
.Y(n_17554)
);

AND2x2_ASAP7_75t_L g17555 ( 
.A(n_17033),
.B(n_8835),
.Y(n_17555)
);

NAND2xp5_ASAP7_75t_L g17556 ( 
.A(n_17354),
.B(n_10143),
.Y(n_17556)
);

AOI22xp5_ASAP7_75t_L g17557 ( 
.A1(n_17293),
.A2(n_8403),
.B1(n_8408),
.B2(n_8390),
.Y(n_17557)
);

INVx1_ASAP7_75t_L g17558 ( 
.A(n_17137),
.Y(n_17558)
);

OR2x2_ASAP7_75t_L g17559 ( 
.A(n_17169),
.B(n_10143),
.Y(n_17559)
);

NAND2xp5_ASAP7_75t_L g17560 ( 
.A(n_17153),
.B(n_10144),
.Y(n_17560)
);

INVx1_ASAP7_75t_L g17561 ( 
.A(n_17140),
.Y(n_17561)
);

INVx4_ASAP7_75t_L g17562 ( 
.A(n_17297),
.Y(n_17562)
);

INVx1_ASAP7_75t_L g17563 ( 
.A(n_17065),
.Y(n_17563)
);

INVx4_ASAP7_75t_L g17564 ( 
.A(n_17162),
.Y(n_17564)
);

AND2x2_ASAP7_75t_L g17565 ( 
.A(n_17143),
.B(n_17170),
.Y(n_17565)
);

BUFx3_ASAP7_75t_L g17566 ( 
.A(n_17045),
.Y(n_17566)
);

AOI22x1_ASAP7_75t_L g17567 ( 
.A1(n_17349),
.A2(n_17346),
.B1(n_17333),
.B2(n_17298),
.Y(n_17567)
);

AND2x4_ASAP7_75t_L g17568 ( 
.A(n_17337),
.B(n_8835),
.Y(n_17568)
);

AND2x2_ASAP7_75t_L g17569 ( 
.A(n_17190),
.B(n_8950),
.Y(n_17569)
);

INVx2_ASAP7_75t_L g17570 ( 
.A(n_17332),
.Y(n_17570)
);

NAND2xp5_ASAP7_75t_L g17571 ( 
.A(n_17052),
.B(n_10144),
.Y(n_17571)
);

AND2x2_ASAP7_75t_L g17572 ( 
.A(n_17194),
.B(n_8950),
.Y(n_17572)
);

OR2x2_ASAP7_75t_L g17573 ( 
.A(n_17300),
.B(n_10147),
.Y(n_17573)
);

AND2x2_ASAP7_75t_L g17574 ( 
.A(n_17056),
.B(n_8950),
.Y(n_17574)
);

NOR2x1p5_ASAP7_75t_SL g17575 ( 
.A(n_17094),
.B(n_10147),
.Y(n_17575)
);

INVx1_ASAP7_75t_L g17576 ( 
.A(n_17117),
.Y(n_17576)
);

INVx1_ASAP7_75t_L g17577 ( 
.A(n_17119),
.Y(n_17577)
);

AND2x2_ASAP7_75t_L g17578 ( 
.A(n_17059),
.B(n_8950),
.Y(n_17578)
);

INVx2_ASAP7_75t_L g17579 ( 
.A(n_17339),
.Y(n_17579)
);

AND2x4_ASAP7_75t_L g17580 ( 
.A(n_17187),
.B(n_8950),
.Y(n_17580)
);

INVx1_ASAP7_75t_SL g17581 ( 
.A(n_17063),
.Y(n_17581)
);

NAND2xp5_ASAP7_75t_L g17582 ( 
.A(n_17038),
.B(n_10152),
.Y(n_17582)
);

AOI22xp5_ASAP7_75t_L g17583 ( 
.A1(n_17100),
.A2(n_8408),
.B1(n_8434),
.B2(n_8403),
.Y(n_17583)
);

INVxp67_ASAP7_75t_L g17584 ( 
.A(n_17068),
.Y(n_17584)
);

NAND2xp5_ASAP7_75t_L g17585 ( 
.A(n_17135),
.B(n_17141),
.Y(n_17585)
);

INVxp67_ASAP7_75t_L g17586 ( 
.A(n_17083),
.Y(n_17586)
);

AND2x2_ASAP7_75t_L g17587 ( 
.A(n_17186),
.B(n_8978),
.Y(n_17587)
);

OR2x2_ASAP7_75t_L g17588 ( 
.A(n_17229),
.B(n_10152),
.Y(n_17588)
);

INVx1_ASAP7_75t_L g17589 ( 
.A(n_17172),
.Y(n_17589)
);

INVx1_ASAP7_75t_SL g17590 ( 
.A(n_17144),
.Y(n_17590)
);

INVx2_ASAP7_75t_L g17591 ( 
.A(n_17329),
.Y(n_17591)
);

OR2x2_ASAP7_75t_L g17592 ( 
.A(n_17233),
.B(n_10155),
.Y(n_17592)
);

INVx1_ASAP7_75t_SL g17593 ( 
.A(n_17152),
.Y(n_17593)
);

BUFx3_ASAP7_75t_L g17594 ( 
.A(n_17296),
.Y(n_17594)
);

AND2x2_ASAP7_75t_L g17595 ( 
.A(n_17182),
.B(n_8978),
.Y(n_17595)
);

NAND2xp33_ASAP7_75t_L g17596 ( 
.A(n_17212),
.B(n_10155),
.Y(n_17596)
);

OAI21x1_ASAP7_75t_L g17597 ( 
.A1(n_17227),
.A2(n_9317),
.B(n_9305),
.Y(n_17597)
);

OAI21x1_ASAP7_75t_L g17598 ( 
.A1(n_17034),
.A2(n_9305),
.B(n_10248),
.Y(n_17598)
);

INVx2_ASAP7_75t_L g17599 ( 
.A(n_17256),
.Y(n_17599)
);

NAND2xp5_ASAP7_75t_L g17600 ( 
.A(n_17174),
.B(n_10161),
.Y(n_17600)
);

INVx1_ASAP7_75t_L g17601 ( 
.A(n_17054),
.Y(n_17601)
);

INVx1_ASAP7_75t_SL g17602 ( 
.A(n_17079),
.Y(n_17602)
);

INVx1_ASAP7_75t_L g17603 ( 
.A(n_17161),
.Y(n_17603)
);

INVx1_ASAP7_75t_L g17604 ( 
.A(n_17031),
.Y(n_17604)
);

INVx1_ASAP7_75t_L g17605 ( 
.A(n_17035),
.Y(n_17605)
);

INVx1_ASAP7_75t_L g17606 ( 
.A(n_17089),
.Y(n_17606)
);

NOR3xp33_ASAP7_75t_L g17607 ( 
.A(n_17206),
.B(n_8288),
.C(n_8270),
.Y(n_17607)
);

INVx1_ASAP7_75t_L g17608 ( 
.A(n_17093),
.Y(n_17608)
);

INVx2_ASAP7_75t_SL g17609 ( 
.A(n_17201),
.Y(n_17609)
);

BUFx2_ASAP7_75t_L g17610 ( 
.A(n_17175),
.Y(n_17610)
);

AO21x2_ASAP7_75t_L g17611 ( 
.A1(n_17220),
.A2(n_10164),
.B(n_10161),
.Y(n_17611)
);

NOR2xp33_ASAP7_75t_L g17612 ( 
.A(n_16999),
.B(n_8270),
.Y(n_17612)
);

INVxp67_ASAP7_75t_L g17613 ( 
.A(n_17134),
.Y(n_17613)
);

AND2x2_ASAP7_75t_L g17614 ( 
.A(n_17163),
.B(n_17273),
.Y(n_17614)
);

INVx1_ASAP7_75t_L g17615 ( 
.A(n_17133),
.Y(n_17615)
);

NAND2xp5_ASAP7_75t_L g17616 ( 
.A(n_17213),
.B(n_10164),
.Y(n_17616)
);

INVx1_ASAP7_75t_L g17617 ( 
.A(n_17139),
.Y(n_17617)
);

NAND2xp5_ASAP7_75t_L g17618 ( 
.A(n_17218),
.B(n_10172),
.Y(n_17618)
);

INVx1_ASAP7_75t_SL g17619 ( 
.A(n_17221),
.Y(n_17619)
);

INVx3_ASAP7_75t_L g17620 ( 
.A(n_17274),
.Y(n_17620)
);

INVx1_ASAP7_75t_L g17621 ( 
.A(n_17284),
.Y(n_17621)
);

NOR2x1_ASAP7_75t_L g17622 ( 
.A(n_17224),
.B(n_10172),
.Y(n_17622)
);

INVx1_ASAP7_75t_L g17623 ( 
.A(n_17204),
.Y(n_17623)
);

INVx1_ASAP7_75t_L g17624 ( 
.A(n_17214),
.Y(n_17624)
);

AOI22xp33_ASAP7_75t_L g17625 ( 
.A1(n_17171),
.A2(n_8550),
.B1(n_8437),
.B2(n_7975),
.Y(n_17625)
);

NAND2xp5_ASAP7_75t_L g17626 ( 
.A(n_17237),
.B(n_10179),
.Y(n_17626)
);

NAND2xp5_ASAP7_75t_L g17627 ( 
.A(n_16997),
.B(n_10179),
.Y(n_17627)
);

INVx2_ASAP7_75t_SL g17628 ( 
.A(n_17196),
.Y(n_17628)
);

OAI22xp5_ASAP7_75t_L g17629 ( 
.A1(n_17291),
.A2(n_10185),
.B1(n_10193),
.B2(n_10182),
.Y(n_17629)
);

OA21x2_ASAP7_75t_L g17630 ( 
.A1(n_17168),
.A2(n_10321),
.B(n_10248),
.Y(n_17630)
);

INVx1_ASAP7_75t_L g17631 ( 
.A(n_17225),
.Y(n_17631)
);

AND2x2_ASAP7_75t_L g17632 ( 
.A(n_17280),
.B(n_17281),
.Y(n_17632)
);

OR2x2_ASAP7_75t_L g17633 ( 
.A(n_17314),
.B(n_10182),
.Y(n_17633)
);

CKINVDCx16_ASAP7_75t_R g17634 ( 
.A(n_17205),
.Y(n_17634)
);

AND2x2_ASAP7_75t_L g17635 ( 
.A(n_17287),
.B(n_8978),
.Y(n_17635)
);

INVx1_ASAP7_75t_SL g17636 ( 
.A(n_17245),
.Y(n_17636)
);

INVx4_ASAP7_75t_L g17637 ( 
.A(n_17262),
.Y(n_17637)
);

INVx1_ASAP7_75t_L g17638 ( 
.A(n_17234),
.Y(n_17638)
);

AND2x2_ASAP7_75t_L g17639 ( 
.A(n_17248),
.B(n_8978),
.Y(n_17639)
);

AND2x2_ASAP7_75t_L g17640 ( 
.A(n_17236),
.B(n_8978),
.Y(n_17640)
);

AND2x4_ASAP7_75t_L g17641 ( 
.A(n_17211),
.B(n_9018),
.Y(n_17641)
);

BUFx2_ASAP7_75t_L g17642 ( 
.A(n_17238),
.Y(n_17642)
);

AND2x2_ASAP7_75t_L g17643 ( 
.A(n_17217),
.B(n_9018),
.Y(n_17643)
);

INVx4_ASAP7_75t_L g17644 ( 
.A(n_17264),
.Y(n_17644)
);

NAND2xp5_ASAP7_75t_L g17645 ( 
.A(n_17252),
.B(n_10185),
.Y(n_17645)
);

AND2x2_ASAP7_75t_L g17646 ( 
.A(n_17244),
.B(n_9018),
.Y(n_17646)
);

INVx1_ASAP7_75t_L g17647 ( 
.A(n_17239),
.Y(n_17647)
);

AOI22xp33_ASAP7_75t_L g17648 ( 
.A1(n_17350),
.A2(n_8437),
.B1(n_7975),
.B2(n_8434),
.Y(n_17648)
);

OAI22xp5_ASAP7_75t_L g17649 ( 
.A1(n_17259),
.A2(n_10195),
.B1(n_10199),
.B2(n_10193),
.Y(n_17649)
);

AND2x2_ASAP7_75t_L g17650 ( 
.A(n_17249),
.B(n_9018),
.Y(n_17650)
);

INVx1_ASAP7_75t_L g17651 ( 
.A(n_17242),
.Y(n_17651)
);

INVx2_ASAP7_75t_L g17652 ( 
.A(n_17247),
.Y(n_17652)
);

INVx1_ASAP7_75t_L g17653 ( 
.A(n_17208),
.Y(n_17653)
);

AND2x4_ASAP7_75t_L g17654 ( 
.A(n_17312),
.B(n_9018),
.Y(n_17654)
);

INVx1_ASAP7_75t_L g17655 ( 
.A(n_17180),
.Y(n_17655)
);

AND2x2_ASAP7_75t_L g17656 ( 
.A(n_17228),
.B(n_9027),
.Y(n_17656)
);

INVx1_ASAP7_75t_L g17657 ( 
.A(n_17191),
.Y(n_17657)
);

AND2x2_ASAP7_75t_L g17658 ( 
.A(n_17104),
.B(n_17197),
.Y(n_17658)
);

CKINVDCx16_ASAP7_75t_R g17659 ( 
.A(n_17286),
.Y(n_17659)
);

NAND2xp5_ASAP7_75t_L g17660 ( 
.A(n_17261),
.B(n_17303),
.Y(n_17660)
);

INVx1_ASAP7_75t_L g17661 ( 
.A(n_17288),
.Y(n_17661)
);

OR2x2_ASAP7_75t_L g17662 ( 
.A(n_17178),
.B(n_10195),
.Y(n_17662)
);

NOR2xp33_ASAP7_75t_L g17663 ( 
.A(n_17352),
.B(n_8270),
.Y(n_17663)
);

HB1xp67_ASAP7_75t_L g17664 ( 
.A(n_17258),
.Y(n_17664)
);

INVxp67_ASAP7_75t_L g17665 ( 
.A(n_17257),
.Y(n_17665)
);

OR2x2_ASAP7_75t_L g17666 ( 
.A(n_17185),
.B(n_10199),
.Y(n_17666)
);

AND2x2_ASAP7_75t_L g17667 ( 
.A(n_17223),
.B(n_9027),
.Y(n_17667)
);

OR2x2_ASAP7_75t_L g17668 ( 
.A(n_17277),
.B(n_10203),
.Y(n_17668)
);

AND2x2_ASAP7_75t_L g17669 ( 
.A(n_17235),
.B(n_9027),
.Y(n_17669)
);

AND2x2_ASAP7_75t_L g17670 ( 
.A(n_17110),
.B(n_9027),
.Y(n_17670)
);

INVx1_ASAP7_75t_L g17671 ( 
.A(n_17294),
.Y(n_17671)
);

INVx1_ASAP7_75t_L g17672 ( 
.A(n_17334),
.Y(n_17672)
);

HB1xp67_ASAP7_75t_L g17673 ( 
.A(n_17338),
.Y(n_17673)
);

INVx2_ASAP7_75t_L g17674 ( 
.A(n_17250),
.Y(n_17674)
);

INVx1_ASAP7_75t_L g17675 ( 
.A(n_17317),
.Y(n_17675)
);

INVx1_ASAP7_75t_L g17676 ( 
.A(n_17311),
.Y(n_17676)
);

AND2x2_ASAP7_75t_L g17677 ( 
.A(n_17289),
.B(n_9027),
.Y(n_17677)
);

INVx1_ASAP7_75t_L g17678 ( 
.A(n_17177),
.Y(n_17678)
);

NOR3xp33_ASAP7_75t_L g17679 ( 
.A(n_17448),
.B(n_17342),
.C(n_17044),
.Y(n_17679)
);

INVx2_ASAP7_75t_L g17680 ( 
.A(n_17371),
.Y(n_17680)
);

OAI21xp5_ASAP7_75t_L g17681 ( 
.A1(n_17393),
.A2(n_17188),
.B(n_17109),
.Y(n_17681)
);

NAND2xp5_ASAP7_75t_L g17682 ( 
.A(n_17449),
.B(n_17092),
.Y(n_17682)
);

INVx2_ASAP7_75t_L g17683 ( 
.A(n_17372),
.Y(n_17683)
);

OAI22xp5_ASAP7_75t_L g17684 ( 
.A1(n_17367),
.A2(n_17263),
.B1(n_17251),
.B2(n_17327),
.Y(n_17684)
);

NAND2xp5_ASAP7_75t_L g17685 ( 
.A(n_17421),
.B(n_17279),
.Y(n_17685)
);

AOI22xp5_ASAP7_75t_L g17686 ( 
.A1(n_17357),
.A2(n_17081),
.B1(n_17072),
.B2(n_17344),
.Y(n_17686)
);

AOI221x1_ASAP7_75t_L g17687 ( 
.A1(n_17395),
.A2(n_17361),
.B1(n_17374),
.B2(n_17463),
.C(n_17382),
.Y(n_17687)
);

INVx1_ASAP7_75t_L g17688 ( 
.A(n_17362),
.Y(n_17688)
);

OAI221xp5_ASAP7_75t_L g17689 ( 
.A1(n_17523),
.A2(n_17269),
.B1(n_17309),
.B2(n_17316),
.C(n_17353),
.Y(n_17689)
);

OR2x2_ASAP7_75t_L g17690 ( 
.A(n_17389),
.B(n_17278),
.Y(n_17690)
);

BUFx2_ASAP7_75t_L g17691 ( 
.A(n_17383),
.Y(n_17691)
);

NAND2xp5_ASAP7_75t_L g17692 ( 
.A(n_17458),
.B(n_17391),
.Y(n_17692)
);

AOI221xp5_ASAP7_75t_L g17693 ( 
.A1(n_17480),
.A2(n_17347),
.B1(n_17226),
.B2(n_17324),
.C(n_17319),
.Y(n_17693)
);

INVx1_ASAP7_75t_L g17694 ( 
.A(n_17370),
.Y(n_17694)
);

NOR2xp67_ASAP7_75t_L g17695 ( 
.A(n_17387),
.B(n_17347),
.Y(n_17695)
);

INVx1_ASAP7_75t_L g17696 ( 
.A(n_17441),
.Y(n_17696)
);

NAND2x1_ASAP7_75t_L g17697 ( 
.A(n_17396),
.B(n_17254),
.Y(n_17697)
);

NAND2xp5_ASAP7_75t_L g17698 ( 
.A(n_17411),
.B(n_17318),
.Y(n_17698)
);

INVx1_ASAP7_75t_SL g17699 ( 
.A(n_17494),
.Y(n_17699)
);

INVx1_ASAP7_75t_L g17700 ( 
.A(n_17528),
.Y(n_17700)
);

NAND2xp5_ASAP7_75t_L g17701 ( 
.A(n_17428),
.B(n_17302),
.Y(n_17701)
);

NAND2xp5_ASAP7_75t_L g17702 ( 
.A(n_17398),
.B(n_17345),
.Y(n_17702)
);

AOI221xp5_ASAP7_75t_L g17703 ( 
.A1(n_17546),
.A2(n_17405),
.B1(n_17478),
.B2(n_17530),
.C(n_17452),
.Y(n_17703)
);

NAND2xp5_ASAP7_75t_L g17704 ( 
.A(n_17416),
.B(n_17328),
.Y(n_17704)
);

OAI32xp33_ASAP7_75t_L g17705 ( 
.A1(n_17502),
.A2(n_17042),
.A3(n_17202),
.B1(n_17157),
.B2(n_17115),
.Y(n_17705)
);

INVx1_ASAP7_75t_SL g17706 ( 
.A(n_17397),
.Y(n_17706)
);

INVx1_ASAP7_75t_L g17707 ( 
.A(n_17551),
.Y(n_17707)
);

INVx2_ASAP7_75t_L g17708 ( 
.A(n_17360),
.Y(n_17708)
);

INVx1_ASAP7_75t_L g17709 ( 
.A(n_17575),
.Y(n_17709)
);

INVxp67_ASAP7_75t_L g17710 ( 
.A(n_17417),
.Y(n_17710)
);

OAI22xp5_ASAP7_75t_L g17711 ( 
.A1(n_17438),
.A2(n_17096),
.B1(n_17209),
.B2(n_17330),
.Y(n_17711)
);

INVx1_ASAP7_75t_SL g17712 ( 
.A(n_17386),
.Y(n_17712)
);

AND2x2_ASAP7_75t_L g17713 ( 
.A(n_17475),
.B(n_17272),
.Y(n_17713)
);

INVx2_ASAP7_75t_L g17714 ( 
.A(n_17364),
.Y(n_17714)
);

OAI22xp5_ASAP7_75t_L g17715 ( 
.A1(n_17454),
.A2(n_17315),
.B1(n_17271),
.B2(n_17095),
.Y(n_17715)
);

HB1xp67_ASAP7_75t_L g17716 ( 
.A(n_17399),
.Y(n_17716)
);

INVx1_ASAP7_75t_L g17717 ( 
.A(n_17455),
.Y(n_17717)
);

OAI22xp5_ASAP7_75t_L g17718 ( 
.A1(n_17419),
.A2(n_17215),
.B1(n_17285),
.B2(n_17078),
.Y(n_17718)
);

AOI21xp5_ASAP7_75t_L g17719 ( 
.A1(n_17489),
.A2(n_17222),
.B(n_17283),
.Y(n_17719)
);

INVx1_ASAP7_75t_L g17720 ( 
.A(n_17658),
.Y(n_17720)
);

INVx2_ASAP7_75t_L g17721 ( 
.A(n_17566),
.Y(n_17721)
);

O2A1O1Ixp33_ASAP7_75t_L g17722 ( 
.A1(n_17420),
.A2(n_17232),
.B(n_17230),
.C(n_17219),
.Y(n_17722)
);

AOI22xp33_ASAP7_75t_L g17723 ( 
.A1(n_17562),
.A2(n_17508),
.B1(n_17594),
.B2(n_17453),
.Y(n_17723)
);

INVx1_ASAP7_75t_L g17724 ( 
.A(n_17565),
.Y(n_17724)
);

AOI222xp33_ASAP7_75t_L g17725 ( 
.A1(n_17434),
.A2(n_17195),
.B1(n_17126),
.B2(n_10208),
.C1(n_10217),
.C2(n_10236),
.Y(n_17725)
);

AOI22xp33_ASAP7_75t_L g17726 ( 
.A1(n_17476),
.A2(n_8434),
.B1(n_8558),
.B2(n_8496),
.Y(n_17726)
);

NAND2xp5_ASAP7_75t_L g17727 ( 
.A(n_17436),
.B(n_17442),
.Y(n_17727)
);

NAND2xp5_ASAP7_75t_L g17728 ( 
.A(n_17481),
.B(n_10203),
.Y(n_17728)
);

OAI21xp33_ASAP7_75t_L g17729 ( 
.A1(n_17471),
.A2(n_8331),
.B(n_8288),
.Y(n_17729)
);

AOI322xp5_ASAP7_75t_L g17730 ( 
.A1(n_17512),
.A2(n_8288),
.A3(n_8331),
.B1(n_8384),
.B2(n_8423),
.C1(n_8421),
.C2(n_8371),
.Y(n_17730)
);

INVx1_ASAP7_75t_L g17731 ( 
.A(n_17457),
.Y(n_17731)
);

XOR2xp5_ASAP7_75t_L g17732 ( 
.A(n_17450),
.B(n_8293),
.Y(n_17732)
);

INVx1_ASAP7_75t_L g17733 ( 
.A(n_17591),
.Y(n_17733)
);

NOR3xp33_ASAP7_75t_L g17734 ( 
.A(n_17634),
.B(n_8331),
.C(n_8288),
.Y(n_17734)
);

OAI32xp33_ASAP7_75t_L g17735 ( 
.A1(n_17545),
.A2(n_8384),
.A3(n_8421),
.B1(n_8371),
.B2(n_8331),
.Y(n_17735)
);

AOI22xp5_ASAP7_75t_L g17736 ( 
.A1(n_17550),
.A2(n_8371),
.B1(n_8384),
.B2(n_8331),
.Y(n_17736)
);

INVx1_ASAP7_75t_SL g17737 ( 
.A(n_17456),
.Y(n_17737)
);

A2O1A1Ixp33_ASAP7_75t_L g17738 ( 
.A1(n_17375),
.A2(n_10321),
.B(n_10248),
.C(n_10217),
.Y(n_17738)
);

NAND2xp5_ASAP7_75t_L g17739 ( 
.A(n_17403),
.B(n_10208),
.Y(n_17739)
);

INVx1_ASAP7_75t_L g17740 ( 
.A(n_17610),
.Y(n_17740)
);

AOI21xp5_ASAP7_75t_L g17741 ( 
.A1(n_17660),
.A2(n_10236),
.B(n_10231),
.Y(n_17741)
);

OAI21x1_ASAP7_75t_SL g17742 ( 
.A1(n_17474),
.A2(n_8558),
.B(n_8496),
.Y(n_17742)
);

AOI32xp33_ASAP7_75t_L g17743 ( 
.A1(n_17612),
.A2(n_8421),
.A3(n_8423),
.B1(n_8384),
.B2(n_8371),
.Y(n_17743)
);

OAI21xp5_ASAP7_75t_L g17744 ( 
.A1(n_17459),
.A2(n_7734),
.B(n_7733),
.Y(n_17744)
);

INVx1_ASAP7_75t_L g17745 ( 
.A(n_17443),
.Y(n_17745)
);

INVx1_ASAP7_75t_L g17746 ( 
.A(n_17400),
.Y(n_17746)
);

AND2x2_ASAP7_75t_L g17747 ( 
.A(n_17486),
.B(n_10231),
.Y(n_17747)
);

AOI222xp33_ASAP7_75t_L g17748 ( 
.A1(n_17498),
.A2(n_17401),
.B1(n_17482),
.B2(n_17533),
.C1(n_17427),
.C2(n_17359),
.Y(n_17748)
);

INVxp67_ASAP7_75t_L g17749 ( 
.A(n_17468),
.Y(n_17749)
);

AOI211xp5_ASAP7_75t_L g17750 ( 
.A1(n_17526),
.A2(n_6757),
.B(n_6781),
.C(n_7198),
.Y(n_17750)
);

AOI22xp5_ASAP7_75t_L g17751 ( 
.A1(n_17466),
.A2(n_8371),
.B1(n_8421),
.B2(n_8384),
.Y(n_17751)
);

O2A1O1Ixp33_ASAP7_75t_SL g17752 ( 
.A1(n_17379),
.A2(n_8558),
.B(n_8676),
.C(n_8496),
.Y(n_17752)
);

OAI21xp5_ASAP7_75t_L g17753 ( 
.A1(n_17409),
.A2(n_17373),
.B(n_17519),
.Y(n_17753)
);

OR2x2_ASAP7_75t_L g17754 ( 
.A(n_17659),
.B(n_10256),
.Y(n_17754)
);

OR2x2_ASAP7_75t_L g17755 ( 
.A(n_17609),
.B(n_10256),
.Y(n_17755)
);

NOR2xp33_ASAP7_75t_L g17756 ( 
.A(n_17564),
.B(n_8421),
.Y(n_17756)
);

INVx1_ASAP7_75t_L g17757 ( 
.A(n_17446),
.Y(n_17757)
);

OAI221xp5_ASAP7_75t_L g17758 ( 
.A1(n_17567),
.A2(n_6781),
.B1(n_8726),
.B2(n_8913),
.C(n_8676),
.Y(n_17758)
);

AND2x2_ASAP7_75t_L g17759 ( 
.A(n_17430),
.B(n_10257),
.Y(n_17759)
);

NOR2xp67_ASAP7_75t_L g17760 ( 
.A(n_17620),
.B(n_10257),
.Y(n_17760)
);

AND2x2_ASAP7_75t_L g17761 ( 
.A(n_17568),
.B(n_10259),
.Y(n_17761)
);

NOR2xp33_ASAP7_75t_L g17762 ( 
.A(n_17541),
.B(n_8423),
.Y(n_17762)
);

AND2x2_ASAP7_75t_L g17763 ( 
.A(n_17547),
.B(n_10259),
.Y(n_17763)
);

O2A1O1Ixp33_ASAP7_75t_L g17764 ( 
.A1(n_17369),
.A2(n_17525),
.B(n_17529),
.C(n_17524),
.Y(n_17764)
);

INVx1_ASAP7_75t_L g17765 ( 
.A(n_17462),
.Y(n_17765)
);

A2O1A1Ixp33_ASAP7_75t_L g17766 ( 
.A1(n_17538),
.A2(n_10321),
.B(n_10261),
.C(n_10270),
.Y(n_17766)
);

INVx1_ASAP7_75t_L g17767 ( 
.A(n_17365),
.Y(n_17767)
);

INVx1_ASAP7_75t_L g17768 ( 
.A(n_17429),
.Y(n_17768)
);

INVx2_ASAP7_75t_L g17769 ( 
.A(n_17552),
.Y(n_17769)
);

INVx1_ASAP7_75t_L g17770 ( 
.A(n_17431),
.Y(n_17770)
);

NAND3xp33_ASAP7_75t_L g17771 ( 
.A(n_17433),
.B(n_10150),
.C(n_10104),
.Y(n_17771)
);

INVx1_ASAP7_75t_L g17772 ( 
.A(n_17410),
.Y(n_17772)
);

OAI33xp33_ASAP7_75t_L g17773 ( 
.A1(n_17366),
.A2(n_10270),
.A3(n_10260),
.B1(n_10275),
.B2(n_10274),
.B3(n_10261),
.Y(n_17773)
);

AOI22xp33_ASAP7_75t_L g17774 ( 
.A1(n_17520),
.A2(n_8726),
.B1(n_8913),
.B2(n_8676),
.Y(n_17774)
);

NAND2xp5_ASAP7_75t_L g17775 ( 
.A(n_17461),
.B(n_10260),
.Y(n_17775)
);

AND2x2_ASAP7_75t_L g17776 ( 
.A(n_17444),
.B(n_17399),
.Y(n_17776)
);

INVx2_ASAP7_75t_L g17777 ( 
.A(n_17531),
.Y(n_17777)
);

AO32x1_ASAP7_75t_L g17778 ( 
.A1(n_17628),
.A2(n_8963),
.A3(n_8913),
.B1(n_8726),
.B2(n_10274),
.Y(n_17778)
);

AOI21xp33_ASAP7_75t_L g17779 ( 
.A1(n_17485),
.A2(n_10150),
.B(n_10104),
.Y(n_17779)
);

INVx1_ASAP7_75t_L g17780 ( 
.A(n_17418),
.Y(n_17780)
);

AND2x2_ASAP7_75t_L g17781 ( 
.A(n_17490),
.B(n_10275),
.Y(n_17781)
);

INVx1_ASAP7_75t_L g17782 ( 
.A(n_17451),
.Y(n_17782)
);

AND2x2_ASAP7_75t_L g17783 ( 
.A(n_17500),
.B(n_10276),
.Y(n_17783)
);

NAND2xp5_ASAP7_75t_L g17784 ( 
.A(n_17590),
.B(n_10276),
.Y(n_17784)
);

HB1xp67_ASAP7_75t_L g17785 ( 
.A(n_17491),
.Y(n_17785)
);

OAI33xp33_ASAP7_75t_L g17786 ( 
.A1(n_17539),
.A2(n_10293),
.A3(n_10281),
.B1(n_10300),
.B2(n_10296),
.B3(n_10285),
.Y(n_17786)
);

XOR2xp5_ASAP7_75t_L g17787 ( 
.A(n_17470),
.B(n_8293),
.Y(n_17787)
);

AOI31xp33_ASAP7_75t_L g17788 ( 
.A1(n_17549),
.A2(n_8569),
.A3(n_8585),
.B(n_8366),
.Y(n_17788)
);

INVxp67_ASAP7_75t_SL g17789 ( 
.A(n_17585),
.Y(n_17789)
);

AOI21xp33_ASAP7_75t_SL g17790 ( 
.A1(n_17493),
.A2(n_8437),
.B(n_8369),
.Y(n_17790)
);

OR2x2_ASAP7_75t_L g17791 ( 
.A(n_17593),
.B(n_10281),
.Y(n_17791)
);

INVx1_ASAP7_75t_L g17792 ( 
.A(n_17487),
.Y(n_17792)
);

INVxp67_ASAP7_75t_L g17793 ( 
.A(n_17358),
.Y(n_17793)
);

AND2x4_ASAP7_75t_L g17794 ( 
.A(n_17652),
.B(n_10285),
.Y(n_17794)
);

OR2x2_ASAP7_75t_L g17795 ( 
.A(n_17619),
.B(n_10293),
.Y(n_17795)
);

NAND2xp5_ASAP7_75t_L g17796 ( 
.A(n_17581),
.B(n_10296),
.Y(n_17796)
);

NAND2xp5_ASAP7_75t_L g17797 ( 
.A(n_17674),
.B(n_10300),
.Y(n_17797)
);

OR2x2_ASAP7_75t_L g17798 ( 
.A(n_17542),
.B(n_10302),
.Y(n_17798)
);

AOI321xp33_ASAP7_75t_L g17799 ( 
.A1(n_17467),
.A2(n_7298),
.A3(n_7081),
.B1(n_7342),
.B2(n_7296),
.C(n_6942),
.Y(n_17799)
);

INVx1_ASAP7_75t_L g17800 ( 
.A(n_17511),
.Y(n_17800)
);

INVx1_ASAP7_75t_L g17801 ( 
.A(n_17514),
.Y(n_17801)
);

OAI32xp33_ASAP7_75t_SL g17802 ( 
.A1(n_17642),
.A2(n_8087),
.A3(n_7874),
.B1(n_8535),
.B2(n_8336),
.Y(n_17802)
);

INVx1_ASAP7_75t_L g17803 ( 
.A(n_17515),
.Y(n_17803)
);

OAI21xp5_ASAP7_75t_L g17804 ( 
.A1(n_17483),
.A2(n_7734),
.B(n_7733),
.Y(n_17804)
);

NAND2xp5_ASAP7_75t_SL g17805 ( 
.A(n_17536),
.B(n_8423),
.Y(n_17805)
);

INVxp33_ASAP7_75t_L g17806 ( 
.A(n_17376),
.Y(n_17806)
);

AND2x2_ASAP7_75t_L g17807 ( 
.A(n_17503),
.B(n_10302),
.Y(n_17807)
);

AOI22xp5_ASAP7_75t_L g17808 ( 
.A1(n_17501),
.A2(n_8423),
.B1(n_8581),
.B2(n_8463),
.Y(n_17808)
);

AOI322xp5_ASAP7_75t_L g17809 ( 
.A1(n_17636),
.A2(n_8463),
.A3(n_8581),
.B1(n_8743),
.B2(n_8943),
.C1(n_8844),
.C2(n_8689),
.Y(n_17809)
);

INVx1_ASAP7_75t_L g17810 ( 
.A(n_17368),
.Y(n_17810)
);

NAND2xp5_ASAP7_75t_L g17811 ( 
.A(n_17558),
.B(n_10307),
.Y(n_17811)
);

INVx1_ASAP7_75t_L g17812 ( 
.A(n_17464),
.Y(n_17812)
);

NAND2xp5_ASAP7_75t_L g17813 ( 
.A(n_17537),
.B(n_10307),
.Y(n_17813)
);

OAI21xp33_ASAP7_75t_L g17814 ( 
.A1(n_17667),
.A2(n_8581),
.B(n_8463),
.Y(n_17814)
);

INVx1_ASAP7_75t_L g17815 ( 
.A(n_17377),
.Y(n_17815)
);

NAND2xp5_ASAP7_75t_SL g17816 ( 
.A(n_17557),
.B(n_17548),
.Y(n_17816)
);

INVx1_ASAP7_75t_L g17817 ( 
.A(n_17472),
.Y(n_17817)
);

OAI33xp33_ASAP7_75t_L g17818 ( 
.A1(n_17518),
.A2(n_10324),
.A3(n_10309),
.B1(n_10330),
.B2(n_10326),
.B3(n_10310),
.Y(n_17818)
);

INVx1_ASAP7_75t_SL g17819 ( 
.A(n_17363),
.Y(n_17819)
);

AOI22xp33_ASAP7_75t_SL g17820 ( 
.A1(n_17473),
.A2(n_8463),
.B1(n_8689),
.B2(n_8581),
.Y(n_17820)
);

INVx1_ASAP7_75t_L g17821 ( 
.A(n_17477),
.Y(n_17821)
);

INVx1_ASAP7_75t_SL g17822 ( 
.A(n_17394),
.Y(n_17822)
);

AND2x2_ASAP7_75t_L g17823 ( 
.A(n_17587),
.B(n_10309),
.Y(n_17823)
);

INVx1_ASAP7_75t_L g17824 ( 
.A(n_17540),
.Y(n_17824)
);

BUFx2_ASAP7_75t_L g17825 ( 
.A(n_17484),
.Y(n_17825)
);

INVx1_ASAP7_75t_L g17826 ( 
.A(n_17544),
.Y(n_17826)
);

NAND2xp33_ASAP7_75t_L g17827 ( 
.A(n_17406),
.B(n_10310),
.Y(n_17827)
);

INVx1_ASAP7_75t_L g17828 ( 
.A(n_17517),
.Y(n_17828)
);

NAND2xp5_ASAP7_75t_L g17829 ( 
.A(n_17570),
.B(n_10324),
.Y(n_17829)
);

NAND2xp5_ASAP7_75t_L g17830 ( 
.A(n_17579),
.B(n_10326),
.Y(n_17830)
);

NAND2xp5_ASAP7_75t_L g17831 ( 
.A(n_17580),
.B(n_10330),
.Y(n_17831)
);

NAND2xp5_ASAP7_75t_L g17832 ( 
.A(n_17595),
.B(n_10331),
.Y(n_17832)
);

OR2x2_ASAP7_75t_L g17833 ( 
.A(n_17506),
.B(n_10331),
.Y(n_17833)
);

AOI22xp5_ASAP7_75t_L g17834 ( 
.A1(n_17654),
.A2(n_8463),
.B1(n_8689),
.B2(n_8581),
.Y(n_17834)
);

AND2x2_ASAP7_75t_L g17835 ( 
.A(n_17635),
.B(n_10334),
.Y(n_17835)
);

AOI21xp33_ASAP7_75t_L g17836 ( 
.A1(n_17554),
.A2(n_10150),
.B(n_10104),
.Y(n_17836)
);

OA21x2_ASAP7_75t_L g17837 ( 
.A1(n_17621),
.A2(n_10036),
.B(n_10334),
.Y(n_17837)
);

OR2x2_ASAP7_75t_L g17838 ( 
.A(n_17424),
.B(n_10335),
.Y(n_17838)
);

INVx2_ASAP7_75t_L g17839 ( 
.A(n_17555),
.Y(n_17839)
);

AOI322xp5_ASAP7_75t_L g17840 ( 
.A1(n_17479),
.A2(n_8689),
.A3(n_8743),
.B1(n_8943),
.B2(n_9004),
.C1(n_8844),
.C2(n_8963),
.Y(n_17840)
);

AND2x2_ASAP7_75t_L g17841 ( 
.A(n_17643),
.B(n_10335),
.Y(n_17841)
);

OAI31xp33_ASAP7_75t_L g17842 ( 
.A1(n_17497),
.A2(n_8963),
.A3(n_8569),
.B(n_8585),
.Y(n_17842)
);

AOI22xp33_ASAP7_75t_L g17843 ( 
.A1(n_17670),
.A2(n_8369),
.B1(n_8317),
.B2(n_8227),
.Y(n_17843)
);

OAI21xp5_ASAP7_75t_L g17844 ( 
.A1(n_17584),
.A2(n_7734),
.B(n_7733),
.Y(n_17844)
);

OAI322xp33_ASAP7_75t_L g17845 ( 
.A1(n_17507),
.A2(n_17513),
.A3(n_17423),
.B1(n_17437),
.B2(n_17378),
.C1(n_17415),
.C2(n_17675),
.Y(n_17845)
);

NAND2xp5_ASAP7_75t_L g17846 ( 
.A(n_17641),
.B(n_10336),
.Y(n_17846)
);

OAI21xp5_ASAP7_75t_SL g17847 ( 
.A1(n_17639),
.A2(n_8569),
.B(n_8366),
.Y(n_17847)
);

OAI21xp33_ASAP7_75t_SL g17848 ( 
.A1(n_17583),
.A2(n_10338),
.B(n_10336),
.Y(n_17848)
);

AND2x2_ASAP7_75t_L g17849 ( 
.A(n_17640),
.B(n_10338),
.Y(n_17849)
);

NOR2xp33_ASAP7_75t_L g17850 ( 
.A(n_17637),
.B(n_8689),
.Y(n_17850)
);

NAND3xp33_ASAP7_75t_SL g17851 ( 
.A(n_17602),
.B(n_8585),
.C(n_8366),
.Y(n_17851)
);

OAI22xp5_ASAP7_75t_L g17852 ( 
.A1(n_17504),
.A2(n_10343),
.B1(n_10346),
.B2(n_10342),
.Y(n_17852)
);

INVx1_ASAP7_75t_SL g17853 ( 
.A(n_17632),
.Y(n_17853)
);

AOI221xp5_ASAP7_75t_L g17854 ( 
.A1(n_17586),
.A2(n_8943),
.B1(n_9004),
.B2(n_8844),
.C(n_8743),
.Y(n_17854)
);

AND2x4_ASAP7_75t_L g17855 ( 
.A(n_17599),
.B(n_10342),
.Y(n_17855)
);

NAND2xp5_ASAP7_75t_L g17856 ( 
.A(n_17646),
.B(n_10343),
.Y(n_17856)
);

INVx1_ASAP7_75t_L g17857 ( 
.A(n_17402),
.Y(n_17857)
);

INVx1_ASAP7_75t_L g17858 ( 
.A(n_17521),
.Y(n_17858)
);

INVx1_ASAP7_75t_L g17859 ( 
.A(n_17380),
.Y(n_17859)
);

NAND2xp5_ASAP7_75t_L g17860 ( 
.A(n_17650),
.B(n_17553),
.Y(n_17860)
);

INVx1_ASAP7_75t_L g17861 ( 
.A(n_17505),
.Y(n_17861)
);

INVx1_ASAP7_75t_L g17862 ( 
.A(n_17532),
.Y(n_17862)
);

INVx1_ASAP7_75t_L g17863 ( 
.A(n_17465),
.Y(n_17863)
);

INVx1_ASAP7_75t_L g17864 ( 
.A(n_17460),
.Y(n_17864)
);

AND2x2_ASAP7_75t_L g17865 ( 
.A(n_17614),
.B(n_10346),
.Y(n_17865)
);

AND2x2_ASAP7_75t_L g17866 ( 
.A(n_17644),
.B(n_10356),
.Y(n_17866)
);

INVxp67_ASAP7_75t_SL g17867 ( 
.A(n_17576),
.Y(n_17867)
);

INVx1_ASAP7_75t_L g17868 ( 
.A(n_17414),
.Y(n_17868)
);

OAI21xp33_ASAP7_75t_L g17869 ( 
.A1(n_17663),
.A2(n_8844),
.B(n_8743),
.Y(n_17869)
);

A2O1A1Ixp33_ASAP7_75t_L g17870 ( 
.A1(n_17577),
.A2(n_10359),
.B(n_10362),
.C(n_10356),
.Y(n_17870)
);

AOI21xp5_ASAP7_75t_L g17871 ( 
.A1(n_17627),
.A2(n_17563),
.B(n_17561),
.Y(n_17871)
);

INVx1_ASAP7_75t_L g17872 ( 
.A(n_17673),
.Y(n_17872)
);

AOI21xp5_ASAP7_75t_L g17873 ( 
.A1(n_17655),
.A2(n_10362),
.B(n_10359),
.Y(n_17873)
);

NAND2xp5_ASAP7_75t_L g17874 ( 
.A(n_17676),
.B(n_10366),
.Y(n_17874)
);

INVx1_ASAP7_75t_L g17875 ( 
.A(n_17381),
.Y(n_17875)
);

OAI22xp5_ASAP7_75t_L g17876 ( 
.A1(n_17439),
.A2(n_10374),
.B1(n_10379),
.B2(n_10366),
.Y(n_17876)
);

O2A1O1Ixp5_ASAP7_75t_L g17877 ( 
.A1(n_17556),
.A2(n_10379),
.B(n_10380),
.C(n_10374),
.Y(n_17877)
);

AND2x2_ASAP7_75t_L g17878 ( 
.A(n_17569),
.B(n_17572),
.Y(n_17878)
);

OAI32xp33_ASAP7_75t_L g17879 ( 
.A1(n_17522),
.A2(n_8943),
.A3(n_9004),
.B1(n_8844),
.B2(n_8743),
.Y(n_17879)
);

AND2x4_ASAP7_75t_L g17880 ( 
.A(n_17589),
.B(n_10380),
.Y(n_17880)
);

AOI22xp5_ASAP7_75t_L g17881 ( 
.A1(n_17677),
.A2(n_9004),
.B1(n_8943),
.B2(n_10381),
.Y(n_17881)
);

NOR2xp33_ASAP7_75t_L g17882 ( 
.A(n_17613),
.B(n_9004),
.Y(n_17882)
);

INVx2_ASAP7_75t_L g17883 ( 
.A(n_17669),
.Y(n_17883)
);

AND2x2_ASAP7_75t_L g17884 ( 
.A(n_17656),
.B(n_10381),
.Y(n_17884)
);

NAND2xp5_ASAP7_75t_L g17885 ( 
.A(n_17496),
.B(n_10104),
.Y(n_17885)
);

OAI32xp33_ASAP7_75t_L g17886 ( 
.A1(n_17534),
.A2(n_8681),
.A3(n_8797),
.B1(n_8661),
.B2(n_8585),
.Y(n_17886)
);

OAI21xp5_ASAP7_75t_L g17887 ( 
.A1(n_17665),
.A2(n_8178),
.B(n_8177),
.Y(n_17887)
);

AND2x2_ASAP7_75t_L g17888 ( 
.A(n_17574),
.B(n_8121),
.Y(n_17888)
);

AOI21xp33_ASAP7_75t_L g17889 ( 
.A1(n_17672),
.A2(n_10150),
.B(n_9808),
.Y(n_17889)
);

NAND2xp5_ASAP7_75t_L g17890 ( 
.A(n_17664),
.B(n_9808),
.Y(n_17890)
);

OAI221xp5_ASAP7_75t_L g17891 ( 
.A1(n_17440),
.A2(n_17407),
.B1(n_17560),
.B2(n_17509),
.C(n_17607),
.Y(n_17891)
);

INVx1_ASAP7_75t_L g17892 ( 
.A(n_17492),
.Y(n_17892)
);

INVx1_ASAP7_75t_L g17893 ( 
.A(n_17488),
.Y(n_17893)
);

NOR3xp33_ASAP7_75t_L g17894 ( 
.A(n_17678),
.B(n_8042),
.C(n_8041),
.Y(n_17894)
);

AOI21xp5_ASAP7_75t_L g17895 ( 
.A1(n_17657),
.A2(n_9808),
.B(n_9757),
.Y(n_17895)
);

AND2x2_ASAP7_75t_L g17896 ( 
.A(n_17578),
.B(n_8121),
.Y(n_17896)
);

INVx1_ASAP7_75t_L g17897 ( 
.A(n_17392),
.Y(n_17897)
);

INVx1_ASAP7_75t_L g17898 ( 
.A(n_17588),
.Y(n_17898)
);

OAI22xp33_ASAP7_75t_L g17899 ( 
.A1(n_17573),
.A2(n_7772),
.B1(n_7872),
.B2(n_7717),
.Y(n_17899)
);

INVx1_ASAP7_75t_L g17900 ( 
.A(n_17445),
.Y(n_17900)
);

NOR2xp33_ASAP7_75t_SL g17901 ( 
.A(n_17661),
.B(n_8661),
.Y(n_17901)
);

INVx1_ASAP7_75t_L g17902 ( 
.A(n_17592),
.Y(n_17902)
);

NAND2xp5_ASAP7_75t_L g17903 ( 
.A(n_17653),
.B(n_9808),
.Y(n_17903)
);

INVx1_ASAP7_75t_L g17904 ( 
.A(n_17447),
.Y(n_17904)
);

INVx1_ASAP7_75t_L g17905 ( 
.A(n_17469),
.Y(n_17905)
);

INVx1_ASAP7_75t_L g17906 ( 
.A(n_17499),
.Y(n_17906)
);

OAI22xp33_ASAP7_75t_L g17907 ( 
.A1(n_17633),
.A2(n_7772),
.B1(n_7925),
.B2(n_7717),
.Y(n_17907)
);

OAI21xp5_ASAP7_75t_L g17908 ( 
.A1(n_17671),
.A2(n_8178),
.B(n_8177),
.Y(n_17908)
);

INVx1_ASAP7_75t_L g17909 ( 
.A(n_17622),
.Y(n_17909)
);

NAND2xp5_ASAP7_75t_L g17910 ( 
.A(n_17601),
.B(n_9484),
.Y(n_17910)
);

NAND3xp33_ASAP7_75t_L g17911 ( 
.A(n_17603),
.B(n_17617),
.C(n_17605),
.Y(n_17911)
);

INVx2_ASAP7_75t_L g17912 ( 
.A(n_17425),
.Y(n_17912)
);

NAND2xp5_ASAP7_75t_L g17913 ( 
.A(n_17606),
.B(n_9484),
.Y(n_17913)
);

NAND2xp5_ASAP7_75t_L g17914 ( 
.A(n_17608),
.B(n_9484),
.Y(n_17914)
);

INVx1_ASAP7_75t_L g17915 ( 
.A(n_17510),
.Y(n_17915)
);

INVx1_ASAP7_75t_L g17916 ( 
.A(n_17516),
.Y(n_17916)
);

HB1xp67_ASAP7_75t_L g17917 ( 
.A(n_17495),
.Y(n_17917)
);

OAI22xp5_ASAP7_75t_L g17918 ( 
.A1(n_17435),
.A2(n_8440),
.B1(n_7929),
.B2(n_7981),
.Y(n_17918)
);

AOI22xp5_ASAP7_75t_L g17919 ( 
.A1(n_17413),
.A2(n_9757),
.B1(n_9484),
.B2(n_8841),
.Y(n_17919)
);

INVxp67_ASAP7_75t_L g17920 ( 
.A(n_17604),
.Y(n_17920)
);

INVx2_ASAP7_75t_L g17921 ( 
.A(n_17426),
.Y(n_17921)
);

NAND2xp5_ASAP7_75t_SL g17922 ( 
.A(n_17384),
.B(n_8440),
.Y(n_17922)
);

AND2x2_ASAP7_75t_L g17923 ( 
.A(n_17615),
.B(n_8121),
.Y(n_17923)
);

NAND3xp33_ASAP7_75t_L g17924 ( 
.A(n_17623),
.B(n_8369),
.C(n_8317),
.Y(n_17924)
);

AND2x2_ASAP7_75t_L g17925 ( 
.A(n_17624),
.B(n_8121),
.Y(n_17925)
);

NAND3xp33_ASAP7_75t_SL g17926 ( 
.A(n_17631),
.B(n_8681),
.C(n_8661),
.Y(n_17926)
);

INVx1_ASAP7_75t_L g17927 ( 
.A(n_17645),
.Y(n_17927)
);

AOI221x1_ASAP7_75t_L g17928 ( 
.A1(n_17638),
.A2(n_8745),
.B1(n_8747),
.B2(n_8740),
.C(n_8735),
.Y(n_17928)
);

OAI21xp33_ASAP7_75t_L g17929 ( 
.A1(n_17422),
.A2(n_7929),
.B(n_7925),
.Y(n_17929)
);

AOI21xp33_ASAP7_75t_L g17930 ( 
.A1(n_17647),
.A2(n_9757),
.B(n_9862),
.Y(n_17930)
);

BUFx2_ASAP7_75t_L g17931 ( 
.A(n_17390),
.Y(n_17931)
);

INVx1_ASAP7_75t_L g17932 ( 
.A(n_17596),
.Y(n_17932)
);

OAI21xp5_ASAP7_75t_L g17933 ( 
.A1(n_17651),
.A2(n_8178),
.B(n_8177),
.Y(n_17933)
);

INVx1_ASAP7_75t_L g17934 ( 
.A(n_17582),
.Y(n_17934)
);

OAI31xp33_ASAP7_75t_L g17935 ( 
.A1(n_17404),
.A2(n_8681),
.A3(n_8797),
.B(n_8661),
.Y(n_17935)
);

OR2x2_ASAP7_75t_L g17936 ( 
.A(n_17559),
.B(n_7874),
.Y(n_17936)
);

AOI21xp33_ASAP7_75t_SL g17937 ( 
.A1(n_17408),
.A2(n_8369),
.B(n_8317),
.Y(n_17937)
);

AOI22xp5_ASAP7_75t_L g17938 ( 
.A1(n_17412),
.A2(n_9757),
.B1(n_8841),
.B2(n_8975),
.Y(n_17938)
);

INVx1_ASAP7_75t_L g17939 ( 
.A(n_17600),
.Y(n_17939)
);

INVx1_ASAP7_75t_SL g17940 ( 
.A(n_17668),
.Y(n_17940)
);

NAND2xp5_ASAP7_75t_L g17941 ( 
.A(n_17616),
.B(n_9862),
.Y(n_17941)
);

INVx2_ASAP7_75t_SL g17942 ( 
.A(n_17611),
.Y(n_17942)
);

INVx1_ASAP7_75t_L g17943 ( 
.A(n_17618),
.Y(n_17943)
);

NAND3xp33_ASAP7_75t_SL g17944 ( 
.A(n_17662),
.B(n_8814),
.C(n_8797),
.Y(n_17944)
);

AOI222xp33_ASAP7_75t_L g17945 ( 
.A1(n_17629),
.A2(n_7805),
.B1(n_7812),
.B2(n_7858),
.C1(n_7852),
.C2(n_7836),
.Y(n_17945)
);

INVx1_ASAP7_75t_L g17946 ( 
.A(n_17626),
.Y(n_17946)
);

AND2x2_ASAP7_75t_L g17947 ( 
.A(n_17571),
.B(n_8121),
.Y(n_17947)
);

NAND4xp25_ASAP7_75t_L g17948 ( 
.A(n_17666),
.B(n_6939),
.C(n_6950),
.D(n_6912),
.Y(n_17948)
);

NOR2xp33_ASAP7_75t_L g17949 ( 
.A(n_17649),
.B(n_7376),
.Y(n_17949)
);

NAND3x2_ASAP7_75t_L g17950 ( 
.A(n_17691),
.B(n_17385),
.C(n_17648),
.Y(n_17950)
);

AOI222xp33_ASAP7_75t_L g17951 ( 
.A1(n_17720),
.A2(n_17625),
.B1(n_17432),
.B2(n_17388),
.C1(n_17597),
.C2(n_17535),
.Y(n_17951)
);

INVxp67_ASAP7_75t_L g17952 ( 
.A(n_17785),
.Y(n_17952)
);

AOI21xp5_ASAP7_75t_L g17953 ( 
.A1(n_17692),
.A2(n_17867),
.B(n_17709),
.Y(n_17953)
);

INVx1_ASAP7_75t_L g17954 ( 
.A(n_17697),
.Y(n_17954)
);

NAND2xp5_ASAP7_75t_L g17955 ( 
.A(n_17724),
.B(n_17543),
.Y(n_17955)
);

O2A1O1Ixp33_ASAP7_75t_SL g17956 ( 
.A1(n_17942),
.A2(n_17630),
.B(n_17527),
.C(n_17598),
.Y(n_17956)
);

INVx1_ASAP7_75t_SL g17957 ( 
.A(n_17737),
.Y(n_17957)
);

NAND2xp5_ASAP7_75t_L g17958 ( 
.A(n_17706),
.B(n_17630),
.Y(n_17958)
);

AOI22xp5_ASAP7_75t_L g17959 ( 
.A1(n_17699),
.A2(n_8841),
.B1(n_8975),
.B2(n_8870),
.Y(n_17959)
);

NAND2xp5_ASAP7_75t_L g17960 ( 
.A(n_17712),
.B(n_9862),
.Y(n_17960)
);

INVx1_ASAP7_75t_L g17961 ( 
.A(n_17680),
.Y(n_17961)
);

OAI22xp5_ASAP7_75t_L g17962 ( 
.A1(n_17723),
.A2(n_7981),
.B1(n_7925),
.B2(n_8797),
.Y(n_17962)
);

OAI21xp5_ASAP7_75t_SL g17963 ( 
.A1(n_17687),
.A2(n_8935),
.B(n_8814),
.Y(n_17963)
);

AOI31xp33_ASAP7_75t_L g17964 ( 
.A1(n_17806),
.A2(n_8973),
.A3(n_9006),
.B(n_8935),
.Y(n_17964)
);

NAND2xp5_ASAP7_75t_L g17965 ( 
.A(n_17810),
.B(n_9862),
.Y(n_17965)
);

AOI221xp5_ASAP7_75t_L g17966 ( 
.A1(n_17705),
.A2(n_6765),
.B1(n_6761),
.B2(n_6749),
.C(n_8609),
.Y(n_17966)
);

OR2x2_ASAP7_75t_L g17967 ( 
.A(n_17721),
.B(n_7874),
.Y(n_17967)
);

AOI22xp5_ASAP7_75t_L g17968 ( 
.A1(n_17710),
.A2(n_8870),
.B1(n_8975),
.B2(n_8369),
.Y(n_17968)
);

NAND3xp33_ASAP7_75t_SL g17969 ( 
.A(n_17703),
.B(n_8973),
.C(n_8935),
.Y(n_17969)
);

AND2x2_ASAP7_75t_L g17970 ( 
.A(n_17714),
.B(n_8121),
.Y(n_17970)
);

INVx1_ASAP7_75t_L g17971 ( 
.A(n_17825),
.Y(n_17971)
);

OA21x2_ASAP7_75t_L g17972 ( 
.A1(n_17909),
.A2(n_10036),
.B(n_8583),
.Y(n_17972)
);

NOR2xp33_ASAP7_75t_R g17973 ( 
.A(n_17731),
.B(n_5834),
.Y(n_17973)
);

NAND2xp5_ASAP7_75t_SL g17974 ( 
.A(n_17695),
.B(n_17740),
.Y(n_17974)
);

INVx2_ASAP7_75t_L g17975 ( 
.A(n_17683),
.Y(n_17975)
);

INVx1_ASAP7_75t_SL g17976 ( 
.A(n_17853),
.Y(n_17976)
);

INVx1_ASAP7_75t_L g17977 ( 
.A(n_17696),
.Y(n_17977)
);

OAI322xp33_ASAP7_75t_L g17978 ( 
.A1(n_17793),
.A2(n_7981),
.A3(n_8763),
.B1(n_8925),
.B2(n_8774),
.C1(n_6749),
.C2(n_6765),
.Y(n_17978)
);

NAND2xp5_ASAP7_75t_SL g17979 ( 
.A(n_17748),
.B(n_8973),
.Y(n_17979)
);

INVx2_ASAP7_75t_L g17980 ( 
.A(n_17708),
.Y(n_17980)
);

INVx1_ASAP7_75t_L g17981 ( 
.A(n_17688),
.Y(n_17981)
);

INVx1_ASAP7_75t_L g17982 ( 
.A(n_17694),
.Y(n_17982)
);

AOI32xp33_ASAP7_75t_L g17983 ( 
.A1(n_17819),
.A2(n_8475),
.A3(n_8482),
.B1(n_8466),
.B2(n_8456),
.Y(n_17983)
);

OAI22xp5_ASAP7_75t_L g17984 ( 
.A1(n_17774),
.A2(n_9006),
.B1(n_8973),
.B2(n_8763),
.Y(n_17984)
);

AOI21xp33_ASAP7_75t_L g17985 ( 
.A1(n_17722),
.A2(n_8522),
.B(n_7812),
.Y(n_17985)
);

NOR2xp33_ASAP7_75t_L g17986 ( 
.A(n_17824),
.B(n_7376),
.Y(n_17986)
);

AND2x2_ASAP7_75t_L g17987 ( 
.A(n_17713),
.B(n_8121),
.Y(n_17987)
);

NAND2xp5_ASAP7_75t_L g17988 ( 
.A(n_17733),
.B(n_8677),
.Y(n_17988)
);

NOR2x1_ASAP7_75t_L g17989 ( 
.A(n_17690),
.B(n_8609),
.Y(n_17989)
);

AND2x2_ASAP7_75t_L g17990 ( 
.A(n_17878),
.B(n_8121),
.Y(n_17990)
);

INVx1_ASAP7_75t_L g17991 ( 
.A(n_17727),
.Y(n_17991)
);

OAI21xp33_ASAP7_75t_L g17992 ( 
.A1(n_17682),
.A2(n_8774),
.B(n_8763),
.Y(n_17992)
);

NOR3xp33_ASAP7_75t_L g17993 ( 
.A(n_17764),
.B(n_5287),
.C(n_5197),
.Y(n_17993)
);

INVx1_ASAP7_75t_L g17994 ( 
.A(n_17704),
.Y(n_17994)
);

INVx1_ASAP7_75t_SL g17995 ( 
.A(n_17776),
.Y(n_17995)
);

INVxp67_ASAP7_75t_L g17996 ( 
.A(n_17716),
.Y(n_17996)
);

OAI22xp5_ASAP7_75t_L g17997 ( 
.A1(n_17746),
.A2(n_9006),
.B1(n_8774),
.B2(n_8925),
.Y(n_17997)
);

INVx1_ASAP7_75t_L g17998 ( 
.A(n_17685),
.Y(n_17998)
);

INVx2_ASAP7_75t_L g17999 ( 
.A(n_17754),
.Y(n_17999)
);

AOI21xp33_ASAP7_75t_SL g18000 ( 
.A1(n_17932),
.A2(n_8317),
.B(n_8227),
.Y(n_18000)
);

AOI32xp33_ASAP7_75t_L g18001 ( 
.A1(n_17772),
.A2(n_8475),
.A3(n_8482),
.B1(n_8466),
.B2(n_8456),
.Y(n_18001)
);

OR2x2_ASAP7_75t_L g18002 ( 
.A(n_17826),
.B(n_7874),
.Y(n_18002)
);

NOR2xp33_ASAP7_75t_L g18003 ( 
.A(n_17780),
.B(n_7376),
.Y(n_18003)
);

NOR2xp33_ASAP7_75t_L g18004 ( 
.A(n_17769),
.B(n_7376),
.Y(n_18004)
);

INVx1_ASAP7_75t_L g18005 ( 
.A(n_17698),
.Y(n_18005)
);

INVx1_ASAP7_75t_SL g18006 ( 
.A(n_17940),
.Y(n_18006)
);

NAND4xp25_ASAP7_75t_SL g18007 ( 
.A(n_17719),
.B(n_8925),
.C(n_7124),
.D(n_7425),
.Y(n_18007)
);

INVx1_ASAP7_75t_L g18008 ( 
.A(n_17701),
.Y(n_18008)
);

NAND3xp33_ASAP7_75t_L g18009 ( 
.A(n_17679),
.B(n_8317),
.C(n_8227),
.Y(n_18009)
);

NAND2xp5_ASAP7_75t_L g18010 ( 
.A(n_17777),
.B(n_8677),
.Y(n_18010)
);

NAND3xp33_ASAP7_75t_L g18011 ( 
.A(n_17700),
.B(n_8317),
.C(n_8227),
.Y(n_18011)
);

OAI221xp5_ASAP7_75t_L g18012 ( 
.A1(n_17686),
.A2(n_9006),
.B1(n_7244),
.B2(n_7570),
.C(n_7301),
.Y(n_18012)
);

OAI21xp5_ASAP7_75t_L g18013 ( 
.A1(n_17871),
.A2(n_8042),
.B(n_8041),
.Y(n_18013)
);

AND2x4_ASAP7_75t_L g18014 ( 
.A(n_17883),
.B(n_7993),
.Y(n_18014)
);

INVx1_ASAP7_75t_L g18015 ( 
.A(n_17757),
.Y(n_18015)
);

INVx1_ASAP7_75t_L g18016 ( 
.A(n_17702),
.Y(n_18016)
);

AOI22xp33_ASAP7_75t_SL g18017 ( 
.A1(n_17789),
.A2(n_8369),
.B1(n_8227),
.B2(n_7376),
.Y(n_18017)
);

OA21x2_ASAP7_75t_L g18018 ( 
.A1(n_17860),
.A2(n_10036),
.B(n_8583),
.Y(n_18018)
);

AND2x2_ASAP7_75t_L g18019 ( 
.A(n_17839),
.B(n_8264),
.Y(n_18019)
);

NOR2xp33_ASAP7_75t_L g18020 ( 
.A(n_17765),
.B(n_7573),
.Y(n_18020)
);

INVx1_ASAP7_75t_L g18021 ( 
.A(n_17931),
.Y(n_18021)
);

INVx1_ASAP7_75t_L g18022 ( 
.A(n_17707),
.Y(n_18022)
);

INVx2_ASAP7_75t_L g18023 ( 
.A(n_17742),
.Y(n_18023)
);

INVx1_ASAP7_75t_L g18024 ( 
.A(n_17755),
.Y(n_18024)
);

AOI32xp33_ASAP7_75t_L g18025 ( 
.A1(n_17767),
.A2(n_8482),
.A3(n_8492),
.B1(n_8475),
.B2(n_8466),
.Y(n_18025)
);

OAI21xp33_ASAP7_75t_L g18026 ( 
.A1(n_17949),
.A2(n_7034),
.B(n_7015),
.Y(n_18026)
);

AOI21xp5_ASAP7_75t_L g18027 ( 
.A1(n_17816),
.A2(n_8522),
.B(n_7812),
.Y(n_18027)
);

OR2x2_ASAP7_75t_L g18028 ( 
.A(n_17812),
.B(n_7874),
.Y(n_18028)
);

NAND2xp5_ASAP7_75t_L g18029 ( 
.A(n_17745),
.B(n_8677),
.Y(n_18029)
);

INVx2_ASAP7_75t_L g18030 ( 
.A(n_17807),
.Y(n_18030)
);

OAI222xp33_ASAP7_75t_L g18031 ( 
.A1(n_17758),
.A2(n_6633),
.B1(n_6627),
.B2(n_6762),
.C1(n_6700),
.C2(n_6630),
.Y(n_18031)
);

INVx1_ASAP7_75t_L g18032 ( 
.A(n_17866),
.Y(n_18032)
);

OR2x2_ASAP7_75t_L g18033 ( 
.A(n_17792),
.B(n_7874),
.Y(n_18033)
);

NOR2xp33_ASAP7_75t_L g18034 ( 
.A(n_17689),
.B(n_7573),
.Y(n_18034)
);

AND2x2_ASAP7_75t_L g18035 ( 
.A(n_17800),
.B(n_8264),
.Y(n_18035)
);

OAI21xp5_ASAP7_75t_L g18036 ( 
.A1(n_17911),
.A2(n_17684),
.B(n_17920),
.Y(n_18036)
);

AOI21xp33_ASAP7_75t_SL g18037 ( 
.A1(n_17715),
.A2(n_8227),
.B(n_7975),
.Y(n_18037)
);

OAI322xp33_ASAP7_75t_L g18038 ( 
.A1(n_17717),
.A2(n_6761),
.A3(n_6700),
.B1(n_6630),
.B2(n_6762),
.C1(n_6633),
.C2(n_6627),
.Y(n_18038)
);

NOR3xp33_ASAP7_75t_SL g18039 ( 
.A(n_17845),
.B(n_6661),
.C(n_6955),
.Y(n_18039)
);

AOI21xp5_ASAP7_75t_L g18040 ( 
.A1(n_17872),
.A2(n_17718),
.B(n_17753),
.Y(n_18040)
);

AOI222xp33_ASAP7_75t_L g18041 ( 
.A1(n_17827),
.A2(n_7805),
.B1(n_7858),
.B2(n_7852),
.C1(n_8583),
.C2(n_7836),
.Y(n_18041)
);

OAI22xp5_ASAP7_75t_L g18042 ( 
.A1(n_17750),
.A2(n_6627),
.B1(n_6633),
.B2(n_6630),
.Y(n_18042)
);

AOI21xp33_ASAP7_75t_SL g18043 ( 
.A1(n_17711),
.A2(n_7975),
.B(n_8609),
.Y(n_18043)
);

AND2x2_ASAP7_75t_L g18044 ( 
.A(n_17801),
.B(n_8264),
.Y(n_18044)
);

NAND2xp5_ASAP7_75t_L g18045 ( 
.A(n_17803),
.B(n_8677),
.Y(n_18045)
);

NOR2xp33_ASAP7_75t_L g18046 ( 
.A(n_17822),
.B(n_7573),
.Y(n_18046)
);

AOI221xp5_ASAP7_75t_L g18047 ( 
.A1(n_17693),
.A2(n_8624),
.B1(n_8609),
.B2(n_8501),
.C(n_8677),
.Y(n_18047)
);

OAI322xp33_ASAP7_75t_L g18048 ( 
.A1(n_17768),
.A2(n_6700),
.A3(n_6630),
.B1(n_6762),
.B2(n_6784),
.C1(n_6633),
.C2(n_6627),
.Y(n_18048)
);

OAI21xp5_ASAP7_75t_L g18049 ( 
.A1(n_17762),
.A2(n_8042),
.B(n_8041),
.Y(n_18049)
);

NAND4xp25_ASAP7_75t_L g18050 ( 
.A(n_17681),
.B(n_6939),
.C(n_6950),
.D(n_6912),
.Y(n_18050)
);

INVx1_ASAP7_75t_L g18051 ( 
.A(n_17763),
.Y(n_18051)
);

INVx1_ASAP7_75t_L g18052 ( 
.A(n_17917),
.Y(n_18052)
);

OR2x2_ASAP7_75t_L g18053 ( 
.A(n_17912),
.B(n_7874),
.Y(n_18053)
);

AND2x2_ASAP7_75t_L g18054 ( 
.A(n_17921),
.B(n_8264),
.Y(n_18054)
);

NAND2xp5_ASAP7_75t_L g18055 ( 
.A(n_17858),
.B(n_8728),
.Y(n_18055)
);

INVx1_ASAP7_75t_L g18056 ( 
.A(n_17865),
.Y(n_18056)
);

NAND3xp33_ASAP7_75t_L g18057 ( 
.A(n_17770),
.B(n_7975),
.C(n_5083),
.Y(n_18057)
);

AOI211xp5_ASAP7_75t_L g18058 ( 
.A1(n_17817),
.A2(n_7244),
.B(n_7301),
.C(n_7198),
.Y(n_18058)
);

AOI21xp5_ASAP7_75t_L g18059 ( 
.A1(n_17857),
.A2(n_8522),
.B(n_7805),
.Y(n_18059)
);

NAND2xp5_ASAP7_75t_L g18060 ( 
.A(n_17821),
.B(n_8728),
.Y(n_18060)
);

AOI32xp33_ASAP7_75t_L g18061 ( 
.A1(n_17782),
.A2(n_8498),
.A3(n_8502),
.B1(n_8493),
.B2(n_8492),
.Y(n_18061)
);

NAND2xp5_ASAP7_75t_L g18062 ( 
.A(n_17761),
.B(n_8728),
.Y(n_18062)
);

OAI22xp5_ASAP7_75t_SL g18063 ( 
.A1(n_17828),
.A2(n_7573),
.B1(n_7244),
.B2(n_7301),
.Y(n_18063)
);

INVx2_ASAP7_75t_L g18064 ( 
.A(n_17781),
.Y(n_18064)
);

NAND2xp5_ASAP7_75t_L g18065 ( 
.A(n_17892),
.B(n_8728),
.Y(n_18065)
);

NAND2xp5_ASAP7_75t_L g18066 ( 
.A(n_17893),
.B(n_8728),
.Y(n_18066)
);

NOR2xp33_ASAP7_75t_L g18067 ( 
.A(n_17732),
.B(n_7573),
.Y(n_18067)
);

AOI21xp33_ASAP7_75t_SL g18068 ( 
.A1(n_17861),
.A2(n_8624),
.B(n_8609),
.Y(n_18068)
);

OR3x2_ASAP7_75t_L g18069 ( 
.A(n_17864),
.B(n_17902),
.C(n_17898),
.Y(n_18069)
);

OR2x2_ASAP7_75t_L g18070 ( 
.A(n_17796),
.B(n_7874),
.Y(n_18070)
);

OAI21xp5_ASAP7_75t_L g18071 ( 
.A1(n_17749),
.A2(n_7724),
.B(n_7706),
.Y(n_18071)
);

INVx1_ASAP7_75t_L g18072 ( 
.A(n_17791),
.Y(n_18072)
);

NOR2xp67_ASAP7_75t_L g18073 ( 
.A(n_17862),
.B(n_8740),
.Y(n_18073)
);

OAI22xp5_ASAP7_75t_L g18074 ( 
.A1(n_17787),
.A2(n_6762),
.B1(n_6784),
.B2(n_6700),
.Y(n_18074)
);

HB1xp67_ASAP7_75t_L g18075 ( 
.A(n_17760),
.Y(n_18075)
);

INVxp67_ASAP7_75t_L g18076 ( 
.A(n_17850),
.Y(n_18076)
);

INVx1_ASAP7_75t_L g18077 ( 
.A(n_17795),
.Y(n_18077)
);

NAND4xp25_ASAP7_75t_L g18078 ( 
.A(n_17756),
.B(n_6939),
.C(n_6950),
.D(n_6912),
.Y(n_18078)
);

INVx1_ASAP7_75t_L g18079 ( 
.A(n_17798),
.Y(n_18079)
);

INVx1_ASAP7_75t_L g18080 ( 
.A(n_17784),
.Y(n_18080)
);

AOI222xp33_ASAP7_75t_L g18081 ( 
.A1(n_17922),
.A2(n_7836),
.B1(n_7847),
.B2(n_7842),
.C1(n_8613),
.C2(n_7987),
.Y(n_18081)
);

INVx1_ASAP7_75t_L g18082 ( 
.A(n_17797),
.Y(n_18082)
);

INVx1_ASAP7_75t_L g18083 ( 
.A(n_17813),
.Y(n_18083)
);

NOR4xp25_ASAP7_75t_L g18084 ( 
.A(n_17891),
.B(n_17863),
.C(n_17815),
.D(n_17859),
.Y(n_18084)
);

AND2x2_ASAP7_75t_L g18085 ( 
.A(n_17897),
.B(n_8264),
.Y(n_18085)
);

NAND2xp5_ASAP7_75t_L g18086 ( 
.A(n_17794),
.B(n_8522),
.Y(n_18086)
);

NOR2xp33_ASAP7_75t_L g18087 ( 
.A(n_17868),
.B(n_7573),
.Y(n_18087)
);

INVx1_ASAP7_75t_L g18088 ( 
.A(n_17739),
.Y(n_18088)
);

INVx1_ASAP7_75t_L g18089 ( 
.A(n_17829),
.Y(n_18089)
);

AOI21xp5_ASAP7_75t_SL g18090 ( 
.A1(n_17906),
.A2(n_7669),
.B(n_6706),
.Y(n_18090)
);

NAND2xp5_ASAP7_75t_L g18091 ( 
.A(n_17794),
.B(n_8522),
.Y(n_18091)
);

NAND4xp25_ASAP7_75t_L g18092 ( 
.A(n_17882),
.B(n_17725),
.C(n_17830),
.D(n_17934),
.Y(n_18092)
);

AOI31xp33_ASAP7_75t_L g18093 ( 
.A1(n_17875),
.A2(n_5350),
.A3(n_5465),
.B(n_5203),
.Y(n_18093)
);

INVx1_ASAP7_75t_L g18094 ( 
.A(n_17811),
.Y(n_18094)
);

INVx1_ASAP7_75t_L g18095 ( 
.A(n_17838),
.Y(n_18095)
);

NOR2xp33_ASAP7_75t_L g18096 ( 
.A(n_17939),
.B(n_7573),
.Y(n_18096)
);

INVx1_ASAP7_75t_L g18097 ( 
.A(n_17855),
.Y(n_18097)
);

NOR2x1_ASAP7_75t_L g18098 ( 
.A(n_17900),
.B(n_8624),
.Y(n_18098)
);

INVx1_ASAP7_75t_L g18099 ( 
.A(n_17855),
.Y(n_18099)
);

OAI22xp5_ASAP7_75t_L g18100 ( 
.A1(n_17726),
.A2(n_6791),
.B1(n_6892),
.B2(n_6784),
.Y(n_18100)
);

INVx1_ASAP7_75t_L g18101 ( 
.A(n_17880),
.Y(n_18101)
);

NOR2xp33_ASAP7_75t_L g18102 ( 
.A(n_17943),
.B(n_6912),
.Y(n_18102)
);

OAI22xp33_ASAP7_75t_L g18103 ( 
.A1(n_17901),
.A2(n_7225),
.B1(n_7254),
.B2(n_7199),
.Y(n_18103)
);

INVx1_ASAP7_75t_L g18104 ( 
.A(n_17880),
.Y(n_18104)
);

AOI22xp5_ASAP7_75t_L g18105 ( 
.A1(n_17734),
.A2(n_8975),
.B1(n_8870),
.B2(n_6784),
.Y(n_18105)
);

OAI32xp33_ASAP7_75t_L g18106 ( 
.A1(n_17874),
.A2(n_17903),
.A3(n_17904),
.B1(n_17915),
.B2(n_17905),
.Y(n_18106)
);

AND2x2_ASAP7_75t_L g18107 ( 
.A(n_17783),
.B(n_8264),
.Y(n_18107)
);

OR2x2_ASAP7_75t_L g18108 ( 
.A(n_17728),
.B(n_8264),
.Y(n_18108)
);

HB1xp67_ASAP7_75t_L g18109 ( 
.A(n_17916),
.Y(n_18109)
);

NAND2xp5_ASAP7_75t_L g18110 ( 
.A(n_17823),
.B(n_8624),
.Y(n_18110)
);

OAI221xp5_ASAP7_75t_L g18111 ( 
.A1(n_17738),
.A2(n_7301),
.B1(n_7570),
.B2(n_7244),
.C(n_7198),
.Y(n_18111)
);

INVx1_ASAP7_75t_L g18112 ( 
.A(n_17833),
.Y(n_18112)
);

OAI22xp5_ASAP7_75t_L g18113 ( 
.A1(n_17820),
.A2(n_6892),
.B1(n_6923),
.B2(n_6791),
.Y(n_18113)
);

OAI21xp33_ASAP7_75t_L g18114 ( 
.A1(n_17948),
.A2(n_7034),
.B(n_7015),
.Y(n_18114)
);

AOI22xp5_ASAP7_75t_L g18115 ( 
.A1(n_17923),
.A2(n_8975),
.B1(n_8870),
.B2(n_6791),
.Y(n_18115)
);

INVx1_ASAP7_75t_L g18116 ( 
.A(n_17832),
.Y(n_18116)
);

AND2x4_ASAP7_75t_L g18117 ( 
.A(n_17946),
.B(n_8557),
.Y(n_18117)
);

NAND2xp5_ASAP7_75t_L g18118 ( 
.A(n_17835),
.B(n_8624),
.Y(n_18118)
);

AOI22xp33_ASAP7_75t_L g18119 ( 
.A1(n_17929),
.A2(n_8975),
.B1(n_8501),
.B2(n_8454),
.Y(n_18119)
);

NAND2xp5_ASAP7_75t_L g18120 ( 
.A(n_17841),
.B(n_8501),
.Y(n_18120)
);

NOR4xp25_ASAP7_75t_SL g18121 ( 
.A(n_17927),
.B(n_6906),
.C(n_7004),
.D(n_7000),
.Y(n_18121)
);

OAI21xp5_ASAP7_75t_L g18122 ( 
.A1(n_17741),
.A2(n_7724),
.B(n_7706),
.Y(n_18122)
);

AND2x2_ASAP7_75t_L g18123 ( 
.A(n_17849),
.B(n_8264),
.Y(n_18123)
);

OAI22xp5_ASAP7_75t_L g18124 ( 
.A1(n_17918),
.A2(n_6892),
.B1(n_6923),
.B2(n_6791),
.Y(n_18124)
);

INVx1_ASAP7_75t_L g18125 ( 
.A(n_17856),
.Y(n_18125)
);

AOI22xp33_ASAP7_75t_L g18126 ( 
.A1(n_17729),
.A2(n_17814),
.B1(n_17869),
.B2(n_17851),
.Y(n_18126)
);

AOI22xp5_ASAP7_75t_L g18127 ( 
.A1(n_17925),
.A2(n_6892),
.B1(n_6928),
.B2(n_6923),
.Y(n_18127)
);

OAI32xp33_ASAP7_75t_L g18128 ( 
.A1(n_17885),
.A2(n_7110),
.A3(n_7132),
.B1(n_7106),
.B2(n_7057),
.Y(n_18128)
);

INVx1_ASAP7_75t_L g18129 ( 
.A(n_17775),
.Y(n_18129)
);

INVx1_ASAP7_75t_SL g18130 ( 
.A(n_17936),
.Y(n_18130)
);

NAND2xp5_ASAP7_75t_L g18131 ( 
.A(n_17759),
.B(n_8480),
.Y(n_18131)
);

AND2x2_ASAP7_75t_L g18132 ( 
.A(n_17747),
.B(n_8276),
.Y(n_18132)
);

NAND2xp5_ASAP7_75t_L g18133 ( 
.A(n_17884),
.B(n_8500),
.Y(n_18133)
);

OAI21xp33_ASAP7_75t_L g18134 ( 
.A1(n_17947),
.A2(n_7034),
.B(n_7015),
.Y(n_18134)
);

OAI22xp33_ASAP7_75t_L g18135 ( 
.A1(n_17831),
.A2(n_7225),
.B1(n_7254),
.B2(n_7199),
.Y(n_18135)
);

OAI32xp33_ASAP7_75t_L g18136 ( 
.A1(n_17890),
.A2(n_7110),
.A3(n_7132),
.B1(n_7106),
.B2(n_7057),
.Y(n_18136)
);

OAI21xp5_ASAP7_75t_SL g18137 ( 
.A1(n_17846),
.A2(n_7523),
.B(n_7081),
.Y(n_18137)
);

INVx2_ASAP7_75t_L g18138 ( 
.A(n_17888),
.Y(n_18138)
);

NAND2x1_ASAP7_75t_L g18139 ( 
.A(n_17837),
.B(n_17896),
.Y(n_18139)
);

AOI22xp5_ASAP7_75t_L g18140 ( 
.A1(n_17773),
.A2(n_6923),
.B1(n_6929),
.B2(n_6928),
.Y(n_18140)
);

NAND3xp33_ASAP7_75t_SL g18141 ( 
.A(n_17910),
.B(n_7425),
.C(n_7364),
.Y(n_18141)
);

INVx1_ASAP7_75t_L g18142 ( 
.A(n_17877),
.Y(n_18142)
);

AOI22xp33_ASAP7_75t_SL g18143 ( 
.A1(n_17735),
.A2(n_7669),
.B1(n_6706),
.B2(n_6929),
.Y(n_18143)
);

AOI22xp5_ASAP7_75t_L g18144 ( 
.A1(n_17805),
.A2(n_6928),
.B1(n_6975),
.B2(n_6929),
.Y(n_18144)
);

NAND2xp5_ASAP7_75t_L g18145 ( 
.A(n_17873),
.B(n_8500),
.Y(n_18145)
);

INVx1_ASAP7_75t_L g18146 ( 
.A(n_17913),
.Y(n_18146)
);

INVx1_ASAP7_75t_L g18147 ( 
.A(n_17914),
.Y(n_18147)
);

INVx1_ASAP7_75t_L g18148 ( 
.A(n_17848),
.Y(n_18148)
);

INVx2_ASAP7_75t_SL g18149 ( 
.A(n_17837),
.Y(n_18149)
);

NAND2xp5_ASAP7_75t_SL g18150 ( 
.A(n_17743),
.B(n_7199),
.Y(n_18150)
);

OAI221xp5_ASAP7_75t_L g18151 ( 
.A1(n_17842),
.A2(n_7301),
.B1(n_7570),
.B2(n_7244),
.C(n_7198),
.Y(n_18151)
);

OAI311xp33_ASAP7_75t_L g18152 ( 
.A1(n_17847),
.A2(n_6959),
.A3(n_6955),
.B1(n_6661),
.C1(n_7610),
.Y(n_18152)
);

NOR2xp67_ASAP7_75t_L g18153 ( 
.A(n_17926),
.B(n_17944),
.Y(n_18153)
);

AND2x2_ASAP7_75t_L g18154 ( 
.A(n_17870),
.B(n_8276),
.Y(n_18154)
);

INVx2_ASAP7_75t_L g18155 ( 
.A(n_17941),
.Y(n_18155)
);

AOI22xp33_ASAP7_75t_L g18156 ( 
.A1(n_17786),
.A2(n_8454),
.B1(n_8646),
.B2(n_8575),
.Y(n_18156)
);

AND2x4_ASAP7_75t_L g18157 ( 
.A(n_17928),
.B(n_8557),
.Y(n_18157)
);

OAI22xp33_ASAP7_75t_L g18158 ( 
.A1(n_17736),
.A2(n_7225),
.B1(n_7254),
.B2(n_7199),
.Y(n_18158)
);

OR2x2_ASAP7_75t_L g18159 ( 
.A(n_17876),
.B(n_8276),
.Y(n_18159)
);

NAND2xp5_ASAP7_75t_L g18160 ( 
.A(n_17899),
.B(n_8500),
.Y(n_18160)
);

INVx1_ASAP7_75t_L g18161 ( 
.A(n_17778),
.Y(n_18161)
);

INVx2_ASAP7_75t_SL g18162 ( 
.A(n_17852),
.Y(n_18162)
);

OAI21xp5_ASAP7_75t_SL g18163 ( 
.A1(n_17935),
.A2(n_7523),
.B(n_7081),
.Y(n_18163)
);

INVx1_ASAP7_75t_L g18164 ( 
.A(n_17778),
.Y(n_18164)
);

INVx1_ASAP7_75t_L g18165 ( 
.A(n_17778),
.Y(n_18165)
);

OAI21xp33_ASAP7_75t_L g18166 ( 
.A1(n_17840),
.A2(n_6929),
.B(n_6928),
.Y(n_18166)
);

NAND2xp5_ASAP7_75t_L g18167 ( 
.A(n_17907),
.B(n_8511),
.Y(n_18167)
);

NAND2xp5_ASAP7_75t_L g18168 ( 
.A(n_17881),
.B(n_8511),
.Y(n_18168)
);

AND2x2_ASAP7_75t_L g18169 ( 
.A(n_17751),
.B(n_8276),
.Y(n_18169)
);

INVx1_ASAP7_75t_L g18170 ( 
.A(n_17766),
.Y(n_18170)
);

NAND2xp5_ASAP7_75t_L g18171 ( 
.A(n_17809),
.B(n_8511),
.Y(n_18171)
);

INVx1_ASAP7_75t_L g18172 ( 
.A(n_17879),
.Y(n_18172)
);

NAND3xp33_ASAP7_75t_SL g18173 ( 
.A(n_17799),
.B(n_7425),
.C(n_7364),
.Y(n_18173)
);

AOI32xp33_ASAP7_75t_L g18174 ( 
.A1(n_17854),
.A2(n_8498),
.A3(n_8502),
.B1(n_8493),
.B2(n_8492),
.Y(n_18174)
);

AOI211xp5_ASAP7_75t_L g18175 ( 
.A1(n_17752),
.A2(n_7570),
.B(n_7198),
.C(n_8613),
.Y(n_18175)
);

INVxp67_ASAP7_75t_SL g18176 ( 
.A(n_17771),
.Y(n_18176)
);

INVxp67_ASAP7_75t_SL g18177 ( 
.A(n_17895),
.Y(n_18177)
);

OAI21xp33_ASAP7_75t_L g18178 ( 
.A1(n_17730),
.A2(n_6978),
.B(n_6975),
.Y(n_18178)
);

NAND2xp5_ASAP7_75t_L g18179 ( 
.A(n_17834),
.B(n_8548),
.Y(n_18179)
);

INVx1_ASAP7_75t_L g18180 ( 
.A(n_17808),
.Y(n_18180)
);

INVxp67_ASAP7_75t_SL g18181 ( 
.A(n_17779),
.Y(n_18181)
);

AND2x2_ASAP7_75t_L g18182 ( 
.A(n_17938),
.B(n_8276),
.Y(n_18182)
);

OAI221xp5_ASAP7_75t_L g18183 ( 
.A1(n_17836),
.A2(n_7570),
.B1(n_8922),
.B2(n_8931),
.C(n_8852),
.Y(n_18183)
);

AND2x2_ASAP7_75t_L g18184 ( 
.A(n_17843),
.B(n_8276),
.Y(n_18184)
);

NAND2xp33_ASAP7_75t_SL g18185 ( 
.A(n_17802),
.B(n_17818),
.Y(n_18185)
);

AOI22xp33_ASAP7_75t_L g18186 ( 
.A1(n_17930),
.A2(n_8454),
.B1(n_8646),
.B2(n_8575),
.Y(n_18186)
);

INVx1_ASAP7_75t_L g18187 ( 
.A(n_17924),
.Y(n_18187)
);

NOR2xp33_ASAP7_75t_L g18188 ( 
.A(n_17788),
.B(n_17886),
.Y(n_18188)
);

NAND3xp33_ASAP7_75t_SL g18189 ( 
.A(n_17919),
.B(n_7434),
.C(n_7364),
.Y(n_18189)
);

INVx1_ASAP7_75t_L g18190 ( 
.A(n_17937),
.Y(n_18190)
);

INVx2_ASAP7_75t_L g18191 ( 
.A(n_17933),
.Y(n_18191)
);

INVx2_ASAP7_75t_L g18192 ( 
.A(n_17908),
.Y(n_18192)
);

AOI221xp5_ASAP7_75t_L g18193 ( 
.A1(n_17889),
.A2(n_6978),
.B1(n_7070),
.B2(n_7058),
.C(n_6975),
.Y(n_18193)
);

INVx1_ASAP7_75t_L g18194 ( 
.A(n_18139),
.Y(n_18194)
);

NAND2xp5_ASAP7_75t_L g18195 ( 
.A(n_17954),
.B(n_17995),
.Y(n_18195)
);

NAND2xp5_ASAP7_75t_L g18196 ( 
.A(n_17957),
.B(n_17887),
.Y(n_18196)
);

INVx1_ASAP7_75t_L g18197 ( 
.A(n_18075),
.Y(n_18197)
);

NOR2xp33_ASAP7_75t_L g18198 ( 
.A(n_17952),
.B(n_17976),
.Y(n_18198)
);

NAND2xp5_ASAP7_75t_L g18199 ( 
.A(n_17961),
.B(n_17790),
.Y(n_18199)
);

INVx1_ASAP7_75t_L g18200 ( 
.A(n_17958),
.Y(n_18200)
);

INVx1_ASAP7_75t_L g18201 ( 
.A(n_17975),
.Y(n_18201)
);

INVx1_ASAP7_75t_L g18202 ( 
.A(n_17980),
.Y(n_18202)
);

NAND2xp5_ASAP7_75t_L g18203 ( 
.A(n_17977),
.B(n_17945),
.Y(n_18203)
);

NAND2x1p5_ASAP7_75t_L g18204 ( 
.A(n_17974),
.B(n_5180),
.Y(n_18204)
);

INVx1_ASAP7_75t_SL g18205 ( 
.A(n_18006),
.Y(n_18205)
);

NAND2xp5_ASAP7_75t_L g18206 ( 
.A(n_18004),
.B(n_17744),
.Y(n_18206)
);

OR2x2_ASAP7_75t_L g18207 ( 
.A(n_17981),
.B(n_17804),
.Y(n_18207)
);

AND2x2_ASAP7_75t_L g18208 ( 
.A(n_18052),
.B(n_17996),
.Y(n_18208)
);

INVx1_ASAP7_75t_L g18209 ( 
.A(n_18149),
.Y(n_18209)
);

INVx2_ASAP7_75t_SL g18210 ( 
.A(n_17999),
.Y(n_18210)
);

NAND2xp5_ASAP7_75t_L g18211 ( 
.A(n_17982),
.B(n_17894),
.Y(n_18211)
);

INVx1_ASAP7_75t_L g18212 ( 
.A(n_18021),
.Y(n_18212)
);

NAND2x1p5_ASAP7_75t_L g18213 ( 
.A(n_17971),
.B(n_5180),
.Y(n_18213)
);

NOR2xp33_ASAP7_75t_L g18214 ( 
.A(n_18051),
.B(n_17844),
.Y(n_18214)
);

INVx2_ASAP7_75t_L g18215 ( 
.A(n_18069),
.Y(n_18215)
);

INVx1_ASAP7_75t_L g18216 ( 
.A(n_18022),
.Y(n_18216)
);

AND2x2_ASAP7_75t_L g18217 ( 
.A(n_17986),
.B(n_8276),
.Y(n_18217)
);

NOR2xp33_ASAP7_75t_L g18218 ( 
.A(n_18015),
.B(n_6939),
.Y(n_18218)
);

INVx1_ASAP7_75t_L g18219 ( 
.A(n_18097),
.Y(n_18219)
);

INVx1_ASAP7_75t_L g18220 ( 
.A(n_18099),
.Y(n_18220)
);

NOR2xp33_ASAP7_75t_L g18221 ( 
.A(n_17979),
.B(n_6950),
.Y(n_18221)
);

INVx1_ASAP7_75t_L g18222 ( 
.A(n_18101),
.Y(n_18222)
);

AND2x2_ASAP7_75t_L g18223 ( 
.A(n_18020),
.B(n_8276),
.Y(n_18223)
);

INVx1_ASAP7_75t_L g18224 ( 
.A(n_18104),
.Y(n_18224)
);

AND2x2_ASAP7_75t_L g18225 ( 
.A(n_18003),
.B(n_8636),
.Y(n_18225)
);

NAND2xp5_ASAP7_75t_L g18226 ( 
.A(n_18034),
.B(n_8548),
.Y(n_18226)
);

BUFx2_ASAP7_75t_L g18227 ( 
.A(n_17973),
.Y(n_18227)
);

NOR2xp33_ASAP7_75t_L g18228 ( 
.A(n_18030),
.B(n_6950),
.Y(n_18228)
);

INVx1_ASAP7_75t_L g18229 ( 
.A(n_18032),
.Y(n_18229)
);

AND2x2_ASAP7_75t_L g18230 ( 
.A(n_18087),
.B(n_8636),
.Y(n_18230)
);

INVx1_ASAP7_75t_L g18231 ( 
.A(n_18109),
.Y(n_18231)
);

AND2x2_ASAP7_75t_L g18232 ( 
.A(n_18005),
.B(n_8636),
.Y(n_18232)
);

NOR2xp33_ASAP7_75t_L g18233 ( 
.A(n_18064),
.B(n_6950),
.Y(n_18233)
);

NAND2xp5_ASAP7_75t_L g18234 ( 
.A(n_17953),
.B(n_8548),
.Y(n_18234)
);

INVx1_ASAP7_75t_L g18235 ( 
.A(n_17955),
.Y(n_18235)
);

NAND2xp5_ASAP7_75t_L g18236 ( 
.A(n_18046),
.B(n_8555),
.Y(n_18236)
);

AOI31xp33_ASAP7_75t_L g18237 ( 
.A1(n_18036),
.A2(n_5465),
.A3(n_5490),
.B(n_5350),
.Y(n_18237)
);

AND2x2_ASAP7_75t_L g18238 ( 
.A(n_17994),
.B(n_8636),
.Y(n_18238)
);

INVx1_ASAP7_75t_L g18239 ( 
.A(n_18056),
.Y(n_18239)
);

INVx2_ASAP7_75t_L g18240 ( 
.A(n_17990),
.Y(n_18240)
);

NOR2xp33_ASAP7_75t_L g18241 ( 
.A(n_18016),
.B(n_6967),
.Y(n_18241)
);

OAI22xp5_ASAP7_75t_L g18242 ( 
.A1(n_18012),
.A2(n_6975),
.B1(n_7058),
.B2(n_6978),
.Y(n_18242)
);

NAND2xp5_ASAP7_75t_L g18243 ( 
.A(n_18096),
.B(n_8555),
.Y(n_18243)
);

NOR2x1_ASAP7_75t_L g18244 ( 
.A(n_18092),
.B(n_8454),
.Y(n_18244)
);

NAND2xp5_ASAP7_75t_L g18245 ( 
.A(n_18148),
.B(n_8555),
.Y(n_18245)
);

NAND2xp5_ASAP7_75t_L g18246 ( 
.A(n_18040),
.B(n_8577),
.Y(n_18246)
);

INVx1_ASAP7_75t_L g18247 ( 
.A(n_17956),
.Y(n_18247)
);

AND2x2_ASAP7_75t_L g18248 ( 
.A(n_18039),
.B(n_8636),
.Y(n_18248)
);

NAND2xp5_ASAP7_75t_L g18249 ( 
.A(n_18024),
.B(n_8577),
.Y(n_18249)
);

INVx1_ASAP7_75t_L g18250 ( 
.A(n_18190),
.Y(n_18250)
);

NAND2xp5_ASAP7_75t_L g18251 ( 
.A(n_18084),
.B(n_8577),
.Y(n_18251)
);

INVx1_ASAP7_75t_L g18252 ( 
.A(n_17998),
.Y(n_18252)
);

INVx1_ASAP7_75t_L g18253 ( 
.A(n_18072),
.Y(n_18253)
);

INVx1_ASAP7_75t_L g18254 ( 
.A(n_18077),
.Y(n_18254)
);

INVx1_ASAP7_75t_L g18255 ( 
.A(n_18142),
.Y(n_18255)
);

NAND2xp5_ASAP7_75t_L g18256 ( 
.A(n_18162),
.B(n_8582),
.Y(n_18256)
);

NAND2xp5_ASAP7_75t_L g18257 ( 
.A(n_18095),
.B(n_8582),
.Y(n_18257)
);

AND2x2_ASAP7_75t_L g18258 ( 
.A(n_18067),
.B(n_8636),
.Y(n_18258)
);

NAND2xp5_ASAP7_75t_L g18259 ( 
.A(n_18138),
.B(n_8582),
.Y(n_18259)
);

HB1xp67_ASAP7_75t_L g18260 ( 
.A(n_18153),
.Y(n_18260)
);

AND2x2_ASAP7_75t_L g18261 ( 
.A(n_18008),
.B(n_8636),
.Y(n_18261)
);

AND2x2_ASAP7_75t_L g18262 ( 
.A(n_17991),
.B(n_8636),
.Y(n_18262)
);

OAI22xp5_ASAP7_75t_L g18263 ( 
.A1(n_17950),
.A2(n_6978),
.B1(n_7070),
.B2(n_7058),
.Y(n_18263)
);

NOR2xp33_ASAP7_75t_L g18264 ( 
.A(n_18130),
.B(n_6967),
.Y(n_18264)
);

AND2x2_ASAP7_75t_L g18265 ( 
.A(n_17970),
.B(n_8557),
.Y(n_18265)
);

INVx1_ASAP7_75t_L g18266 ( 
.A(n_18161),
.Y(n_18266)
);

AND2x2_ASAP7_75t_L g18267 ( 
.A(n_17987),
.B(n_8561),
.Y(n_18267)
);

AOI22xp33_ASAP7_75t_L g18268 ( 
.A1(n_18007),
.A2(n_8646),
.B1(n_8575),
.B2(n_7058),
.Y(n_18268)
);

INVx1_ASAP7_75t_L g18269 ( 
.A(n_18164),
.Y(n_18269)
);

INVx2_ASAP7_75t_L g18270 ( 
.A(n_18019),
.Y(n_18270)
);

INVx1_ASAP7_75t_L g18271 ( 
.A(n_18165),
.Y(n_18271)
);

NAND2xp5_ASAP7_75t_L g18272 ( 
.A(n_18079),
.B(n_8589),
.Y(n_18272)
);

NAND2xp5_ASAP7_75t_L g18273 ( 
.A(n_17963),
.B(n_8589),
.Y(n_18273)
);

INVx1_ASAP7_75t_L g18274 ( 
.A(n_18176),
.Y(n_18274)
);

INVx1_ASAP7_75t_SL g18275 ( 
.A(n_18185),
.Y(n_18275)
);

AND2x2_ASAP7_75t_L g18276 ( 
.A(n_18102),
.B(n_8561),
.Y(n_18276)
);

INVx1_ASAP7_75t_L g18277 ( 
.A(n_18187),
.Y(n_18277)
);

NAND2xp5_ASAP7_75t_L g18278 ( 
.A(n_18181),
.B(n_8589),
.Y(n_18278)
);

NAND2xp5_ASAP7_75t_L g18279 ( 
.A(n_18172),
.B(n_18188),
.Y(n_18279)
);

NAND2xp5_ASAP7_75t_L g18280 ( 
.A(n_18080),
.B(n_8602),
.Y(n_18280)
);

INVx1_ASAP7_75t_L g18281 ( 
.A(n_18028),
.Y(n_18281)
);

INVx1_ASAP7_75t_L g18282 ( 
.A(n_18023),
.Y(n_18282)
);

INVx1_ASAP7_75t_L g18283 ( 
.A(n_18002),
.Y(n_18283)
);

OR2x2_ASAP7_75t_L g18284 ( 
.A(n_18173),
.B(n_8097),
.Y(n_18284)
);

INVx1_ASAP7_75t_L g18285 ( 
.A(n_18073),
.Y(n_18285)
);

INVxp67_ASAP7_75t_L g18286 ( 
.A(n_18112),
.Y(n_18286)
);

INVx1_ASAP7_75t_SL g18287 ( 
.A(n_17967),
.Y(n_18287)
);

INVx1_ASAP7_75t_L g18288 ( 
.A(n_18170),
.Y(n_18288)
);

OR2x2_ASAP7_75t_L g18289 ( 
.A(n_17969),
.B(n_8097),
.Y(n_18289)
);

NAND2xp5_ASAP7_75t_L g18290 ( 
.A(n_17951),
.B(n_8602),
.Y(n_18290)
);

NAND2xp5_ASAP7_75t_L g18291 ( 
.A(n_18035),
.B(n_8602),
.Y(n_18291)
);

NOR2xp33_ASAP7_75t_L g18292 ( 
.A(n_18106),
.B(n_18116),
.Y(n_18292)
);

INVx1_ASAP7_75t_L g18293 ( 
.A(n_18177),
.Y(n_18293)
);

NAND2xp5_ASAP7_75t_SL g18294 ( 
.A(n_17966),
.B(n_7199),
.Y(n_18294)
);

NAND2xp5_ASAP7_75t_L g18295 ( 
.A(n_18044),
.B(n_8607),
.Y(n_18295)
);

NAND2xp5_ASAP7_75t_L g18296 ( 
.A(n_18155),
.B(n_18125),
.Y(n_18296)
);

NOR2xp33_ASAP7_75t_L g18297 ( 
.A(n_18180),
.B(n_6967),
.Y(n_18297)
);

INVx1_ASAP7_75t_L g18298 ( 
.A(n_18033),
.Y(n_18298)
);

INVx1_ASAP7_75t_L g18299 ( 
.A(n_18129),
.Y(n_18299)
);

INVx1_ASAP7_75t_L g18300 ( 
.A(n_18082),
.Y(n_18300)
);

AND2x2_ASAP7_75t_L g18301 ( 
.A(n_18085),
.B(n_8561),
.Y(n_18301)
);

INVx1_ASAP7_75t_L g18302 ( 
.A(n_18083),
.Y(n_18302)
);

INVx1_ASAP7_75t_L g18303 ( 
.A(n_18089),
.Y(n_18303)
);

NAND2xp5_ASAP7_75t_L g18304 ( 
.A(n_18094),
.B(n_18088),
.Y(n_18304)
);

AOI22xp5_ASAP7_75t_L g18305 ( 
.A1(n_17992),
.A2(n_7070),
.B1(n_7107),
.B2(n_7104),
.Y(n_18305)
);

AND2x2_ASAP7_75t_L g18306 ( 
.A(n_18054),
.B(n_18126),
.Y(n_18306)
);

NAND2xp5_ASAP7_75t_L g18307 ( 
.A(n_17993),
.B(n_8607),
.Y(n_18307)
);

OAI22xp5_ASAP7_75t_L g18308 ( 
.A1(n_18183),
.A2(n_7104),
.B1(n_7107),
.B2(n_7070),
.Y(n_18308)
);

INVx2_ASAP7_75t_L g18309 ( 
.A(n_18157),
.Y(n_18309)
);

NOR2xp33_ASAP7_75t_L g18310 ( 
.A(n_18076),
.B(n_6967),
.Y(n_18310)
);

NAND2xp5_ASAP7_75t_L g18311 ( 
.A(n_18191),
.B(n_18192),
.Y(n_18311)
);

INVx1_ASAP7_75t_SL g18312 ( 
.A(n_18053),
.Y(n_18312)
);

NAND2xp5_ASAP7_75t_L g18313 ( 
.A(n_17965),
.B(n_8607),
.Y(n_18313)
);

INVx1_ASAP7_75t_SL g18314 ( 
.A(n_17960),
.Y(n_18314)
);

INVx1_ASAP7_75t_L g18315 ( 
.A(n_18146),
.Y(n_18315)
);

NAND2xp5_ASAP7_75t_L g18316 ( 
.A(n_18154),
.B(n_8623),
.Y(n_18316)
);

OR2x2_ASAP7_75t_L g18317 ( 
.A(n_18070),
.B(n_8097),
.Y(n_18317)
);

NAND2xp5_ASAP7_75t_L g18318 ( 
.A(n_18147),
.B(n_8623),
.Y(n_18318)
);

INVx2_ASAP7_75t_SL g18319 ( 
.A(n_18150),
.Y(n_18319)
);

NOR2xp33_ASAP7_75t_L g18320 ( 
.A(n_18141),
.B(n_6967),
.Y(n_18320)
);

AOI22xp33_ASAP7_75t_L g18321 ( 
.A1(n_18063),
.A2(n_18050),
.B1(n_18184),
.B2(n_17962),
.Y(n_18321)
);

AND2x2_ASAP7_75t_L g18322 ( 
.A(n_18107),
.B(n_8566),
.Y(n_18322)
);

NAND2xp5_ASAP7_75t_L g18323 ( 
.A(n_18159),
.B(n_8623),
.Y(n_18323)
);

NAND2xp5_ASAP7_75t_L g18324 ( 
.A(n_18121),
.B(n_8647),
.Y(n_18324)
);

INVxp67_ASAP7_75t_SL g18325 ( 
.A(n_17988),
.Y(n_18325)
);

NAND2xp5_ASAP7_75t_L g18326 ( 
.A(n_18123),
.B(n_8647),
.Y(n_18326)
);

INVx1_ASAP7_75t_L g18327 ( 
.A(n_18145),
.Y(n_18327)
);

NAND2xp5_ASAP7_75t_L g18328 ( 
.A(n_18132),
.B(n_8647),
.Y(n_18328)
);

INVx1_ASAP7_75t_SL g18329 ( 
.A(n_18060),
.Y(n_18329)
);

AND2x2_ASAP7_75t_SL g18330 ( 
.A(n_18010),
.B(n_5470),
.Y(n_18330)
);

INVx1_ASAP7_75t_L g18331 ( 
.A(n_18029),
.Y(n_18331)
);

BUFx2_ASAP7_75t_L g18332 ( 
.A(n_18045),
.Y(n_18332)
);

NOR2xp33_ASAP7_75t_L g18333 ( 
.A(n_18090),
.B(n_6967),
.Y(n_18333)
);

NAND2xp5_ASAP7_75t_L g18334 ( 
.A(n_18143),
.B(n_8651),
.Y(n_18334)
);

NAND2xp5_ASAP7_75t_L g18335 ( 
.A(n_18137),
.B(n_8651),
.Y(n_18335)
);

INVx1_ASAP7_75t_SL g18336 ( 
.A(n_18055),
.Y(n_18336)
);

INVx1_ASAP7_75t_SL g18337 ( 
.A(n_18065),
.Y(n_18337)
);

INVx1_ASAP7_75t_L g18338 ( 
.A(n_18066),
.Y(n_18338)
);

INVx1_ASAP7_75t_L g18339 ( 
.A(n_18108),
.Y(n_18339)
);

NAND2xp5_ASAP7_75t_L g18340 ( 
.A(n_18133),
.B(n_8651),
.Y(n_18340)
);

INVx1_ASAP7_75t_L g18341 ( 
.A(n_18131),
.Y(n_18341)
);

AO22x2_ASAP7_75t_L g18342 ( 
.A1(n_18189),
.A2(n_8668),
.B1(n_8672),
.B2(n_8656),
.Y(n_18342)
);

OAI221xp5_ASAP7_75t_L g18343 ( 
.A1(n_18171),
.A2(n_8931),
.B1(n_8922),
.B2(n_8852),
.C(n_7109),
.Y(n_18343)
);

INVx1_ASAP7_75t_L g18344 ( 
.A(n_18160),
.Y(n_18344)
);

HB1xp67_ASAP7_75t_L g18345 ( 
.A(n_17989),
.Y(n_18345)
);

AND2x2_ASAP7_75t_L g18346 ( 
.A(n_18182),
.B(n_8566),
.Y(n_18346)
);

NAND2xp5_ASAP7_75t_L g18347 ( 
.A(n_18134),
.B(n_8656),
.Y(n_18347)
);

AND2x2_ASAP7_75t_L g18348 ( 
.A(n_18169),
.B(n_8566),
.Y(n_18348)
);

NAND2xp5_ASAP7_75t_L g18349 ( 
.A(n_18163),
.B(n_8656),
.Y(n_18349)
);

NAND2xp5_ASAP7_75t_L g18350 ( 
.A(n_18093),
.B(n_18026),
.Y(n_18350)
);

OR2x2_ASAP7_75t_L g18351 ( 
.A(n_18078),
.B(n_8097),
.Y(n_18351)
);

NAND2xp5_ASAP7_75t_L g18352 ( 
.A(n_18167),
.B(n_8668),
.Y(n_18352)
);

NAND2xp5_ASAP7_75t_L g18353 ( 
.A(n_18114),
.B(n_8668),
.Y(n_18353)
);

INVx1_ASAP7_75t_L g18354 ( 
.A(n_18086),
.Y(n_18354)
);

INVx1_ASAP7_75t_L g18355 ( 
.A(n_18091),
.Y(n_18355)
);

NAND2xp5_ASAP7_75t_L g18356 ( 
.A(n_18058),
.B(n_8672),
.Y(n_18356)
);

NAND2xp5_ASAP7_75t_L g18357 ( 
.A(n_18124),
.B(n_8672),
.Y(n_18357)
);

INVx1_ASAP7_75t_SL g18358 ( 
.A(n_18168),
.Y(n_18358)
);

HB1xp67_ASAP7_75t_L g18359 ( 
.A(n_18157),
.Y(n_18359)
);

AND2x2_ASAP7_75t_L g18360 ( 
.A(n_18115),
.B(n_8336),
.Y(n_18360)
);

AND2x2_ASAP7_75t_L g18361 ( 
.A(n_18140),
.B(n_8336),
.Y(n_18361)
);

NAND2xp5_ASAP7_75t_L g18362 ( 
.A(n_18179),
.B(n_8675),
.Y(n_18362)
);

HB1xp67_ASAP7_75t_L g18363 ( 
.A(n_18098),
.Y(n_18363)
);

INVx1_ASAP7_75t_L g18364 ( 
.A(n_18062),
.Y(n_18364)
);

OR2x2_ASAP7_75t_L g18365 ( 
.A(n_17997),
.B(n_8097),
.Y(n_18365)
);

INVx1_ASAP7_75t_L g18366 ( 
.A(n_18110),
.Y(n_18366)
);

INVx1_ASAP7_75t_L g18367 ( 
.A(n_18118),
.Y(n_18367)
);

NAND2xp5_ASAP7_75t_L g18368 ( 
.A(n_18103),
.B(n_8675),
.Y(n_18368)
);

INVx1_ASAP7_75t_L g18369 ( 
.A(n_18120),
.Y(n_18369)
);

AND2x2_ASAP7_75t_L g18370 ( 
.A(n_18105),
.B(n_8336),
.Y(n_18370)
);

AND2x2_ASAP7_75t_L g18371 ( 
.A(n_17959),
.B(n_8336),
.Y(n_18371)
);

NAND2xp5_ASAP7_75t_L g18372 ( 
.A(n_18175),
.B(n_8675),
.Y(n_18372)
);

INVx2_ASAP7_75t_SL g18373 ( 
.A(n_18014),
.Y(n_18373)
);

NOR2xp33_ASAP7_75t_L g18374 ( 
.A(n_18151),
.B(n_7007),
.Y(n_18374)
);

NOR2xp33_ASAP7_75t_L g18375 ( 
.A(n_18111),
.B(n_18031),
.Y(n_18375)
);

INVx1_ASAP7_75t_L g18376 ( 
.A(n_18128),
.Y(n_18376)
);

INVx2_ASAP7_75t_L g18377 ( 
.A(n_18014),
.Y(n_18377)
);

CKINVDCx16_ASAP7_75t_R g18378 ( 
.A(n_17984),
.Y(n_18378)
);

AND2x2_ASAP7_75t_L g18379 ( 
.A(n_18127),
.B(n_8336),
.Y(n_18379)
);

NAND2xp5_ASAP7_75t_L g18380 ( 
.A(n_18174),
.B(n_8683),
.Y(n_18380)
);

AOI22xp5_ASAP7_75t_L g18381 ( 
.A1(n_18166),
.A2(n_18178),
.B1(n_18158),
.B2(n_17985),
.Y(n_18381)
);

OR2x6_ASAP7_75t_L g18382 ( 
.A(n_18027),
.B(n_5498),
.Y(n_18382)
);

INVx1_ASAP7_75t_SL g18383 ( 
.A(n_18042),
.Y(n_18383)
);

NOR2xp33_ASAP7_75t_L g18384 ( 
.A(n_17978),
.B(n_7007),
.Y(n_18384)
);

AND2x4_ASAP7_75t_L g18385 ( 
.A(n_18057),
.B(n_8204),
.Y(n_18385)
);

NAND2xp5_ASAP7_75t_L g18386 ( 
.A(n_18037),
.B(n_8683),
.Y(n_18386)
);

INVx1_ASAP7_75t_L g18387 ( 
.A(n_18136),
.Y(n_18387)
);

INVx1_ASAP7_75t_L g18388 ( 
.A(n_18038),
.Y(n_18388)
);

NAND2xp5_ASAP7_75t_L g18389 ( 
.A(n_18193),
.B(n_8683),
.Y(n_18389)
);

INVx1_ASAP7_75t_L g18390 ( 
.A(n_18048),
.Y(n_18390)
);

NAND2xp5_ASAP7_75t_L g18391 ( 
.A(n_18135),
.B(n_8704),
.Y(n_18391)
);

NOR2x1_ASAP7_75t_L g18392 ( 
.A(n_18009),
.B(n_8454),
.Y(n_18392)
);

AND2x2_ASAP7_75t_L g18393 ( 
.A(n_18156),
.B(n_8336),
.Y(n_18393)
);

OAI21xp5_ASAP7_75t_L g18394 ( 
.A1(n_18152),
.A2(n_7724),
.B(n_7706),
.Y(n_18394)
);

INVx1_ASAP7_75t_L g18395 ( 
.A(n_18043),
.Y(n_18395)
);

NAND2xp5_ASAP7_75t_L g18396 ( 
.A(n_18186),
.B(n_8704),
.Y(n_18396)
);

INVx1_ASAP7_75t_L g18397 ( 
.A(n_18068),
.Y(n_18397)
);

INVx1_ASAP7_75t_L g18398 ( 
.A(n_18047),
.Y(n_18398)
);

NAND2xp5_ASAP7_75t_L g18399 ( 
.A(n_18119),
.B(n_8704),
.Y(n_18399)
);

INVx1_ASAP7_75t_L g18400 ( 
.A(n_17972),
.Y(n_18400)
);

NOR2x1_ASAP7_75t_L g18401 ( 
.A(n_18011),
.B(n_8206),
.Y(n_18401)
);

NAND2xp5_ASAP7_75t_SL g18402 ( 
.A(n_17983),
.B(n_7199),
.Y(n_18402)
);

NAND2xp5_ASAP7_75t_L g18403 ( 
.A(n_18061),
.B(n_8718),
.Y(n_18403)
);

NAND2xp5_ASAP7_75t_L g18404 ( 
.A(n_18025),
.B(n_8718),
.Y(n_18404)
);

AND2x2_ASAP7_75t_L g18405 ( 
.A(n_18074),
.B(n_8336),
.Y(n_18405)
);

INVx1_ASAP7_75t_L g18406 ( 
.A(n_17972),
.Y(n_18406)
);

NAND2xp5_ASAP7_75t_L g18407 ( 
.A(n_18059),
.B(n_8718),
.Y(n_18407)
);

INVx1_ASAP7_75t_L g18408 ( 
.A(n_18018),
.Y(n_18408)
);

NAND2xp5_ASAP7_75t_L g18409 ( 
.A(n_18001),
.B(n_8733),
.Y(n_18409)
);

OR2x2_ASAP7_75t_L g18410 ( 
.A(n_18100),
.B(n_17964),
.Y(n_18410)
);

NOR2x1_ASAP7_75t_L g18411 ( 
.A(n_18018),
.B(n_8206),
.Y(n_18411)
);

INVxp67_ASAP7_75t_L g18412 ( 
.A(n_18113),
.Y(n_18412)
);

OR2x2_ASAP7_75t_L g18413 ( 
.A(n_18144),
.B(n_17968),
.Y(n_18413)
);

INVx2_ASAP7_75t_L g18414 ( 
.A(n_18117),
.Y(n_18414)
);

INVx1_ASAP7_75t_L g18415 ( 
.A(n_18117),
.Y(n_18415)
);

AND2x2_ASAP7_75t_L g18416 ( 
.A(n_18017),
.B(n_8535),
.Y(n_18416)
);

HB1xp67_ASAP7_75t_L g18417 ( 
.A(n_18013),
.Y(n_18417)
);

NAND2x1_ASAP7_75t_L g18418 ( 
.A(n_18122),
.B(n_9947),
.Y(n_18418)
);

NAND2xp5_ASAP7_75t_L g18419 ( 
.A(n_18000),
.B(n_8733),
.Y(n_18419)
);

INVx1_ASAP7_75t_L g18420 ( 
.A(n_18041),
.Y(n_18420)
);

OR2x2_ASAP7_75t_L g18421 ( 
.A(n_18071),
.B(n_8097),
.Y(n_18421)
);

NAND2xp5_ASAP7_75t_SL g18422 ( 
.A(n_18049),
.B(n_7199),
.Y(n_18422)
);

INVx1_ASAP7_75t_L g18423 ( 
.A(n_18081),
.Y(n_18423)
);

NOR2xp33_ASAP7_75t_L g18424 ( 
.A(n_17995),
.B(n_7007),
.Y(n_18424)
);

AOI222xp33_ASAP7_75t_SL g18425 ( 
.A1(n_17957),
.A2(n_7124),
.B1(n_7524),
.B2(n_7588),
.C1(n_7548),
.C2(n_7451),
.Y(n_18425)
);

AND2x2_ASAP7_75t_L g18426 ( 
.A(n_17995),
.B(n_8535),
.Y(n_18426)
);

NAND2xp5_ASAP7_75t_L g18427 ( 
.A(n_17954),
.B(n_8733),
.Y(n_18427)
);

NAND2xp5_ASAP7_75t_L g18428 ( 
.A(n_17954),
.B(n_8773),
.Y(n_18428)
);

NAND2xp5_ASAP7_75t_L g18429 ( 
.A(n_17954),
.B(n_8773),
.Y(n_18429)
);

NAND2xp5_ASAP7_75t_SL g18430 ( 
.A(n_17954),
.B(n_7199),
.Y(n_18430)
);

INVx1_ASAP7_75t_L g18431 ( 
.A(n_18139),
.Y(n_18431)
);

INVx1_ASAP7_75t_L g18432 ( 
.A(n_18139),
.Y(n_18432)
);

NOR2xp33_ASAP7_75t_L g18433 ( 
.A(n_17995),
.B(n_7007),
.Y(n_18433)
);

INVx1_ASAP7_75t_L g18434 ( 
.A(n_18139),
.Y(n_18434)
);

INVx1_ASAP7_75t_L g18435 ( 
.A(n_18139),
.Y(n_18435)
);

NAND2xp5_ASAP7_75t_L g18436 ( 
.A(n_17954),
.B(n_8773),
.Y(n_18436)
);

INVx1_ASAP7_75t_L g18437 ( 
.A(n_18139),
.Y(n_18437)
);

INVx3_ASAP7_75t_SL g18438 ( 
.A(n_17974),
.Y(n_18438)
);

NOR2xp33_ASAP7_75t_L g18439 ( 
.A(n_17995),
.B(n_7007),
.Y(n_18439)
);

NAND2xp5_ASAP7_75t_L g18440 ( 
.A(n_17954),
.B(n_8780),
.Y(n_18440)
);

NOR2x1p5_ASAP7_75t_L g18441 ( 
.A(n_18195),
.B(n_5453),
.Y(n_18441)
);

AND2x2_ASAP7_75t_L g18442 ( 
.A(n_18208),
.B(n_8535),
.Y(n_18442)
);

OR2x2_ASAP7_75t_L g18443 ( 
.A(n_18275),
.B(n_8097),
.Y(n_18443)
);

AOI22xp5_ASAP7_75t_L g18444 ( 
.A1(n_18205),
.A2(n_7104),
.B1(n_7109),
.B2(n_7107),
.Y(n_18444)
);

INVx1_ASAP7_75t_SL g18445 ( 
.A(n_18438),
.Y(n_18445)
);

AND2x2_ASAP7_75t_L g18446 ( 
.A(n_18222),
.B(n_8535),
.Y(n_18446)
);

AND2x2_ASAP7_75t_L g18447 ( 
.A(n_18224),
.B(n_8535),
.Y(n_18447)
);

AOI221xp5_ASAP7_75t_SL g18448 ( 
.A1(n_18247),
.A2(n_7656),
.B1(n_7611),
.B2(n_7124),
.C(n_6670),
.Y(n_18448)
);

INVx1_ASAP7_75t_L g18449 ( 
.A(n_18359),
.Y(n_18449)
);

INVxp67_ASAP7_75t_L g18450 ( 
.A(n_18198),
.Y(n_18450)
);

INVx1_ASAP7_75t_L g18451 ( 
.A(n_18194),
.Y(n_18451)
);

INVx1_ASAP7_75t_L g18452 ( 
.A(n_18431),
.Y(n_18452)
);

NOR3xp33_ASAP7_75t_L g18453 ( 
.A(n_18212),
.B(n_5287),
.C(n_5197),
.Y(n_18453)
);

INVx2_ASAP7_75t_L g18454 ( 
.A(n_18309),
.Y(n_18454)
);

NAND2x1_ASAP7_75t_L g18455 ( 
.A(n_18432),
.B(n_4865),
.Y(n_18455)
);

NAND2xp5_ASAP7_75t_L g18456 ( 
.A(n_18266),
.B(n_18269),
.Y(n_18456)
);

NOR4xp25_ASAP7_75t_SL g18457 ( 
.A(n_18434),
.B(n_6906),
.C(n_7004),
.D(n_7000),
.Y(n_18457)
);

INVx1_ASAP7_75t_L g18458 ( 
.A(n_18435),
.Y(n_18458)
);

INVx1_ASAP7_75t_L g18459 ( 
.A(n_18437),
.Y(n_18459)
);

OR2x2_ASAP7_75t_L g18460 ( 
.A(n_18231),
.B(n_8097),
.Y(n_18460)
);

INVx1_ASAP7_75t_L g18461 ( 
.A(n_18251),
.Y(n_18461)
);

INVx2_ASAP7_75t_L g18462 ( 
.A(n_18210),
.Y(n_18462)
);

AND2x2_ASAP7_75t_L g18463 ( 
.A(n_18239),
.B(n_8535),
.Y(n_18463)
);

NAND2xp5_ASAP7_75t_L g18464 ( 
.A(n_18271),
.B(n_8780),
.Y(n_18464)
);

OR2x2_ASAP7_75t_L g18465 ( 
.A(n_18219),
.B(n_7707),
.Y(n_18465)
);

OR2x2_ASAP7_75t_L g18466 ( 
.A(n_18220),
.B(n_7707),
.Y(n_18466)
);

INVxp67_ASAP7_75t_L g18467 ( 
.A(n_18260),
.Y(n_18467)
);

INVx1_ASAP7_75t_L g18468 ( 
.A(n_18209),
.Y(n_18468)
);

OAI21xp33_ASAP7_75t_L g18469 ( 
.A1(n_18279),
.A2(n_7107),
.B(n_7104),
.Y(n_18469)
);

INVxp67_ASAP7_75t_L g18470 ( 
.A(n_18292),
.Y(n_18470)
);

INVx1_ASAP7_75t_L g18471 ( 
.A(n_18229),
.Y(n_18471)
);

INVx1_ASAP7_75t_SL g18472 ( 
.A(n_18306),
.Y(n_18472)
);

NAND2xp5_ASAP7_75t_L g18473 ( 
.A(n_18255),
.B(n_8780),
.Y(n_18473)
);

OAI22xp5_ASAP7_75t_L g18474 ( 
.A1(n_18215),
.A2(n_7118),
.B1(n_7187),
.B2(n_7109),
.Y(n_18474)
);

INVxp33_ASAP7_75t_L g18475 ( 
.A(n_18424),
.Y(n_18475)
);

INVx1_ASAP7_75t_SL g18476 ( 
.A(n_18216),
.Y(n_18476)
);

INVx3_ASAP7_75t_SL g18477 ( 
.A(n_18253),
.Y(n_18477)
);

NOR3xp33_ASAP7_75t_L g18478 ( 
.A(n_18197),
.B(n_5363),
.C(n_5287),
.Y(n_18478)
);

INVx1_ASAP7_75t_SL g18479 ( 
.A(n_18246),
.Y(n_18479)
);

NOR2xp33_ASAP7_75t_L g18480 ( 
.A(n_18286),
.B(n_6706),
.Y(n_18480)
);

INVx3_ASAP7_75t_SL g18481 ( 
.A(n_18254),
.Y(n_18481)
);

AND2x2_ASAP7_75t_L g18482 ( 
.A(n_18201),
.B(n_8535),
.Y(n_18482)
);

AND2x2_ASAP7_75t_L g18483 ( 
.A(n_18202),
.B(n_6623),
.Y(n_18483)
);

INVx1_ASAP7_75t_L g18484 ( 
.A(n_18433),
.Y(n_18484)
);

AND3x2_ASAP7_75t_L g18485 ( 
.A(n_18400),
.B(n_5492),
.C(n_7207),
.Y(n_18485)
);

INVx1_ASAP7_75t_L g18486 ( 
.A(n_18439),
.Y(n_18486)
);

AND2x2_ASAP7_75t_L g18487 ( 
.A(n_18228),
.B(n_6623),
.Y(n_18487)
);

NAND2x1_ASAP7_75t_L g18488 ( 
.A(n_18285),
.B(n_4865),
.Y(n_18488)
);

INVx1_ASAP7_75t_L g18489 ( 
.A(n_18282),
.Y(n_18489)
);

AND2x2_ASAP7_75t_L g18490 ( 
.A(n_18233),
.B(n_18218),
.Y(n_18490)
);

INVx1_ASAP7_75t_SL g18491 ( 
.A(n_18312),
.Y(n_18491)
);

INVx1_ASAP7_75t_L g18492 ( 
.A(n_18415),
.Y(n_18492)
);

INVx2_ASAP7_75t_L g18493 ( 
.A(n_18204),
.Y(n_18493)
);

OAI22xp5_ASAP7_75t_L g18494 ( 
.A1(n_18321),
.A2(n_18284),
.B1(n_18268),
.B2(n_18412),
.Y(n_18494)
);

INVxp67_ASAP7_75t_L g18495 ( 
.A(n_18199),
.Y(n_18495)
);

NAND2xp5_ASAP7_75t_L g18496 ( 
.A(n_18200),
.B(n_8799),
.Y(n_18496)
);

INVx2_ASAP7_75t_L g18497 ( 
.A(n_18213),
.Y(n_18497)
);

NAND2xp33_ASAP7_75t_R g18498 ( 
.A(n_18227),
.B(n_5228),
.Y(n_18498)
);

OR2x2_ASAP7_75t_L g18499 ( 
.A(n_18290),
.B(n_18250),
.Y(n_18499)
);

INVx2_ASAP7_75t_L g18500 ( 
.A(n_18426),
.Y(n_18500)
);

INVx1_ASAP7_75t_L g18501 ( 
.A(n_18414),
.Y(n_18501)
);

NAND2xp5_ASAP7_75t_L g18502 ( 
.A(n_18297),
.B(n_8799),
.Y(n_18502)
);

NOR2xp33_ASAP7_75t_R g18503 ( 
.A(n_18235),
.B(n_5834),
.Y(n_18503)
);

XNOR2xp5_ASAP7_75t_L g18504 ( 
.A(n_18381),
.B(n_8852),
.Y(n_18504)
);

INVx1_ASAP7_75t_L g18505 ( 
.A(n_18245),
.Y(n_18505)
);

INVx2_ASAP7_75t_SL g18506 ( 
.A(n_18410),
.Y(n_18506)
);

XOR2x2_ASAP7_75t_L g18507 ( 
.A(n_18196),
.B(n_5513),
.Y(n_18507)
);

NOR2xp33_ASAP7_75t_L g18508 ( 
.A(n_18378),
.B(n_6706),
.Y(n_18508)
);

NAND2xp5_ASAP7_75t_L g18509 ( 
.A(n_18264),
.B(n_8799),
.Y(n_18509)
);

OAI21xp33_ASAP7_75t_SL g18510 ( 
.A1(n_18324),
.A2(n_8498),
.B(n_8493),
.Y(n_18510)
);

CKINVDCx5p33_ASAP7_75t_R g18511 ( 
.A(n_18252),
.Y(n_18511)
);

INVx1_ASAP7_75t_SL g18512 ( 
.A(n_18287),
.Y(n_18512)
);

INVx3_ASAP7_75t_L g18513 ( 
.A(n_18240),
.Y(n_18513)
);

AOI21xp33_ASAP7_75t_SL g18514 ( 
.A1(n_18288),
.A2(n_7847),
.B(n_7842),
.Y(n_18514)
);

NOR3xp33_ASAP7_75t_SL g18515 ( 
.A(n_18311),
.B(n_7522),
.C(n_7491),
.Y(n_18515)
);

XNOR2x2_ASAP7_75t_L g18516 ( 
.A(n_18314),
.B(n_8613),
.Y(n_18516)
);

INVx1_ASAP7_75t_L g18517 ( 
.A(n_18377),
.Y(n_18517)
);

NAND3xp33_ASAP7_75t_L g18518 ( 
.A(n_18277),
.B(n_5083),
.C(n_8575),
.Y(n_18518)
);

NOR4xp25_ASAP7_75t_SL g18519 ( 
.A(n_18406),
.B(n_7000),
.C(n_7004),
.D(n_8745),
.Y(n_18519)
);

INVx1_ASAP7_75t_SL g18520 ( 
.A(n_18207),
.Y(n_18520)
);

NOR3xp33_ASAP7_75t_SL g18521 ( 
.A(n_18203),
.B(n_7522),
.C(n_7491),
.Y(n_18521)
);

AOI21xp33_ASAP7_75t_L g18522 ( 
.A1(n_18274),
.A2(n_9947),
.B(n_6024),
.Y(n_18522)
);

INVx2_ASAP7_75t_L g18523 ( 
.A(n_18373),
.Y(n_18523)
);

NAND2xp33_ASAP7_75t_SL g18524 ( 
.A(n_18256),
.B(n_6706),
.Y(n_18524)
);

OAI221xp5_ASAP7_75t_L g18525 ( 
.A1(n_18388),
.A2(n_8931),
.B1(n_8922),
.B2(n_8852),
.C(n_7109),
.Y(n_18525)
);

INVx1_ASAP7_75t_L g18526 ( 
.A(n_18234),
.Y(n_18526)
);

NAND2xp5_ASAP7_75t_L g18527 ( 
.A(n_18241),
.B(n_8811),
.Y(n_18527)
);

XNOR2x2_ASAP7_75t_L g18528 ( 
.A(n_18211),
.B(n_8217),
.Y(n_18528)
);

INVx1_ASAP7_75t_SL g18529 ( 
.A(n_18358),
.Y(n_18529)
);

BUFx2_ASAP7_75t_L g18530 ( 
.A(n_18244),
.Y(n_18530)
);

HB1xp67_ASAP7_75t_L g18531 ( 
.A(n_18382),
.Y(n_18531)
);

OAI22xp5_ASAP7_75t_L g18532 ( 
.A1(n_18390),
.A2(n_7118),
.B1(n_7231),
.B2(n_7187),
.Y(n_18532)
);

XOR2xp5_ASAP7_75t_L g18533 ( 
.A(n_18299),
.B(n_6623),
.Y(n_18533)
);

OR2x2_ASAP7_75t_L g18534 ( 
.A(n_18296),
.B(n_7707),
.Y(n_18534)
);

INVxp67_ASAP7_75t_SL g18535 ( 
.A(n_18408),
.Y(n_18535)
);

INVxp67_ASAP7_75t_SL g18536 ( 
.A(n_18293),
.Y(n_18536)
);

NAND3xp33_ASAP7_75t_L g18537 ( 
.A(n_18214),
.B(n_5083),
.C(n_8575),
.Y(n_18537)
);

AOI21xp33_ASAP7_75t_SL g18538 ( 
.A1(n_18319),
.A2(n_18420),
.B(n_18302),
.Y(n_18538)
);

OAI21xp5_ASAP7_75t_L g18539 ( 
.A1(n_18375),
.A2(n_7847),
.B(n_7842),
.Y(n_18539)
);

NAND4xp25_ASAP7_75t_L g18540 ( 
.A(n_18310),
.B(n_7039),
.C(n_7007),
.D(n_7504),
.Y(n_18540)
);

NOR3xp33_ASAP7_75t_SL g18541 ( 
.A(n_18304),
.B(n_7567),
.C(n_7522),
.Y(n_18541)
);

NOR2xp33_ASAP7_75t_SL g18542 ( 
.A(n_18383),
.B(n_7039),
.Y(n_18542)
);

INVx2_ASAP7_75t_L g18543 ( 
.A(n_18342),
.Y(n_18543)
);

OAI21xp5_ASAP7_75t_L g18544 ( 
.A1(n_18300),
.A2(n_7726),
.B(n_7739),
.Y(n_18544)
);

INVx1_ASAP7_75t_SL g18545 ( 
.A(n_18303),
.Y(n_18545)
);

INVxp67_ASAP7_75t_L g18546 ( 
.A(n_18298),
.Y(n_18546)
);

INVx1_ASAP7_75t_L g18547 ( 
.A(n_18427),
.Y(n_18547)
);

INVx2_ASAP7_75t_L g18548 ( 
.A(n_18342),
.Y(n_18548)
);

NOR2xp33_ASAP7_75t_L g18549 ( 
.A(n_18270),
.B(n_6706),
.Y(n_18549)
);

AND2x2_ASAP7_75t_L g18550 ( 
.A(n_18232),
.B(n_6623),
.Y(n_18550)
);

INVx1_ASAP7_75t_L g18551 ( 
.A(n_18428),
.Y(n_18551)
);

INVx1_ASAP7_75t_SL g18552 ( 
.A(n_18278),
.Y(n_18552)
);

OR2x2_ASAP7_75t_L g18553 ( 
.A(n_18226),
.B(n_7707),
.Y(n_18553)
);

INVx1_ASAP7_75t_L g18554 ( 
.A(n_18429),
.Y(n_18554)
);

NAND2xp5_ASAP7_75t_L g18555 ( 
.A(n_18238),
.B(n_8811),
.Y(n_18555)
);

AND2x2_ASAP7_75t_L g18556 ( 
.A(n_18261),
.B(n_6623),
.Y(n_18556)
);

NOR2xp67_ASAP7_75t_L g18557 ( 
.A(n_18281),
.B(n_5465),
.Y(n_18557)
);

NAND2xp5_ASAP7_75t_L g18558 ( 
.A(n_18221),
.B(n_8811),
.Y(n_18558)
);

INVx1_ASAP7_75t_L g18559 ( 
.A(n_18436),
.Y(n_18559)
);

INVx1_ASAP7_75t_L g18560 ( 
.A(n_18440),
.Y(n_18560)
);

INVx1_ASAP7_75t_L g18561 ( 
.A(n_18283),
.Y(n_18561)
);

OAI22xp33_ASAP7_75t_SL g18562 ( 
.A1(n_18395),
.A2(n_8922),
.B1(n_8931),
.B2(n_8852),
.Y(n_18562)
);

AND2x2_ASAP7_75t_L g18563 ( 
.A(n_18262),
.B(n_6623),
.Y(n_18563)
);

HB1xp67_ASAP7_75t_L g18564 ( 
.A(n_18382),
.Y(n_18564)
);

OAI21xp5_ASAP7_75t_L g18565 ( 
.A1(n_18384),
.A2(n_7726),
.B(n_7739),
.Y(n_18565)
);

INVx1_ASAP7_75t_L g18566 ( 
.A(n_18350),
.Y(n_18566)
);

NOR4xp25_ASAP7_75t_SL g18567 ( 
.A(n_18332),
.B(n_8760),
.C(n_8783),
.D(n_8747),
.Y(n_18567)
);

AOI22xp33_ASAP7_75t_L g18568 ( 
.A1(n_18393),
.A2(n_8646),
.B1(n_8575),
.B2(n_7187),
.Y(n_18568)
);

OAI222xp33_ASAP7_75t_L g18569 ( 
.A1(n_18387),
.A2(n_18376),
.B1(n_18413),
.B2(n_18423),
.C1(n_18315),
.C2(n_18344),
.Y(n_18569)
);

CKINVDCx5p33_ASAP7_75t_R g18570 ( 
.A(n_18341),
.Y(n_18570)
);

INVx2_ASAP7_75t_L g18571 ( 
.A(n_18416),
.Y(n_18571)
);

NOR2xp33_ASAP7_75t_L g18572 ( 
.A(n_18206),
.B(n_7669),
.Y(n_18572)
);

AND2x2_ASAP7_75t_L g18573 ( 
.A(n_18258),
.B(n_6625),
.Y(n_18573)
);

NOR2xp33_ASAP7_75t_R g18574 ( 
.A(n_18327),
.B(n_5834),
.Y(n_18574)
);

NOR2x1_ASAP7_75t_L g18575 ( 
.A(n_18397),
.B(n_8206),
.Y(n_18575)
);

AND2x4_ASAP7_75t_L g18576 ( 
.A(n_18339),
.B(n_7039),
.Y(n_18576)
);

INVxp33_ASAP7_75t_L g18577 ( 
.A(n_18417),
.Y(n_18577)
);

OAI22xp5_ASAP7_75t_L g18578 ( 
.A1(n_18343),
.A2(n_7118),
.B1(n_7231),
.B2(n_7187),
.Y(n_18578)
);

INVxp67_ASAP7_75t_SL g18579 ( 
.A(n_18345),
.Y(n_18579)
);

INVx2_ASAP7_75t_L g18580 ( 
.A(n_18289),
.Y(n_18580)
);

NOR2xp33_ASAP7_75t_L g18581 ( 
.A(n_18249),
.B(n_7669),
.Y(n_18581)
);

INVx1_ASAP7_75t_L g18582 ( 
.A(n_18272),
.Y(n_18582)
);

INVx1_ASAP7_75t_L g18583 ( 
.A(n_18257),
.Y(n_18583)
);

OAI21xp5_ASAP7_75t_L g18584 ( 
.A1(n_18259),
.A2(n_7726),
.B(n_7739),
.Y(n_18584)
);

INVx1_ASAP7_75t_L g18585 ( 
.A(n_18363),
.Y(n_18585)
);

NOR3xp33_ASAP7_75t_L g18586 ( 
.A(n_18369),
.B(n_5400),
.C(n_5363),
.Y(n_18586)
);

NAND2xp5_ASAP7_75t_L g18587 ( 
.A(n_18330),
.B(n_8824),
.Y(n_18587)
);

NAND2xp5_ASAP7_75t_L g18588 ( 
.A(n_18320),
.B(n_18248),
.Y(n_18588)
);

INVx2_ASAP7_75t_L g18589 ( 
.A(n_18365),
.Y(n_18589)
);

AOI22xp5_ASAP7_75t_L g18590 ( 
.A1(n_18374),
.A2(n_7231),
.B1(n_7258),
.B2(n_7118),
.Y(n_18590)
);

INVx1_ASAP7_75t_L g18591 ( 
.A(n_18280),
.Y(n_18591)
);

NOR2xp33_ASAP7_75t_L g18592 ( 
.A(n_18398),
.B(n_18333),
.Y(n_18592)
);

INVx6_ASAP7_75t_L g18593 ( 
.A(n_18317),
.Y(n_18593)
);

HB1xp67_ASAP7_75t_L g18594 ( 
.A(n_18318),
.Y(n_18594)
);

INVx1_ASAP7_75t_L g18595 ( 
.A(n_18325),
.Y(n_18595)
);

NAND2xp5_ASAP7_75t_L g18596 ( 
.A(n_18336),
.B(n_8824),
.Y(n_18596)
);

NAND2xp5_ASAP7_75t_L g18597 ( 
.A(n_18337),
.B(n_8824),
.Y(n_18597)
);

AND2x2_ASAP7_75t_L g18598 ( 
.A(n_18223),
.B(n_6625),
.Y(n_18598)
);

XOR2x2_ASAP7_75t_L g18599 ( 
.A(n_18294),
.B(n_5871),
.Y(n_18599)
);

NAND2xp5_ASAP7_75t_L g18600 ( 
.A(n_18329),
.B(n_8858),
.Y(n_18600)
);

AND2x2_ASAP7_75t_L g18601 ( 
.A(n_18230),
.B(n_6625),
.Y(n_18601)
);

NAND2xp5_ASAP7_75t_L g18602 ( 
.A(n_18366),
.B(n_8858),
.Y(n_18602)
);

INVx1_ASAP7_75t_SL g18603 ( 
.A(n_18367),
.Y(n_18603)
);

AND2x2_ASAP7_75t_L g18604 ( 
.A(n_18217),
.B(n_18225),
.Y(n_18604)
);

INVx1_ASAP7_75t_L g18605 ( 
.A(n_18338),
.Y(n_18605)
);

INVxp67_ASAP7_75t_L g18606 ( 
.A(n_18364),
.Y(n_18606)
);

AND2x2_ASAP7_75t_L g18607 ( 
.A(n_18361),
.B(n_6625),
.Y(n_18607)
);

INVx1_ASAP7_75t_L g18608 ( 
.A(n_18331),
.Y(n_18608)
);

OAI21xp5_ASAP7_75t_SL g18609 ( 
.A1(n_18237),
.A2(n_18236),
.B(n_18356),
.Y(n_18609)
);

NOR2xp33_ASAP7_75t_L g18610 ( 
.A(n_18243),
.B(n_7669),
.Y(n_18610)
);

AND2x2_ASAP7_75t_L g18611 ( 
.A(n_18371),
.B(n_6625),
.Y(n_18611)
);

INVx3_ASAP7_75t_L g18612 ( 
.A(n_18265),
.Y(n_18612)
);

OAI22xp5_ASAP7_75t_L g18613 ( 
.A1(n_18351),
.A2(n_7258),
.B1(n_7260),
.B2(n_7231),
.Y(n_18613)
);

INVx1_ASAP7_75t_L g18614 ( 
.A(n_18354),
.Y(n_18614)
);

OR2x2_ASAP7_75t_L g18615 ( 
.A(n_18349),
.B(n_7707),
.Y(n_18615)
);

AND2x2_ASAP7_75t_L g18616 ( 
.A(n_18346),
.B(n_6625),
.Y(n_18616)
);

NAND2xp5_ASAP7_75t_L g18617 ( 
.A(n_18355),
.B(n_18402),
.Y(n_18617)
);

INVxp67_ASAP7_75t_L g18618 ( 
.A(n_18323),
.Y(n_18618)
);

AND2x2_ASAP7_75t_L g18619 ( 
.A(n_18360),
.B(n_18348),
.Y(n_18619)
);

NAND2xp5_ASAP7_75t_L g18620 ( 
.A(n_18291),
.B(n_8858),
.Y(n_18620)
);

NAND2xp5_ASAP7_75t_L g18621 ( 
.A(n_18295),
.B(n_8861),
.Y(n_18621)
);

NAND2xp5_ASAP7_75t_L g18622 ( 
.A(n_18273),
.B(n_8861),
.Y(n_18622)
);

INVx1_ASAP7_75t_L g18623 ( 
.A(n_18316),
.Y(n_18623)
);

OAI32xp33_ASAP7_75t_L g18624 ( 
.A1(n_18334),
.A2(n_8882),
.A3(n_8889),
.B1(n_8881),
.B2(n_8861),
.Y(n_18624)
);

INVx1_ASAP7_75t_L g18625 ( 
.A(n_18352),
.Y(n_18625)
);

XNOR2xp5_ASAP7_75t_L g18626 ( 
.A(n_18430),
.B(n_8922),
.Y(n_18626)
);

AND2x2_ASAP7_75t_L g18627 ( 
.A(n_18370),
.B(n_6646),
.Y(n_18627)
);

O2A1O1Ixp5_ASAP7_75t_L g18628 ( 
.A1(n_18418),
.A2(n_8882),
.B(n_8889),
.C(n_8881),
.Y(n_18628)
);

CKINVDCx14_ASAP7_75t_R g18629 ( 
.A(n_18308),
.Y(n_18629)
);

INVx3_ASAP7_75t_L g18630 ( 
.A(n_18276),
.Y(n_18630)
);

INVx1_ASAP7_75t_L g18631 ( 
.A(n_18372),
.Y(n_18631)
);

INVx1_ASAP7_75t_L g18632 ( 
.A(n_18362),
.Y(n_18632)
);

AOI22xp5_ASAP7_75t_L g18633 ( 
.A1(n_18425),
.A2(n_7260),
.B1(n_7295),
.B2(n_7258),
.Y(n_18633)
);

AND2x2_ASAP7_75t_L g18634 ( 
.A(n_18301),
.B(n_6646),
.Y(n_18634)
);

AND2x2_ASAP7_75t_L g18635 ( 
.A(n_18267),
.B(n_6646),
.Y(n_18635)
);

NAND2xp5_ASAP7_75t_L g18636 ( 
.A(n_18335),
.B(n_18307),
.Y(n_18636)
);

AND2x4_ASAP7_75t_L g18637 ( 
.A(n_18353),
.B(n_7039),
.Y(n_18637)
);

OR2x2_ASAP7_75t_L g18638 ( 
.A(n_18380),
.B(n_7707),
.Y(n_18638)
);

AND2x2_ASAP7_75t_L g18639 ( 
.A(n_18405),
.B(n_6646),
.Y(n_18639)
);

OR2x2_ASAP7_75t_L g18640 ( 
.A(n_18404),
.B(n_7707),
.Y(n_18640)
);

INVxp67_ASAP7_75t_L g18641 ( 
.A(n_18403),
.Y(n_18641)
);

NAND2xp5_ASAP7_75t_L g18642 ( 
.A(n_18326),
.B(n_8881),
.Y(n_18642)
);

AND2x4_ASAP7_75t_SL g18643 ( 
.A(n_18322),
.B(n_7272),
.Y(n_18643)
);

AOI221xp5_ASAP7_75t_L g18644 ( 
.A1(n_18422),
.A2(n_7258),
.B1(n_7326),
.B2(n_7295),
.C(n_7260),
.Y(n_18644)
);

NOR2xp33_ASAP7_75t_L g18645 ( 
.A(n_18409),
.B(n_7669),
.Y(n_18645)
);

NAND2xp5_ASAP7_75t_L g18646 ( 
.A(n_18328),
.B(n_8882),
.Y(n_18646)
);

INVx1_ASAP7_75t_L g18647 ( 
.A(n_18313),
.Y(n_18647)
);

AOI22xp5_ASAP7_75t_L g18648 ( 
.A1(n_18263),
.A2(n_7295),
.B1(n_7326),
.B2(n_7260),
.Y(n_18648)
);

NOR2x1_ASAP7_75t_L g18649 ( 
.A(n_18392),
.B(n_8206),
.Y(n_18649)
);

AOI22xp5_ASAP7_75t_L g18650 ( 
.A1(n_18542),
.A2(n_18242),
.B1(n_18401),
.B2(n_18396),
.Y(n_18650)
);

OA22x2_ASAP7_75t_L g18651 ( 
.A1(n_18472),
.A2(n_18389),
.B1(n_18391),
.B2(n_18407),
.Y(n_18651)
);

NOR3xp33_ASAP7_75t_SL g18652 ( 
.A(n_18569),
.B(n_18368),
.C(n_18340),
.Y(n_18652)
);

INVx2_ASAP7_75t_L g18653 ( 
.A(n_18528),
.Y(n_18653)
);

AOI22xp5_ASAP7_75t_L g18654 ( 
.A1(n_18467),
.A2(n_18385),
.B1(n_18399),
.B2(n_18386),
.Y(n_18654)
);

NAND2xp5_ASAP7_75t_L g18655 ( 
.A(n_18445),
.B(n_18347),
.Y(n_18655)
);

OA22x2_ASAP7_75t_L g18656 ( 
.A1(n_18504),
.A2(n_18419),
.B1(n_18357),
.B2(n_18385),
.Y(n_18656)
);

NAND2xp5_ASAP7_75t_L g18657 ( 
.A(n_18470),
.B(n_18379),
.Y(n_18657)
);

OA22x2_ASAP7_75t_L g18658 ( 
.A1(n_18451),
.A2(n_18305),
.B1(n_18394),
.B2(n_18411),
.Y(n_18658)
);

AOI21xp5_ASAP7_75t_L g18659 ( 
.A1(n_18579),
.A2(n_18421),
.B(n_8931),
.Y(n_18659)
);

AOI22xp5_ASAP7_75t_SL g18660 ( 
.A1(n_18536),
.A2(n_8320),
.B1(n_8188),
.B2(n_8646),
.Y(n_18660)
);

AOI21xp5_ASAP7_75t_L g18661 ( 
.A1(n_18535),
.A2(n_8931),
.B(n_8922),
.Y(n_18661)
);

NOR3x1_ASAP7_75t_L g18662 ( 
.A(n_18494),
.B(n_8515),
.C(n_8502),
.Y(n_18662)
);

INVx1_ASAP7_75t_L g18663 ( 
.A(n_18533),
.Y(n_18663)
);

AO22x2_ASAP7_75t_L g18664 ( 
.A1(n_18452),
.A2(n_18459),
.B1(n_18458),
.B2(n_18449),
.Y(n_18664)
);

INVx1_ASAP7_75t_L g18665 ( 
.A(n_18456),
.Y(n_18665)
);

AO22x2_ASAP7_75t_L g18666 ( 
.A1(n_18501),
.A2(n_18492),
.B1(n_18468),
.B2(n_18476),
.Y(n_18666)
);

AOI22xp5_ASAP7_75t_L g18667 ( 
.A1(n_18508),
.A2(n_7326),
.B1(n_7330),
.B2(n_7295),
.Y(n_18667)
);

INVx1_ASAP7_75t_L g18668 ( 
.A(n_18462),
.Y(n_18668)
);

OA22x2_ASAP7_75t_L g18669 ( 
.A1(n_18545),
.A2(n_7330),
.B1(n_7338),
.B2(n_7326),
.Y(n_18669)
);

INVx2_ASAP7_75t_SL g18670 ( 
.A(n_18441),
.Y(n_18670)
);

AND2x2_ASAP7_75t_L g18671 ( 
.A(n_18483),
.B(n_6646),
.Y(n_18671)
);

NOR3x1_ASAP7_75t_L g18672 ( 
.A(n_18506),
.B(n_8523),
.C(n_8515),
.Y(n_18672)
);

NAND2x1p5_ASAP7_75t_L g18673 ( 
.A(n_18529),
.B(n_5180),
.Y(n_18673)
);

AOI21xp5_ASAP7_75t_L g18674 ( 
.A1(n_18588),
.A2(n_8931),
.B(n_8922),
.Y(n_18674)
);

OAI21xp33_ASAP7_75t_SL g18675 ( 
.A1(n_18568),
.A2(n_8523),
.B(n_8515),
.Y(n_18675)
);

AOI21xp5_ASAP7_75t_L g18676 ( 
.A1(n_18577),
.A2(n_9947),
.B(n_7059),
.Y(n_18676)
);

NOR2x1_ASAP7_75t_L g18677 ( 
.A(n_18454),
.B(n_5363),
.Y(n_18677)
);

INVx1_ASAP7_75t_SL g18678 ( 
.A(n_18477),
.Y(n_18678)
);

AOI211x1_ASAP7_75t_L g18679 ( 
.A1(n_18565),
.A2(n_8783),
.B(n_8789),
.C(n_8760),
.Y(n_18679)
);

AOI21xp5_ASAP7_75t_SL g18680 ( 
.A1(n_18471),
.A2(n_5960),
.B(n_5891),
.Y(n_18680)
);

NOR2x1_ASAP7_75t_L g18681 ( 
.A(n_18530),
.B(n_5400),
.Y(n_18681)
);

NOR2x1_ASAP7_75t_L g18682 ( 
.A(n_18513),
.B(n_5400),
.Y(n_18682)
);

AND2x2_ASAP7_75t_L g18683 ( 
.A(n_18481),
.B(n_6646),
.Y(n_18683)
);

OAI21xp33_ASAP7_75t_SL g18684 ( 
.A1(n_18649),
.A2(n_8523),
.B(n_8233),
.Y(n_18684)
);

NAND2xp5_ASAP7_75t_L g18685 ( 
.A(n_18576),
.B(n_8889),
.Y(n_18685)
);

INVx2_ASAP7_75t_L g18686 ( 
.A(n_18485),
.Y(n_18686)
);

AOI22xp5_ASAP7_75t_L g18687 ( 
.A1(n_18491),
.A2(n_18512),
.B1(n_18520),
.B2(n_18480),
.Y(n_18687)
);

NOR3x1_ASAP7_75t_L g18688 ( 
.A(n_18609),
.B(n_18489),
.C(n_18517),
.Y(n_18688)
);

AOI22xp5_ASAP7_75t_L g18689 ( 
.A1(n_18511),
.A2(n_7338),
.B1(n_7403),
.B2(n_7330),
.Y(n_18689)
);

INVx1_ASAP7_75t_L g18690 ( 
.A(n_18531),
.Y(n_18690)
);

AO22x2_ASAP7_75t_L g18691 ( 
.A1(n_18461),
.A2(n_8910),
.B1(n_8914),
.B2(n_8905),
.Y(n_18691)
);

AOI21xp5_ASAP7_75t_L g18692 ( 
.A1(n_18617),
.A2(n_9947),
.B(n_7059),
.Y(n_18692)
);

OA22x2_ASAP7_75t_L g18693 ( 
.A1(n_18590),
.A2(n_7338),
.B1(n_7403),
.B2(n_7330),
.Y(n_18693)
);

NAND3xp33_ASAP7_75t_L g18694 ( 
.A(n_18538),
.B(n_5083),
.C(n_5180),
.Y(n_18694)
);

NAND4xp75_ASAP7_75t_L g18695 ( 
.A(n_18561),
.B(n_8320),
.C(n_8646),
.D(n_8188),
.Y(n_18695)
);

AOI22xp5_ASAP7_75t_L g18696 ( 
.A1(n_18549),
.A2(n_7403),
.B1(n_7414),
.B2(n_7338),
.Y(n_18696)
);

OAI211xp5_ASAP7_75t_SL g18697 ( 
.A1(n_18546),
.A2(n_5490),
.B(n_4598),
.C(n_4618),
.Y(n_18697)
);

NAND2xp5_ASAP7_75t_L g18698 ( 
.A(n_18576),
.B(n_8905),
.Y(n_18698)
);

NAND2xp5_ASAP7_75t_L g18699 ( 
.A(n_18523),
.B(n_8905),
.Y(n_18699)
);

INVx2_ASAP7_75t_L g18700 ( 
.A(n_18499),
.Y(n_18700)
);

CKINVDCx5p33_ASAP7_75t_R g18701 ( 
.A(n_18570),
.Y(n_18701)
);

AOI22xp5_ASAP7_75t_L g18702 ( 
.A1(n_18450),
.A2(n_7414),
.B1(n_7423),
.B2(n_7403),
.Y(n_18702)
);

NAND2xp5_ASAP7_75t_L g18703 ( 
.A(n_18571),
.B(n_8910),
.Y(n_18703)
);

NOR2xp67_ASAP7_75t_L g18704 ( 
.A(n_18612),
.B(n_5490),
.Y(n_18704)
);

AOI211x1_ASAP7_75t_SL g18705 ( 
.A1(n_18532),
.A2(n_8914),
.B(n_8920),
.C(n_8910),
.Y(n_18705)
);

INVx1_ASAP7_75t_L g18706 ( 
.A(n_18564),
.Y(n_18706)
);

INVx1_ASAP7_75t_L g18707 ( 
.A(n_18464),
.Y(n_18707)
);

NAND2xp5_ASAP7_75t_L g18708 ( 
.A(n_18585),
.B(n_8914),
.Y(n_18708)
);

AOI211x1_ASAP7_75t_L g18709 ( 
.A1(n_18525),
.A2(n_8804),
.B(n_8808),
.C(n_8789),
.Y(n_18709)
);

NOR2xp33_ASAP7_75t_L g18710 ( 
.A(n_18475),
.B(n_7039),
.Y(n_18710)
);

OAI21xp33_ASAP7_75t_L g18711 ( 
.A1(n_18572),
.A2(n_7423),
.B(n_7414),
.Y(n_18711)
);

OAI21xp5_ASAP7_75t_L g18712 ( 
.A1(n_18495),
.A2(n_7743),
.B(n_7878),
.Y(n_18712)
);

OAI211xp5_ASAP7_75t_L g18713 ( 
.A1(n_18629),
.A2(n_7207),
.B(n_7239),
.C(n_7230),
.Y(n_18713)
);

INVx1_ASAP7_75t_L g18714 ( 
.A(n_18619),
.Y(n_18714)
);

AOI21xp5_ASAP7_75t_L g18715 ( 
.A1(n_18524),
.A2(n_7059),
.B(n_7040),
.Y(n_18715)
);

AND4x1_ASAP7_75t_L g18716 ( 
.A(n_18592),
.B(n_7567),
.C(n_7568),
.D(n_7040),
.Y(n_18716)
);

NAND2xp5_ASAP7_75t_L g18717 ( 
.A(n_18630),
.B(n_8920),
.Y(n_18717)
);

NAND4xp25_ASAP7_75t_L g18718 ( 
.A(n_18566),
.B(n_4967),
.C(n_5045),
.D(n_4933),
.Y(n_18718)
);

INVx2_ASAP7_75t_L g18719 ( 
.A(n_18637),
.Y(n_18719)
);

INVx2_ASAP7_75t_L g18720 ( 
.A(n_18637),
.Y(n_18720)
);

OAI21xp5_ASAP7_75t_SL g18721 ( 
.A1(n_18603),
.A2(n_5470),
.B(n_7523),
.Y(n_18721)
);

NAND2xp5_ASAP7_75t_SL g18722 ( 
.A(n_18500),
.B(n_6670),
.Y(n_18722)
);

NOR2xp33_ASAP7_75t_L g18723 ( 
.A(n_18479),
.B(n_7039),
.Y(n_18723)
);

NAND2xp5_ASAP7_75t_L g18724 ( 
.A(n_18552),
.B(n_8920),
.Y(n_18724)
);

NAND4xp25_ASAP7_75t_SL g18725 ( 
.A(n_18448),
.B(n_7434),
.C(n_7524),
.D(n_7451),
.Y(n_18725)
);

OAI22xp5_ASAP7_75t_L g18726 ( 
.A1(n_18443),
.A2(n_7423),
.B1(n_7428),
.B2(n_7414),
.Y(n_18726)
);

NOR3x1_ASAP7_75t_L g18727 ( 
.A(n_18595),
.B(n_7916),
.C(n_8217),
.Y(n_18727)
);

AOI22xp5_ASAP7_75t_L g18728 ( 
.A1(n_18645),
.A2(n_7428),
.B1(n_7442),
.B2(n_7423),
.Y(n_18728)
);

NOR2xp67_ASAP7_75t_SL g18729 ( 
.A(n_18614),
.B(n_5453),
.Y(n_18729)
);

OAI21xp5_ASAP7_75t_L g18730 ( 
.A1(n_18606),
.A2(n_7743),
.B(n_7878),
.Y(n_18730)
);

AOI211xp5_ASAP7_75t_L g18731 ( 
.A1(n_18641),
.A2(n_8204),
.B(n_8207),
.C(n_7916),
.Y(n_18731)
);

AOI22xp5_ASAP7_75t_L g18732 ( 
.A1(n_18581),
.A2(n_7442),
.B1(n_7466),
.B2(n_7428),
.Y(n_18732)
);

INVx1_ASAP7_75t_L g18733 ( 
.A(n_18557),
.Y(n_18733)
);

NAND4xp25_ASAP7_75t_L g18734 ( 
.A(n_18498),
.B(n_4967),
.C(n_5045),
.D(n_4933),
.Y(n_18734)
);

AOI21xp5_ASAP7_75t_L g18735 ( 
.A1(n_18636),
.A2(n_7040),
.B(n_7567),
.Y(n_18735)
);

O2A1O1Ixp33_ASAP7_75t_L g18736 ( 
.A1(n_18497),
.A2(n_4601),
.B(n_4618),
.C(n_4598),
.Y(n_18736)
);

NAND4xp75_ASAP7_75t_L g18737 ( 
.A(n_18605),
.B(n_8320),
.C(n_8188),
.D(n_4953),
.Y(n_18737)
);

INVx1_ASAP7_75t_L g18738 ( 
.A(n_18496),
.Y(n_18738)
);

OAI211xp5_ASAP7_75t_L g18739 ( 
.A1(n_18589),
.A2(n_7230),
.B(n_7285),
.C(n_7239),
.Y(n_18739)
);

AOI211xp5_ASAP7_75t_L g18740 ( 
.A1(n_18608),
.A2(n_8204),
.B(n_8207),
.C(n_7916),
.Y(n_18740)
);

O2A1O1Ixp33_ASAP7_75t_SL g18741 ( 
.A1(n_18543),
.A2(n_7442),
.B(n_7466),
.C(n_7428),
.Y(n_18741)
);

NAND2xp5_ASAP7_75t_L g18742 ( 
.A(n_18493),
.B(n_8924),
.Y(n_18742)
);

NOR2xp33_ASAP7_75t_L g18743 ( 
.A(n_18484),
.B(n_18486),
.Y(n_18743)
);

INVx1_ASAP7_75t_L g18744 ( 
.A(n_18604),
.Y(n_18744)
);

OR2x2_ASAP7_75t_L g18745 ( 
.A(n_18460),
.B(n_7707),
.Y(n_18745)
);

INVx1_ASAP7_75t_L g18746 ( 
.A(n_18473),
.Y(n_18746)
);

XNOR2x1_ASAP7_75t_SL g18747 ( 
.A(n_18505),
.B(n_4946),
.Y(n_18747)
);

AOI22xp33_ASAP7_75t_L g18748 ( 
.A1(n_18442),
.A2(n_7466),
.B1(n_7528),
.B2(n_7442),
.Y(n_18748)
);

AOI21xp5_ASAP7_75t_L g18749 ( 
.A1(n_18618),
.A2(n_7568),
.B(n_7354),
.Y(n_18749)
);

NOR3xp33_ASAP7_75t_L g18750 ( 
.A(n_18631),
.B(n_5400),
.C(n_4967),
.Y(n_18750)
);

NOR2x1_ASAP7_75t_L g18751 ( 
.A(n_18548),
.B(n_5400),
.Y(n_18751)
);

AOI21xp5_ASAP7_75t_L g18752 ( 
.A1(n_18580),
.A2(n_7568),
.B(n_7354),
.Y(n_18752)
);

NAND2xp5_ASAP7_75t_L g18753 ( 
.A(n_18526),
.B(n_8924),
.Y(n_18753)
);

AND2x2_ASAP7_75t_L g18754 ( 
.A(n_18521),
.B(n_18550),
.Y(n_18754)
);

NOR3xp33_ASAP7_75t_L g18755 ( 
.A(n_18625),
.B(n_5400),
.C(n_4967),
.Y(n_18755)
);

AOI31xp33_ASAP7_75t_L g18756 ( 
.A1(n_18594),
.A2(n_4953),
.A3(n_4957),
.B(n_4946),
.Y(n_18756)
);

INVx1_ASAP7_75t_L g18757 ( 
.A(n_18593),
.Y(n_18757)
);

NOR2x1_ASAP7_75t_L g18758 ( 
.A(n_18547),
.B(n_8206),
.Y(n_18758)
);

XNOR2x1_ASAP7_75t_SL g18759 ( 
.A(n_18623),
.B(n_4946),
.Y(n_18759)
);

AOI22xp5_ASAP7_75t_L g18760 ( 
.A1(n_18610),
.A2(n_7528),
.B1(n_7581),
.B2(n_7466),
.Y(n_18760)
);

NOR2xp33_ASAP7_75t_L g18761 ( 
.A(n_18593),
.B(n_18632),
.Y(n_18761)
);

NAND4xp25_ASAP7_75t_L g18762 ( 
.A(n_18490),
.B(n_5045),
.C(n_5078),
.D(n_4933),
.Y(n_18762)
);

INVx1_ASAP7_75t_L g18763 ( 
.A(n_18507),
.Y(n_18763)
);

AOI211x1_ASAP7_75t_L g18764 ( 
.A1(n_18469),
.A2(n_8808),
.B(n_8819),
.C(n_8804),
.Y(n_18764)
);

NOR3xp33_ASAP7_75t_SL g18765 ( 
.A(n_18551),
.B(n_7344),
.C(n_7421),
.Y(n_18765)
);

INVx2_ASAP7_75t_L g18766 ( 
.A(n_18446),
.Y(n_18766)
);

NOR2x1_ASAP7_75t_L g18767 ( 
.A(n_18554),
.B(n_8258),
.Y(n_18767)
);

NAND2xp5_ASAP7_75t_SL g18768 ( 
.A(n_18503),
.B(n_6670),
.Y(n_18768)
);

OA22x2_ASAP7_75t_L g18769 ( 
.A1(n_18643),
.A2(n_7581),
.B1(n_7587),
.B2(n_7528),
.Y(n_18769)
);

INVx2_ASAP7_75t_SL g18770 ( 
.A(n_18574),
.Y(n_18770)
);

NOR2x1_ASAP7_75t_L g18771 ( 
.A(n_18559),
.B(n_8258),
.Y(n_18771)
);

NAND4xp25_ASAP7_75t_L g18772 ( 
.A(n_18596),
.B(n_5045),
.C(n_5078),
.D(n_4933),
.Y(n_18772)
);

INVx1_ASAP7_75t_L g18773 ( 
.A(n_18560),
.Y(n_18773)
);

NAND2xp5_ASAP7_75t_L g18774 ( 
.A(n_18582),
.B(n_18583),
.Y(n_18774)
);

INVx2_ASAP7_75t_L g18775 ( 
.A(n_18447),
.Y(n_18775)
);

INVxp33_ASAP7_75t_SL g18776 ( 
.A(n_18647),
.Y(n_18776)
);

INVx1_ASAP7_75t_L g18777 ( 
.A(n_18591),
.Y(n_18777)
);

HB1xp67_ASAP7_75t_SL g18778 ( 
.A(n_18534),
.Y(n_18778)
);

NOR3xp33_ASAP7_75t_L g18779 ( 
.A(n_18602),
.B(n_5078),
.C(n_5045),
.Y(n_18779)
);

NAND2xp5_ASAP7_75t_L g18780 ( 
.A(n_18556),
.B(n_8924),
.Y(n_18780)
);

OAI22xp5_ASAP7_75t_L g18781 ( 
.A1(n_18537),
.A2(n_7581),
.B1(n_7587),
.B2(n_7528),
.Y(n_18781)
);

NOR3x1_ASAP7_75t_L g18782 ( 
.A(n_18597),
.B(n_8233),
.C(n_8217),
.Y(n_18782)
);

AND2x2_ASAP7_75t_L g18783 ( 
.A(n_18563),
.B(n_6853),
.Y(n_18783)
);

NAND2xp5_ASAP7_75t_L g18784 ( 
.A(n_18607),
.B(n_8930),
.Y(n_18784)
);

NAND2xp5_ASAP7_75t_SL g18785 ( 
.A(n_18613),
.B(n_6670),
.Y(n_18785)
);

NOR3xp33_ASAP7_75t_L g18786 ( 
.A(n_18600),
.B(n_5078),
.C(n_5045),
.Y(n_18786)
);

AOI221xp5_ASAP7_75t_L g18787 ( 
.A1(n_18510),
.A2(n_8956),
.B1(n_8967),
.B2(n_8946),
.C(n_8930),
.Y(n_18787)
);

NOR3xp33_ASAP7_75t_L g18788 ( 
.A(n_18465),
.B(n_5125),
.C(n_5078),
.Y(n_18788)
);

NOR3xp33_ASAP7_75t_L g18789 ( 
.A(n_18466),
.B(n_5125),
.C(n_5078),
.Y(n_18789)
);

NOR2x1_ASAP7_75t_L g18790 ( 
.A(n_18488),
.B(n_18640),
.Y(n_18790)
);

OAI211xp5_ASAP7_75t_SL g18791 ( 
.A1(n_18558),
.A2(n_4598),
.B(n_4618),
.C(n_4601),
.Y(n_18791)
);

XNOR2x1_ASAP7_75t_L g18792 ( 
.A(n_18599),
.B(n_7931),
.Y(n_18792)
);

INVx1_ASAP7_75t_L g18793 ( 
.A(n_18622),
.Y(n_18793)
);

NOR2xp33_ASAP7_75t_L g18794 ( 
.A(n_18626),
.B(n_7272),
.Y(n_18794)
);

AOI21xp5_ASAP7_75t_L g18795 ( 
.A1(n_18628),
.A2(n_5470),
.B(n_7581),
.Y(n_18795)
);

AOI22xp5_ASAP7_75t_L g18796 ( 
.A1(n_18482),
.A2(n_7591),
.B1(n_7654),
.B2(n_7587),
.Y(n_18796)
);

NAND2xp5_ASAP7_75t_L g18797 ( 
.A(n_18541),
.B(n_8930),
.Y(n_18797)
);

NOR2xp33_ASAP7_75t_L g18798 ( 
.A(n_18509),
.B(n_7272),
.Y(n_18798)
);

OAI21xp5_ASAP7_75t_SL g18799 ( 
.A1(n_18463),
.A2(n_5470),
.B(n_7523),
.Y(n_18799)
);

AOI22xp5_ASAP7_75t_L g18800 ( 
.A1(n_18586),
.A2(n_7591),
.B1(n_7654),
.B2(n_7587),
.Y(n_18800)
);

NOR2xp33_ASAP7_75t_L g18801 ( 
.A(n_18502),
.B(n_7272),
.Y(n_18801)
);

AOI22xp5_ASAP7_75t_L g18802 ( 
.A1(n_18639),
.A2(n_7654),
.B1(n_7671),
.B2(n_7591),
.Y(n_18802)
);

NAND2xp5_ASAP7_75t_L g18803 ( 
.A(n_18487),
.B(n_8946),
.Y(n_18803)
);

AOI21xp5_ASAP7_75t_L g18804 ( 
.A1(n_18527),
.A2(n_7654),
.B(n_7591),
.Y(n_18804)
);

NAND2xp5_ASAP7_75t_L g18805 ( 
.A(n_18515),
.B(n_8946),
.Y(n_18805)
);

INVx2_ASAP7_75t_SL g18806 ( 
.A(n_18455),
.Y(n_18806)
);

AND2x2_ASAP7_75t_L g18807 ( 
.A(n_18573),
.B(n_6853),
.Y(n_18807)
);

NAND4xp75_ASAP7_75t_L g18808 ( 
.A(n_18575),
.B(n_8320),
.C(n_8188),
.D(n_5011),
.Y(n_18808)
);

INVx2_ASAP7_75t_L g18809 ( 
.A(n_18615),
.Y(n_18809)
);

NOR2x1_ASAP7_75t_L g18810 ( 
.A(n_18638),
.B(n_8258),
.Y(n_18810)
);

NAND2x1_ASAP7_75t_SL g18811 ( 
.A(n_18598),
.B(n_8956),
.Y(n_18811)
);

OAI22xp5_ASAP7_75t_R g18812 ( 
.A1(n_18519),
.A2(n_7075),
.B1(n_8821),
.B2(n_8819),
.Y(n_18812)
);

AOI21xp5_ASAP7_75t_SL g18813 ( 
.A1(n_18587),
.A2(n_5960),
.B(n_5891),
.Y(n_18813)
);

AOI211x1_ASAP7_75t_L g18814 ( 
.A1(n_18555),
.A2(n_8828),
.B(n_8831),
.C(n_8821),
.Y(n_18814)
);

AND4x1_ASAP7_75t_L g18815 ( 
.A(n_18478),
.B(n_7421),
.C(n_7441),
.D(n_7422),
.Y(n_18815)
);

AOI211x1_ASAP7_75t_L g18816 ( 
.A1(n_18522),
.A2(n_18578),
.B(n_18621),
.C(n_18620),
.Y(n_18816)
);

INVx1_ASAP7_75t_L g18817 ( 
.A(n_18642),
.Y(n_18817)
);

AOI211xp5_ASAP7_75t_L g18818 ( 
.A1(n_18562),
.A2(n_8207),
.B(n_7878),
.C(n_7894),
.Y(n_18818)
);

HB1xp67_ASAP7_75t_L g18819 ( 
.A(n_18516),
.Y(n_18819)
);

OA22x2_ASAP7_75t_L g18820 ( 
.A1(n_18648),
.A2(n_7671),
.B1(n_8967),
.B2(n_8956),
.Y(n_18820)
);

INVx1_ASAP7_75t_L g18821 ( 
.A(n_18646),
.Y(n_18821)
);

INVx1_ASAP7_75t_L g18822 ( 
.A(n_18601),
.Y(n_18822)
);

NOR3xp33_ASAP7_75t_SL g18823 ( 
.A(n_18540),
.B(n_7441),
.C(n_7422),
.Y(n_18823)
);

AOI22xp5_ASAP7_75t_SL g18824 ( 
.A1(n_18611),
.A2(n_18627),
.B1(n_18616),
.B2(n_18634),
.Y(n_18824)
);

AOI22xp5_ASAP7_75t_SL g18825 ( 
.A1(n_18474),
.A2(n_8320),
.B1(n_8188),
.B2(n_5180),
.Y(n_18825)
);

OAI21xp5_ASAP7_75t_L g18826 ( 
.A1(n_18518),
.A2(n_7743),
.B(n_7885),
.Y(n_18826)
);

INVx2_ASAP7_75t_L g18827 ( 
.A(n_18553),
.Y(n_18827)
);

AOI211x1_ASAP7_75t_L g18828 ( 
.A1(n_18624),
.A2(n_8831),
.B(n_8848),
.C(n_8828),
.Y(n_18828)
);

NOR2x1_ASAP7_75t_L g18829 ( 
.A(n_18635),
.B(n_8258),
.Y(n_18829)
);

INVx1_ASAP7_75t_L g18830 ( 
.A(n_18453),
.Y(n_18830)
);

HB1xp67_ASAP7_75t_L g18831 ( 
.A(n_18759),
.Y(n_18831)
);

XNOR2x2_ASAP7_75t_L g18832 ( 
.A(n_18666),
.B(n_18444),
.Y(n_18832)
);

O2A1O1Ixp33_ASAP7_75t_L g18833 ( 
.A1(n_18819),
.A2(n_18714),
.B(n_18690),
.C(n_18706),
.Y(n_18833)
);

OAI22xp5_ASAP7_75t_L g18834 ( 
.A1(n_18687),
.A2(n_18457),
.B1(n_18567),
.B2(n_18633),
.Y(n_18834)
);

OAI21xp5_ASAP7_75t_L g18835 ( 
.A1(n_18659),
.A2(n_18761),
.B(n_18757),
.Y(n_18835)
);

XNOR2x1_ASAP7_75t_L g18836 ( 
.A(n_18666),
.B(n_18539),
.Y(n_18836)
);

INVx2_ASAP7_75t_SL g18837 ( 
.A(n_18664),
.Y(n_18837)
);

NAND2xp5_ASAP7_75t_L g18838 ( 
.A(n_18683),
.B(n_18664),
.Y(n_18838)
);

AOI22xp5_ASAP7_75t_L g18839 ( 
.A1(n_18744),
.A2(n_18644),
.B1(n_18544),
.B2(n_18584),
.Y(n_18839)
);

AOI21xp33_ASAP7_75t_L g18840 ( 
.A1(n_18678),
.A2(n_18514),
.B(n_6024),
.Y(n_18840)
);

NAND2xp5_ASAP7_75t_SL g18841 ( 
.A(n_18668),
.B(n_6688),
.Y(n_18841)
);

OAI22xp33_ASAP7_75t_SL g18842 ( 
.A1(n_18778),
.A2(n_8848),
.B1(n_8855),
.B2(n_8853),
.Y(n_18842)
);

OAI221xp5_ASAP7_75t_L g18843 ( 
.A1(n_18654),
.A2(n_7671),
.B1(n_7166),
.B2(n_7142),
.C(n_8967),
.Y(n_18843)
);

OAI22xp33_ASAP7_75t_SL g18844 ( 
.A1(n_18686),
.A2(n_8853),
.B1(n_8860),
.B2(n_8855),
.Y(n_18844)
);

BUFx2_ASAP7_75t_L g18845 ( 
.A(n_18673),
.Y(n_18845)
);

NOR4xp25_ASAP7_75t_SL g18846 ( 
.A(n_18701),
.B(n_8871),
.C(n_8879),
.D(n_8860),
.Y(n_18846)
);

AOI22xp5_ASAP7_75t_L g18847 ( 
.A1(n_18710),
.A2(n_7671),
.B1(n_7081),
.B2(n_7296),
.Y(n_18847)
);

AOI211x1_ASAP7_75t_L g18848 ( 
.A1(n_18729),
.A2(n_8879),
.B(n_8883),
.C(n_8871),
.Y(n_18848)
);

NAND2xp5_ASAP7_75t_L g18849 ( 
.A(n_18824),
.B(n_8982),
.Y(n_18849)
);

NOR3xp33_ASAP7_75t_L g18850 ( 
.A(n_18657),
.B(n_5125),
.C(n_4632),
.Y(n_18850)
);

AOI211xp5_ASAP7_75t_SL g18851 ( 
.A1(n_18743),
.A2(n_5353),
.B(n_5390),
.C(n_5228),
.Y(n_18851)
);

INVx1_ASAP7_75t_L g18852 ( 
.A(n_18747),
.Y(n_18852)
);

INVx1_ASAP7_75t_L g18853 ( 
.A(n_18754),
.Y(n_18853)
);

OAI22xp5_ASAP7_75t_L g18854 ( 
.A1(n_18694),
.A2(n_7656),
.B1(n_7611),
.B2(n_8982),
.Y(n_18854)
);

INVx1_ASAP7_75t_L g18855 ( 
.A(n_18658),
.Y(n_18855)
);

AOI221xp5_ASAP7_75t_L g18856 ( 
.A1(n_18723),
.A2(n_8885),
.B1(n_8886),
.B2(n_8884),
.C(n_8883),
.Y(n_18856)
);

AOI21xp5_ASAP7_75t_L g18857 ( 
.A1(n_18655),
.A2(n_7480),
.B(n_8258),
.Y(n_18857)
);

NOR2x1_ASAP7_75t_L g18858 ( 
.A(n_18653),
.B(n_5125),
.Y(n_18858)
);

NOR2xp33_ASAP7_75t_L g18859 ( 
.A(n_18776),
.B(n_18822),
.Y(n_18859)
);

OAI21xp5_ASAP7_75t_SL g18860 ( 
.A1(n_18665),
.A2(n_5180),
.B(n_5453),
.Y(n_18860)
);

INVx1_ASAP7_75t_L g18861 ( 
.A(n_18656),
.Y(n_18861)
);

INVx2_ASAP7_75t_L g18862 ( 
.A(n_18811),
.Y(n_18862)
);

OAI21xp5_ASAP7_75t_SL g18863 ( 
.A1(n_18773),
.A2(n_5180),
.B(n_5453),
.Y(n_18863)
);

A2O1A1Ixp33_ASAP7_75t_L g18864 ( 
.A1(n_18794),
.A2(n_8240),
.B(n_8244),
.C(n_8233),
.Y(n_18864)
);

AOI21xp5_ASAP7_75t_L g18865 ( 
.A1(n_18774),
.A2(n_7480),
.B(n_8352),
.Y(n_18865)
);

INVx1_ASAP7_75t_L g18866 ( 
.A(n_18699),
.Y(n_18866)
);

AOI322xp5_ASAP7_75t_L g18867 ( 
.A1(n_18770),
.A2(n_7434),
.A3(n_7548),
.B1(n_7588),
.B2(n_7596),
.C1(n_7524),
.C2(n_7451),
.Y(n_18867)
);

OAI21xp5_ASAP7_75t_L g18868 ( 
.A1(n_18722),
.A2(n_7894),
.B(n_7885),
.Y(n_18868)
);

AND2x2_ASAP7_75t_L g18869 ( 
.A(n_18700),
.B(n_6658),
.Y(n_18869)
);

NAND2xp5_ASAP7_75t_SL g18870 ( 
.A(n_18766),
.B(n_6688),
.Y(n_18870)
);

OAI221xp5_ASAP7_75t_SL g18871 ( 
.A1(n_18650),
.A2(n_7596),
.B1(n_7608),
.B2(n_7588),
.C(n_7548),
.Y(n_18871)
);

OAI221xp5_ASAP7_75t_L g18872 ( 
.A1(n_18652),
.A2(n_7166),
.B1(n_7142),
.B2(n_8982),
.C(n_5995),
.Y(n_18872)
);

OAI22xp5_ASAP7_75t_L g18873 ( 
.A1(n_18775),
.A2(n_18777),
.B1(n_18663),
.B2(n_18661),
.Y(n_18873)
);

INVx1_ASAP7_75t_L g18874 ( 
.A(n_18651),
.Y(n_18874)
);

AOI22xp33_ASAP7_75t_L g18875 ( 
.A1(n_18725),
.A2(n_6688),
.B1(n_6733),
.B2(n_6718),
.Y(n_18875)
);

AOI22xp5_ASAP7_75t_L g18876 ( 
.A1(n_18798),
.A2(n_7081),
.B1(n_7296),
.B2(n_6942),
.Y(n_18876)
);

NAND2xp33_ASAP7_75t_R g18877 ( 
.A(n_18733),
.B(n_5228),
.Y(n_18877)
);

AOI22xp5_ASAP7_75t_L g18878 ( 
.A1(n_18801),
.A2(n_18768),
.B1(n_18763),
.B2(n_18719),
.Y(n_18878)
);

AOI22xp5_ASAP7_75t_L g18879 ( 
.A1(n_18720),
.A2(n_7081),
.B1(n_7296),
.B2(n_6942),
.Y(n_18879)
);

AOI21xp5_ASAP7_75t_L g18880 ( 
.A1(n_18670),
.A2(n_8352),
.B(n_7779),
.Y(n_18880)
);

AOI21xp33_ASAP7_75t_L g18881 ( 
.A1(n_18830),
.A2(n_6024),
.B(n_5083),
.Y(n_18881)
);

NOR3x1_ASAP7_75t_L g18882 ( 
.A(n_18806),
.B(n_7894),
.C(n_7885),
.Y(n_18882)
);

A2O1A1Ixp33_ASAP7_75t_L g18883 ( 
.A1(n_18704),
.A2(n_8244),
.B(n_8245),
.C(n_8240),
.Y(n_18883)
);

CKINVDCx20_ASAP7_75t_R g18884 ( 
.A(n_18793),
.Y(n_18884)
);

INVxp67_ASAP7_75t_L g18885 ( 
.A(n_18790),
.Y(n_18885)
);

OAI311xp33_ASAP7_75t_L g18886 ( 
.A1(n_18703),
.A2(n_18708),
.A3(n_18717),
.B1(n_18724),
.C1(n_18711),
.Y(n_18886)
);

AOI22xp5_ASAP7_75t_L g18887 ( 
.A1(n_18788),
.A2(n_7296),
.B1(n_7298),
.B2(n_6942),
.Y(n_18887)
);

BUFx2_ASAP7_75t_L g18888 ( 
.A(n_18751),
.Y(n_18888)
);

AOI32xp33_ASAP7_75t_L g18889 ( 
.A1(n_18681),
.A2(n_7298),
.A3(n_7342),
.B1(n_7296),
.B2(n_6942),
.Y(n_18889)
);

OAI21xp33_ASAP7_75t_L g18890 ( 
.A1(n_18792),
.A2(n_7298),
.B(n_6942),
.Y(n_18890)
);

OAI221xp5_ASAP7_75t_SL g18891 ( 
.A1(n_18799),
.A2(n_18742),
.B1(n_18721),
.B2(n_18713),
.C(n_18680),
.Y(n_18891)
);

AOI221xp5_ASAP7_75t_L g18892 ( 
.A1(n_18816),
.A2(n_8886),
.B1(n_8890),
.B2(n_8885),
.C(n_8884),
.Y(n_18892)
);

AOI32xp33_ASAP7_75t_L g18893 ( 
.A1(n_18677),
.A2(n_7510),
.A3(n_7569),
.B1(n_7342),
.B2(n_7298),
.Y(n_18893)
);

AOI221xp5_ASAP7_75t_L g18894 ( 
.A1(n_18789),
.A2(n_8902),
.B1(n_8908),
.B2(n_8900),
.C(n_8890),
.Y(n_18894)
);

AOI221x1_ASAP7_75t_L g18895 ( 
.A1(n_18707),
.A2(n_8908),
.B1(n_8909),
.B2(n_8902),
.C(n_8900),
.Y(n_18895)
);

INVx1_ASAP7_75t_L g18896 ( 
.A(n_18688),
.Y(n_18896)
);

OAI322xp33_ASAP7_75t_L g18897 ( 
.A1(n_18746),
.A2(n_8949),
.A3(n_8932),
.B1(n_8951),
.B2(n_8960),
.C1(n_8936),
.C2(n_8909),
.Y(n_18897)
);

OAI22xp5_ASAP7_75t_L g18898 ( 
.A1(n_18689),
.A2(n_7320),
.B1(n_7363),
.B2(n_7285),
.Y(n_18898)
);

AOI21xp5_ASAP7_75t_L g18899 ( 
.A1(n_18809),
.A2(n_8352),
.B(n_7779),
.Y(n_18899)
);

OAI21xp33_ASAP7_75t_L g18900 ( 
.A1(n_18674),
.A2(n_7342),
.B(n_7298),
.Y(n_18900)
);

AOI322xp5_ASAP7_75t_L g18901 ( 
.A1(n_18817),
.A2(n_18821),
.A3(n_18738),
.B1(n_18827),
.B2(n_18750),
.C1(n_18755),
.C2(n_18682),
.Y(n_18901)
);

AOI31xp33_ASAP7_75t_L g18902 ( 
.A1(n_18753),
.A2(n_18797),
.A3(n_18805),
.B(n_18739),
.Y(n_18902)
);

INVx2_ASAP7_75t_L g18903 ( 
.A(n_18662),
.Y(n_18903)
);

AOI22xp5_ASAP7_75t_L g18904 ( 
.A1(n_18779),
.A2(n_7510),
.B1(n_7569),
.B2(n_7342),
.Y(n_18904)
);

AOI221xp5_ASAP7_75t_L g18905 ( 
.A1(n_18726),
.A2(n_18741),
.B1(n_18813),
.B2(n_18709),
.C(n_18734),
.Y(n_18905)
);

NAND2xp5_ASAP7_75t_L g18906 ( 
.A(n_18823),
.B(n_8352),
.Y(n_18906)
);

INVx1_ASAP7_75t_L g18907 ( 
.A(n_18812),
.Y(n_18907)
);

NAND2xp5_ASAP7_75t_L g18908 ( 
.A(n_18679),
.B(n_8352),
.Y(n_18908)
);

AOI221x1_ASAP7_75t_L g18909 ( 
.A1(n_18786),
.A2(n_8949),
.B1(n_8951),
.B2(n_8936),
.C(n_8932),
.Y(n_18909)
);

INVx1_ASAP7_75t_L g18910 ( 
.A(n_18685),
.Y(n_18910)
);

INVx1_ASAP7_75t_L g18911 ( 
.A(n_18698),
.Y(n_18911)
);

INVx1_ASAP7_75t_L g18912 ( 
.A(n_18820),
.Y(n_18912)
);

XNOR2xp5_ASAP7_75t_L g18913 ( 
.A(n_18671),
.B(n_6911),
.Y(n_18913)
);

AOI221xp5_ASAP7_75t_L g18914 ( 
.A1(n_18756),
.A2(n_8971),
.B1(n_8987),
.B2(n_8968),
.C(n_8960),
.Y(n_18914)
);

OAI21xp33_ASAP7_75t_SL g18915 ( 
.A1(n_18785),
.A2(n_8244),
.B(n_8240),
.Y(n_18915)
);

INVx1_ASAP7_75t_L g18916 ( 
.A(n_18745),
.Y(n_18916)
);

NAND2xp5_ASAP7_75t_L g18917 ( 
.A(n_18715),
.B(n_18764),
.Y(n_18917)
);

NOR2x1_ASAP7_75t_L g18918 ( 
.A(n_18810),
.B(n_5125),
.Y(n_18918)
);

INVx1_ASAP7_75t_L g18919 ( 
.A(n_18705),
.Y(n_18919)
);

BUFx2_ASAP7_75t_L g18920 ( 
.A(n_18684),
.Y(n_18920)
);

AOI221xp5_ASAP7_75t_L g18921 ( 
.A1(n_18718),
.A2(n_18675),
.B1(n_18772),
.B2(n_18828),
.C(n_18762),
.Y(n_18921)
);

INVx2_ASAP7_75t_L g18922 ( 
.A(n_18769),
.Y(n_18922)
);

O2A1O1Ixp33_ASAP7_75t_L g18923 ( 
.A1(n_18803),
.A2(n_4632),
.B(n_4647),
.C(n_4601),
.Y(n_18923)
);

OAI21xp33_ASAP7_75t_SL g18924 ( 
.A1(n_18669),
.A2(n_8247),
.B(n_8245),
.Y(n_18924)
);

INVx1_ASAP7_75t_L g18925 ( 
.A(n_18780),
.Y(n_18925)
);

O2A1O1Ixp33_ASAP7_75t_L g18926 ( 
.A1(n_18784),
.A2(n_4632),
.B(n_4683),
.C(n_4647),
.Y(n_18926)
);

AOI21xp5_ASAP7_75t_L g18927 ( 
.A1(n_18692),
.A2(n_7779),
.B(n_7686),
.Y(n_18927)
);

OAI21xp33_ASAP7_75t_L g18928 ( 
.A1(n_18783),
.A2(n_7510),
.B(n_7342),
.Y(n_18928)
);

OAI322xp33_ASAP7_75t_L g18929 ( 
.A1(n_18693),
.A2(n_8998),
.A3(n_8971),
.B1(n_8999),
.B2(n_9005),
.C1(n_8987),
.C2(n_8968),
.Y(n_18929)
);

INVx1_ASAP7_75t_L g18930 ( 
.A(n_18807),
.Y(n_18930)
);

OAI211xp5_ASAP7_75t_L g18931 ( 
.A1(n_18728),
.A2(n_5125),
.B(n_7363),
.C(n_7320),
.Y(n_18931)
);

INVx2_ASAP7_75t_L g18932 ( 
.A(n_18814),
.Y(n_18932)
);

OAI21xp5_ASAP7_75t_L g18933 ( 
.A1(n_18752),
.A2(n_7895),
.B(n_8245),
.Y(n_18933)
);

OR2x2_ASAP7_75t_L g18934 ( 
.A(n_18749),
.B(n_8790),
.Y(n_18934)
);

AOI22xp5_ASAP7_75t_L g18935 ( 
.A1(n_18702),
.A2(n_7569),
.B1(n_7680),
.B2(n_7510),
.Y(n_18935)
);

INVx2_ASAP7_75t_L g18936 ( 
.A(n_18691),
.Y(n_18936)
);

INVx1_ASAP7_75t_L g18937 ( 
.A(n_18765),
.Y(n_18937)
);

INVx1_ASAP7_75t_SL g18938 ( 
.A(n_18676),
.Y(n_18938)
);

AOI21xp5_ASAP7_75t_L g18939 ( 
.A1(n_18736),
.A2(n_18735),
.B(n_18791),
.Y(n_18939)
);

AOI221xp5_ASAP7_75t_L g18940 ( 
.A1(n_18697),
.A2(n_9005),
.B1(n_9013),
.B2(n_8999),
.C(n_8998),
.Y(n_18940)
);

AOI211x1_ASAP7_75t_SL g18941 ( 
.A1(n_18795),
.A2(n_6718),
.B(n_6733),
.C(n_6688),
.Y(n_18941)
);

INVxp67_ASAP7_75t_L g18942 ( 
.A(n_18815),
.Y(n_18942)
);

NOR2xp33_ASAP7_75t_SL g18943 ( 
.A(n_18829),
.B(n_5180),
.Y(n_18943)
);

O2A1O1Ixp33_ASAP7_75t_L g18944 ( 
.A1(n_18781),
.A2(n_4647),
.B(n_4683),
.C(n_4957),
.Y(n_18944)
);

OAI211xp5_ASAP7_75t_L g18945 ( 
.A1(n_18800),
.A2(n_7372),
.B(n_7467),
.C(n_7368),
.Y(n_18945)
);

INVx2_ASAP7_75t_L g18946 ( 
.A(n_18691),
.Y(n_18946)
);

NAND3xp33_ASAP7_75t_L g18947 ( 
.A(n_18716),
.B(n_7372),
.C(n_7368),
.Y(n_18947)
);

INVx2_ASAP7_75t_L g18948 ( 
.A(n_18782),
.Y(n_18948)
);

NOR2x1_ASAP7_75t_L g18949 ( 
.A(n_18808),
.B(n_8320),
.Y(n_18949)
);

OAI22xp5_ASAP7_75t_L g18950 ( 
.A1(n_18760),
.A2(n_7576),
.B1(n_7652),
.B2(n_7467),
.Y(n_18950)
);

OAI21xp5_ASAP7_75t_SL g18951 ( 
.A1(n_18732),
.A2(n_5459),
.B(n_5453),
.Y(n_18951)
);

XOR2x2_ASAP7_75t_L g18952 ( 
.A(n_18667),
.B(n_5871),
.Y(n_18952)
);

INVxp67_ASAP7_75t_L g18953 ( 
.A(n_18804),
.Y(n_18953)
);

NAND2xp5_ASAP7_75t_L g18954 ( 
.A(n_18696),
.B(n_18796),
.Y(n_18954)
);

XNOR2x1_ASAP7_75t_L g18955 ( 
.A(n_18826),
.B(n_7895),
.Y(n_18955)
);

NAND2xp33_ASAP7_75t_R g18956 ( 
.A(n_18712),
.B(n_5228),
.Y(n_18956)
);

AOI22xp5_ASAP7_75t_L g18957 ( 
.A1(n_18802),
.A2(n_18818),
.B1(n_18748),
.B2(n_18767),
.Y(n_18957)
);

AOI22xp5_ASAP7_75t_L g18958 ( 
.A1(n_18758),
.A2(n_7569),
.B1(n_7680),
.B2(n_7510),
.Y(n_18958)
);

A2O1A1Ixp33_ASAP7_75t_L g18959 ( 
.A1(n_18771),
.A2(n_8250),
.B(n_8252),
.C(n_8247),
.Y(n_18959)
);

O2A1O1Ixp33_ASAP7_75t_L g18960 ( 
.A1(n_18730),
.A2(n_4683),
.B(n_5011),
.C(n_4957),
.Y(n_18960)
);

NAND3xp33_ASAP7_75t_SL g18961 ( 
.A(n_18787),
.B(n_5553),
.C(n_5541),
.Y(n_18961)
);

INVx1_ASAP7_75t_SL g18962 ( 
.A(n_18695),
.Y(n_18962)
);

OAI21xp33_ASAP7_75t_SL g18963 ( 
.A1(n_18737),
.A2(n_8250),
.B(n_8247),
.Y(n_18963)
);

OAI21xp33_ASAP7_75t_L g18964 ( 
.A1(n_18731),
.A2(n_7569),
.B(n_7510),
.Y(n_18964)
);

INVx3_ASAP7_75t_L g18965 ( 
.A(n_18672),
.Y(n_18965)
);

INVx1_ASAP7_75t_L g18966 ( 
.A(n_18727),
.Y(n_18966)
);

INVx2_ASAP7_75t_L g18967 ( 
.A(n_18825),
.Y(n_18967)
);

NOR2x1_ASAP7_75t_L g18968 ( 
.A(n_18660),
.B(n_8188),
.Y(n_18968)
);

INVx2_ASAP7_75t_L g18969 ( 
.A(n_18740),
.Y(n_18969)
);

OAI22xp5_ASAP7_75t_L g18970 ( 
.A1(n_18714),
.A2(n_7652),
.B1(n_7659),
.B2(n_7576),
.Y(n_18970)
);

INVxp67_ASAP7_75t_L g18971 ( 
.A(n_18664),
.Y(n_18971)
);

NOR3xp33_ASAP7_75t_L g18972 ( 
.A(n_18714),
.B(n_5353),
.C(n_5228),
.Y(n_18972)
);

AOI21xp5_ASAP7_75t_L g18973 ( 
.A1(n_18666),
.A2(n_7686),
.B(n_7780),
.Y(n_18973)
);

OAI22xp33_ASAP7_75t_L g18974 ( 
.A1(n_18714),
.A2(n_7254),
.B1(n_7262),
.B2(n_7225),
.Y(n_18974)
);

OAI21xp5_ASAP7_75t_L g18975 ( 
.A1(n_18659),
.A2(n_7895),
.B(n_8250),
.Y(n_18975)
);

AOI22xp5_ASAP7_75t_L g18976 ( 
.A1(n_18714),
.A2(n_7680),
.B1(n_7569),
.B2(n_7608),
.Y(n_18976)
);

AOI221xp5_ASAP7_75t_L g18977 ( 
.A1(n_18664),
.A2(n_9023),
.B1(n_9031),
.B2(n_9016),
.C(n_9013),
.Y(n_18977)
);

OAI221xp5_ASAP7_75t_SL g18978 ( 
.A1(n_18687),
.A2(n_7673),
.B1(n_7608),
.B2(n_7596),
.C(n_7215),
.Y(n_18978)
);

AOI221xp5_ASAP7_75t_L g18979 ( 
.A1(n_18664),
.A2(n_9023),
.B1(n_9021),
.B2(n_9016),
.C(n_9031),
.Y(n_18979)
);

AOI22xp33_ASAP7_75t_SL g18980 ( 
.A1(n_18714),
.A2(n_6688),
.B1(n_6733),
.B2(n_6718),
.Y(n_18980)
);

OAI221xp5_ASAP7_75t_L g18981 ( 
.A1(n_18971),
.A2(n_5033),
.B1(n_5112),
.B2(n_5050),
.C(n_5011),
.Y(n_18981)
);

OAI21xp33_ASAP7_75t_SL g18982 ( 
.A1(n_18968),
.A2(n_8256),
.B(n_8252),
.Y(n_18982)
);

AOI221xp5_ASAP7_75t_L g18983 ( 
.A1(n_18833),
.A2(n_9021),
.B1(n_7682),
.B2(n_7696),
.C(n_7659),
.Y(n_18983)
);

AO211x2_ASAP7_75t_L g18984 ( 
.A1(n_18835),
.A2(n_7208),
.B(n_7237),
.C(n_7232),
.Y(n_18984)
);

AOI21xp5_ASAP7_75t_L g18985 ( 
.A1(n_18838),
.A2(n_7781),
.B(n_7780),
.Y(n_18985)
);

NAND2xp33_ASAP7_75t_R g18986 ( 
.A(n_18845),
.B(n_5353),
.Y(n_18986)
);

AOI321xp33_ASAP7_75t_L g18987 ( 
.A1(n_18873),
.A2(n_7680),
.A3(n_6916),
.B1(n_7037),
.B2(n_7087),
.C(n_7085),
.Y(n_18987)
);

NAND2xp33_ASAP7_75t_SL g18988 ( 
.A(n_18837),
.B(n_5459),
.Y(n_18988)
);

AOI221xp5_ASAP7_75t_L g18989 ( 
.A1(n_18834),
.A2(n_7682),
.B1(n_7696),
.B2(n_7680),
.C(n_7221),
.Y(n_18989)
);

OAI211xp5_ASAP7_75t_SL g18990 ( 
.A1(n_18901),
.A2(n_5390),
.B(n_5452),
.C(n_5353),
.Y(n_18990)
);

NOR2x1_ASAP7_75t_L g18991 ( 
.A(n_18836),
.B(n_5984),
.Y(n_18991)
);

INVx1_ASAP7_75t_L g18992 ( 
.A(n_18849),
.Y(n_18992)
);

OAI321xp33_ASAP7_75t_L g18993 ( 
.A1(n_18885),
.A2(n_6772),
.A3(n_6688),
.B1(n_6785),
.B2(n_6733),
.C(n_6718),
.Y(n_18993)
);

BUFx3_ASAP7_75t_L g18994 ( 
.A(n_18930),
.Y(n_18994)
);

AOI22xp33_ASAP7_75t_L g18995 ( 
.A1(n_18896),
.A2(n_6688),
.B1(n_6733),
.B2(n_6718),
.Y(n_18995)
);

AOI221xp5_ASAP7_75t_L g18996 ( 
.A1(n_18840),
.A2(n_7680),
.B1(n_7221),
.B2(n_7282),
.C(n_7019),
.Y(n_18996)
);

AOI22xp5_ASAP7_75t_L g18997 ( 
.A1(n_18859),
.A2(n_7673),
.B1(n_6718),
.B2(n_6733),
.Y(n_18997)
);

INVx1_ASAP7_75t_L g18998 ( 
.A(n_18869),
.Y(n_18998)
);

OAI21xp33_ASAP7_75t_L g18999 ( 
.A1(n_18853),
.A2(n_7242),
.B(n_7215),
.Y(n_18999)
);

AOI22xp33_ASAP7_75t_L g19000 ( 
.A1(n_18855),
.A2(n_6688),
.B1(n_6733),
.B2(n_6718),
.Y(n_19000)
);

OAI22xp5_ASAP7_75t_L g19001 ( 
.A1(n_18861),
.A2(n_7673),
.B1(n_6718),
.B2(n_6733),
.Y(n_19001)
);

AOI221xp5_ASAP7_75t_L g19002 ( 
.A1(n_18902),
.A2(n_18966),
.B1(n_18907),
.B2(n_18962),
.C(n_18874),
.Y(n_19002)
);

AOI211xp5_ASAP7_75t_L g19003 ( 
.A1(n_18886),
.A2(n_18891),
.B(n_18912),
.C(n_18919),
.Y(n_19003)
);

O2A1O1Ixp33_ASAP7_75t_L g19004 ( 
.A1(n_18831),
.A2(n_5050),
.B(n_5112),
.C(n_5033),
.Y(n_19004)
);

OAI221xp5_ASAP7_75t_L g19005 ( 
.A1(n_18878),
.A2(n_5050),
.B1(n_5112),
.B2(n_5033),
.C(n_7142),
.Y(n_19005)
);

OAI221xp5_ASAP7_75t_L g19006 ( 
.A1(n_18921),
.A2(n_7166),
.B1(n_7142),
.B2(n_5995),
.C(n_5917),
.Y(n_19006)
);

AOI221xp5_ASAP7_75t_L g19007 ( 
.A1(n_18965),
.A2(n_18852),
.B1(n_18870),
.B2(n_18841),
.C(n_18938),
.Y(n_19007)
);

AOI21xp5_ASAP7_75t_L g19008 ( 
.A1(n_18920),
.A2(n_7781),
.B(n_7780),
.Y(n_19008)
);

AOI322xp5_ASAP7_75t_L g19009 ( 
.A1(n_18937),
.A2(n_7242),
.A3(n_7245),
.B1(n_7257),
.B2(n_7014),
.C1(n_6981),
.C2(n_7158),
.Y(n_19009)
);

OAI21xp5_ASAP7_75t_L g19010 ( 
.A1(n_18942),
.A2(n_8578),
.B(n_8571),
.Y(n_19010)
);

AOI21xp5_ASAP7_75t_SL g19011 ( 
.A1(n_18862),
.A2(n_5960),
.B(n_5891),
.Y(n_19011)
);

NOR2x1p5_ASAP7_75t_L g19012 ( 
.A(n_18965),
.B(n_5453),
.Y(n_19012)
);

AOI22xp5_ASAP7_75t_L g19013 ( 
.A1(n_18884),
.A2(n_6718),
.B1(n_6733),
.B2(n_6688),
.Y(n_19013)
);

A2O1A1Ixp33_ASAP7_75t_L g19014 ( 
.A1(n_18903),
.A2(n_8256),
.B(n_8262),
.C(n_8252),
.Y(n_19014)
);

XNOR2xp5_ASAP7_75t_L g19015 ( 
.A(n_18832),
.B(n_4472),
.Y(n_19015)
);

NOR2xp33_ASAP7_75t_R g19016 ( 
.A(n_18888),
.B(n_6157),
.Y(n_19016)
);

NOR2x1_ASAP7_75t_L g19017 ( 
.A(n_18858),
.B(n_18936),
.Y(n_19017)
);

AOI221xp5_ASAP7_75t_L g19018 ( 
.A1(n_18905),
.A2(n_7431),
.B1(n_7437),
.B2(n_7019),
.C(n_6833),
.Y(n_19018)
);

CKINVDCx16_ASAP7_75t_R g19019 ( 
.A(n_18925),
.Y(n_19019)
);

OAI211xp5_ASAP7_75t_L g19020 ( 
.A1(n_18953),
.A2(n_18839),
.B(n_18916),
.C(n_18948),
.Y(n_19020)
);

OAI211xp5_ASAP7_75t_L g19021 ( 
.A1(n_18910),
.A2(n_5459),
.B(n_5484),
.C(n_5453),
.Y(n_19021)
);

OAI211xp5_ASAP7_75t_SL g19022 ( 
.A1(n_18866),
.A2(n_18911),
.B(n_18969),
.C(n_18932),
.Y(n_19022)
);

AOI211xp5_ASAP7_75t_SL g19023 ( 
.A1(n_18881),
.A2(n_5390),
.B(n_5452),
.C(n_5353),
.Y(n_19023)
);

AOI21xp33_ASAP7_75t_L g19024 ( 
.A1(n_18917),
.A2(n_5459),
.B(n_5453),
.Y(n_19024)
);

INVx2_ASAP7_75t_SL g19025 ( 
.A(n_18922),
.Y(n_19025)
);

INVx1_ASAP7_75t_SL g19026 ( 
.A(n_18967),
.Y(n_19026)
);

O2A1O1Ixp33_ASAP7_75t_SL g19027 ( 
.A1(n_18946),
.A2(n_7014),
.B(n_6981),
.C(n_7128),
.Y(n_19027)
);

NAND4xp75_ASAP7_75t_L g19028 ( 
.A(n_18918),
.B(n_7715),
.C(n_7336),
.D(n_7501),
.Y(n_19028)
);

NOR2xp67_ASAP7_75t_L g19029 ( 
.A(n_18957),
.B(n_5453),
.Y(n_19029)
);

AOI221xp5_ASAP7_75t_L g19030 ( 
.A1(n_18872),
.A2(n_7366),
.B1(n_7527),
.B2(n_7136),
.C(n_6941),
.Y(n_19030)
);

NOR2x1_ASAP7_75t_L g19031 ( 
.A(n_18954),
.B(n_5984),
.Y(n_19031)
);

INVx1_ASAP7_75t_L g19032 ( 
.A(n_18939),
.Y(n_19032)
);

OAI211xp5_ASAP7_75t_L g19033 ( 
.A1(n_18951),
.A2(n_5484),
.B(n_5489),
.C(n_5459),
.Y(n_19033)
);

AOI222xp33_ASAP7_75t_L g19034 ( 
.A1(n_18961),
.A2(n_6575),
.B1(n_5960),
.B2(n_6916),
.C1(n_7037),
.C2(n_6969),
.Y(n_19034)
);

AOI221xp5_ASAP7_75t_L g19035 ( 
.A1(n_18973),
.A2(n_7141),
.B1(n_7206),
.B2(n_6989),
.C(n_6951),
.Y(n_19035)
);

AOI31xp33_ASAP7_75t_L g19036 ( 
.A1(n_18877),
.A2(n_7134),
.A3(n_7145),
.B(n_7128),
.Y(n_19036)
);

AND2x2_ASAP7_75t_L g19037 ( 
.A(n_18913),
.B(n_18972),
.Y(n_19037)
);

AOI22xp33_ASAP7_75t_L g19038 ( 
.A1(n_18850),
.A2(n_6772),
.B1(n_6806),
.B2(n_6785),
.Y(n_19038)
);

O2A1O1Ixp5_ASAP7_75t_L g19039 ( 
.A1(n_18871),
.A2(n_7564),
.B(n_7166),
.C(n_7142),
.Y(n_19039)
);

AOI221xp5_ASAP7_75t_L g19040 ( 
.A1(n_18842),
.A2(n_7141),
.B1(n_7206),
.B2(n_6989),
.C(n_6951),
.Y(n_19040)
);

XNOR2x2_ASAP7_75t_L g19041 ( 
.A(n_18952),
.B(n_8256),
.Y(n_19041)
);

NOR3xp33_ASAP7_75t_L g19042 ( 
.A(n_18945),
.B(n_5452),
.C(n_5390),
.Y(n_19042)
);

AOI221xp5_ASAP7_75t_L g19043 ( 
.A1(n_18844),
.A2(n_18944),
.B1(n_18863),
.B2(n_18960),
.C(n_18860),
.Y(n_19043)
);

OAI21xp5_ASAP7_75t_L g19044 ( 
.A1(n_18927),
.A2(n_8578),
.B(n_8571),
.Y(n_19044)
);

OAI21xp5_ASAP7_75t_L g19045 ( 
.A1(n_18949),
.A2(n_8578),
.B(n_8571),
.Y(n_19045)
);

INVx1_ASAP7_75t_SL g19046 ( 
.A(n_18943),
.Y(n_19046)
);

OAI21xp33_ASAP7_75t_SL g19047 ( 
.A1(n_18875),
.A2(n_8266),
.B(n_8262),
.Y(n_19047)
);

A2O1A1Ixp33_ASAP7_75t_L g19048 ( 
.A1(n_18947),
.A2(n_18931),
.B(n_18963),
.C(n_18923),
.Y(n_19048)
);

INVx1_ASAP7_75t_L g19049 ( 
.A(n_18941),
.Y(n_19049)
);

NOR3xp33_ASAP7_75t_L g19050 ( 
.A(n_18978),
.B(n_5452),
.C(n_5390),
.Y(n_19050)
);

OR2x2_ASAP7_75t_L g19051 ( 
.A(n_18970),
.B(n_8790),
.Y(n_19051)
);

OAI21xp5_ASAP7_75t_L g19052 ( 
.A1(n_18854),
.A2(n_8597),
.B(n_8591),
.Y(n_19052)
);

AOI322xp5_ASAP7_75t_L g19053 ( 
.A1(n_18890),
.A2(n_7245),
.A3(n_7257),
.B1(n_7242),
.B2(n_7014),
.C1(n_6981),
.C2(n_7110),
.Y(n_19053)
);

AOI221xp5_ASAP7_75t_L g19054 ( 
.A1(n_18950),
.A2(n_7169),
.B1(n_7221),
.B2(n_7094),
.C(n_6785),
.Y(n_19054)
);

OAI22xp33_ASAP7_75t_L g19055 ( 
.A1(n_18976),
.A2(n_18956),
.B1(n_18906),
.B2(n_18851),
.Y(n_19055)
);

O2A1O1Ixp33_ASAP7_75t_L g19056 ( 
.A1(n_18908),
.A2(n_5452),
.B(n_5917),
.C(n_5871),
.Y(n_19056)
);

INVx1_ASAP7_75t_L g19057 ( 
.A(n_18848),
.Y(n_19057)
);

NAND2xp5_ASAP7_75t_SL g19058 ( 
.A(n_18980),
.B(n_6772),
.Y(n_19058)
);

OAI22xp5_ASAP7_75t_L g19059 ( 
.A1(n_18934),
.A2(n_6785),
.B1(n_6806),
.B2(n_6772),
.Y(n_19059)
);

OAI211xp5_ASAP7_75t_SL g19060 ( 
.A1(n_18926),
.A2(n_5282),
.B(n_5288),
.C(n_5244),
.Y(n_19060)
);

OAI22xp33_ASAP7_75t_L g19061 ( 
.A1(n_18843),
.A2(n_7254),
.B1(n_7262),
.B2(n_7225),
.Y(n_19061)
);

NOR3xp33_ASAP7_75t_SL g19062 ( 
.A(n_18898),
.B(n_7208),
.C(n_7134),
.Y(n_19062)
);

AND2x2_ASAP7_75t_L g19063 ( 
.A(n_18846),
.B(n_6658),
.Y(n_19063)
);

INVx1_ASAP7_75t_SL g19064 ( 
.A(n_18955),
.Y(n_19064)
);

AOI21xp5_ASAP7_75t_L g19065 ( 
.A1(n_18975),
.A2(n_7781),
.B(n_8262),
.Y(n_19065)
);

AOI221xp5_ASAP7_75t_L g19066 ( 
.A1(n_18929),
.A2(n_7527),
.B1(n_7535),
.B2(n_7366),
.C(n_7019),
.Y(n_19066)
);

AOI211xp5_ASAP7_75t_L g19067 ( 
.A1(n_18924),
.A2(n_5484),
.B(n_5489),
.C(n_5459),
.Y(n_19067)
);

AOI22xp5_ASAP7_75t_L g19068 ( 
.A1(n_18900),
.A2(n_18915),
.B1(n_18964),
.B2(n_18928),
.Y(n_19068)
);

OAI221xp5_ASAP7_75t_L g19069 ( 
.A1(n_18894),
.A2(n_7166),
.B1(n_7142),
.B2(n_5995),
.C(n_5917),
.Y(n_19069)
);

INVx1_ASAP7_75t_L g19070 ( 
.A(n_18909),
.Y(n_19070)
);

NOR2xp33_ASAP7_75t_L g19071 ( 
.A(n_18879),
.B(n_5459),
.Y(n_19071)
);

INVx1_ASAP7_75t_SL g19072 ( 
.A(n_18865),
.Y(n_19072)
);

OAI22xp5_ASAP7_75t_L g19073 ( 
.A1(n_18958),
.A2(n_6785),
.B1(n_6806),
.B2(n_6772),
.Y(n_19073)
);

OAI221xp5_ASAP7_75t_L g19074 ( 
.A1(n_18856),
.A2(n_7166),
.B1(n_5995),
.B2(n_5917),
.C(n_5871),
.Y(n_19074)
);

AOI221xp5_ASAP7_75t_L g19075 ( 
.A1(n_18977),
.A2(n_6772),
.B1(n_7282),
.B2(n_6844),
.C(n_6806),
.Y(n_19075)
);

AOI21xp33_ASAP7_75t_L g19076 ( 
.A1(n_18974),
.A2(n_5484),
.B(n_5459),
.Y(n_19076)
);

AOI31xp33_ASAP7_75t_L g19077 ( 
.A1(n_18979),
.A2(n_18892),
.A3(n_18857),
.B(n_18876),
.Y(n_19077)
);

OAI21xp33_ASAP7_75t_L g19078 ( 
.A1(n_18867),
.A2(n_7257),
.B(n_7245),
.Y(n_19078)
);

NOR3xp33_ASAP7_75t_L g19079 ( 
.A(n_18897),
.B(n_18864),
.C(n_18914),
.Y(n_19079)
);

OAI222xp33_ASAP7_75t_L g19080 ( 
.A1(n_18847),
.A2(n_7254),
.B1(n_7303),
.B2(n_7429),
.C1(n_7306),
.C2(n_7225),
.Y(n_19080)
);

OAI211xp5_ASAP7_75t_SL g19081 ( 
.A1(n_18933),
.A2(n_5282),
.B(n_5288),
.C(n_5244),
.Y(n_19081)
);

OAI21xp33_ASAP7_75t_L g19082 ( 
.A1(n_18887),
.A2(n_7505),
.B(n_7504),
.Y(n_19082)
);

O2A1O1Ixp33_ASAP7_75t_L g19083 ( 
.A1(n_18959),
.A2(n_5282),
.B(n_5288),
.C(n_5244),
.Y(n_19083)
);

AOI21xp33_ASAP7_75t_L g19084 ( 
.A1(n_18904),
.A2(n_5484),
.B(n_5459),
.Y(n_19084)
);

AOI22xp5_ASAP7_75t_SL g19085 ( 
.A1(n_18899),
.A2(n_4748),
.B1(n_4608),
.B2(n_5484),
.Y(n_19085)
);

AOI211xp5_ASAP7_75t_L g19086 ( 
.A1(n_18868),
.A2(n_18940),
.B(n_18883),
.C(n_18880),
.Y(n_19086)
);

O2A1O1Ixp33_ASAP7_75t_L g19087 ( 
.A1(n_18882),
.A2(n_5282),
.B(n_5288),
.C(n_5244),
.Y(n_19087)
);

OAI221xp5_ASAP7_75t_L g19088 ( 
.A1(n_18889),
.A2(n_7564),
.B1(n_7508),
.B2(n_7521),
.C(n_7505),
.Y(n_19088)
);

INVx1_ASAP7_75t_L g19089 ( 
.A(n_18895),
.Y(n_19089)
);

AOI21xp5_ASAP7_75t_L g19090 ( 
.A1(n_18935),
.A2(n_18893),
.B(n_8271),
.Y(n_19090)
);

AND2x2_ASAP7_75t_L g19091 ( 
.A(n_18869),
.B(n_6658),
.Y(n_19091)
);

NAND2xp5_ASAP7_75t_SL g19092 ( 
.A(n_18833),
.B(n_6772),
.Y(n_19092)
);

NOR3xp33_ASAP7_75t_L g19093 ( 
.A(n_18833),
.B(n_5282),
.C(n_5244),
.Y(n_19093)
);

NAND4xp25_ASAP7_75t_L g19094 ( 
.A(n_18833),
.B(n_7505),
.C(n_7508),
.D(n_7504),
.Y(n_19094)
);

OAI211xp5_ASAP7_75t_SL g19095 ( 
.A1(n_18971),
.A2(n_5282),
.B(n_5288),
.C(n_5244),
.Y(n_19095)
);

AOI22xp5_ASAP7_75t_L g19096 ( 
.A1(n_18859),
.A2(n_6772),
.B1(n_6806),
.B2(n_6785),
.Y(n_19096)
);

XNOR2x1_ASAP7_75t_SL g19097 ( 
.A(n_18837),
.B(n_5288),
.Y(n_19097)
);

AOI221xp5_ASAP7_75t_L g19098 ( 
.A1(n_18971),
.A2(n_7453),
.B1(n_7492),
.B2(n_7094),
.C(n_6785),
.Y(n_19098)
);

AOI221x1_ASAP7_75t_L g19099 ( 
.A1(n_18855),
.A2(n_7110),
.B1(n_7132),
.B2(n_7106),
.C(n_7057),
.Y(n_19099)
);

NAND3xp33_ASAP7_75t_L g19100 ( 
.A(n_18971),
.B(n_5489),
.C(n_5484),
.Y(n_19100)
);

O2A1O1Ixp33_ASAP7_75t_L g19101 ( 
.A1(n_18971),
.A2(n_5403),
.B(n_5411),
.C(n_5323),
.Y(n_19101)
);

AOI21xp5_ASAP7_75t_L g19102 ( 
.A1(n_18971),
.A2(n_8271),
.B(n_8266),
.Y(n_19102)
);

AOI22xp33_ASAP7_75t_L g19103 ( 
.A1(n_18837),
.A2(n_6772),
.B1(n_6806),
.B2(n_6785),
.Y(n_19103)
);

NAND2xp5_ASAP7_75t_L g19104 ( 
.A(n_18837),
.B(n_7997),
.Y(n_19104)
);

NAND3xp33_ASAP7_75t_SL g19105 ( 
.A(n_18833),
.B(n_5564),
.C(n_5553),
.Y(n_19105)
);

AOI221xp5_ASAP7_75t_L g19106 ( 
.A1(n_18971),
.A2(n_7586),
.B1(n_7657),
.B2(n_7147),
.C(n_7019),
.Y(n_19106)
);

AOI221xp5_ASAP7_75t_L g19107 ( 
.A1(n_18971),
.A2(n_7586),
.B1(n_7657),
.B2(n_7147),
.C(n_7019),
.Y(n_19107)
);

AO221x1_ASAP7_75t_L g19108 ( 
.A1(n_18971),
.A2(n_6785),
.B1(n_6844),
.B2(n_6833),
.C(n_6806),
.Y(n_19108)
);

OAI21xp33_ASAP7_75t_SL g19109 ( 
.A1(n_18968),
.A2(n_8271),
.B(n_8266),
.Y(n_19109)
);

AOI221xp5_ASAP7_75t_L g19110 ( 
.A1(n_18971),
.A2(n_7175),
.B1(n_7282),
.B2(n_7073),
.C(n_6936),
.Y(n_19110)
);

AOI221xp5_ASAP7_75t_L g19111 ( 
.A1(n_18971),
.A2(n_7175),
.B1(n_7282),
.B2(n_7073),
.C(n_6936),
.Y(n_19111)
);

INVxp67_ASAP7_75t_SL g19112 ( 
.A(n_18971),
.Y(n_19112)
);

NAND2xp5_ASAP7_75t_L g19113 ( 
.A(n_18837),
.B(n_7997),
.Y(n_19113)
);

OAI221xp5_ASAP7_75t_L g19114 ( 
.A1(n_18971),
.A2(n_7564),
.B1(n_7526),
.B2(n_7532),
.C(n_7521),
.Y(n_19114)
);

NAND4xp25_ASAP7_75t_L g19115 ( 
.A(n_18833),
.B(n_7521),
.C(n_7526),
.D(n_7508),
.Y(n_19115)
);

AOI221xp5_ASAP7_75t_L g19116 ( 
.A1(n_18971),
.A2(n_7175),
.B1(n_7282),
.B2(n_7073),
.C(n_6936),
.Y(n_19116)
);

OAI211xp5_ASAP7_75t_L g19117 ( 
.A1(n_18971),
.A2(n_5489),
.B(n_5484),
.C(n_6161),
.Y(n_19117)
);

NOR3xp33_ASAP7_75t_L g19118 ( 
.A(n_18833),
.B(n_5403),
.C(n_5323),
.Y(n_19118)
);

AND2x2_ASAP7_75t_L g19119 ( 
.A(n_18869),
.B(n_6658),
.Y(n_19119)
);

OAI22xp5_ASAP7_75t_L g19120 ( 
.A1(n_18971),
.A2(n_6833),
.B1(n_6844),
.B2(n_6806),
.Y(n_19120)
);

NAND3xp33_ASAP7_75t_L g19121 ( 
.A(n_18971),
.B(n_5489),
.C(n_5484),
.Y(n_19121)
);

NOR2x1_ASAP7_75t_L g19122 ( 
.A(n_19017),
.B(n_6161),
.Y(n_19122)
);

NOR3xp33_ASAP7_75t_L g19123 ( 
.A(n_19020),
.B(n_5403),
.C(n_5323),
.Y(n_19123)
);

NOR3xp33_ASAP7_75t_L g19124 ( 
.A(n_19022),
.B(n_5403),
.C(n_5323),
.Y(n_19124)
);

NOR2x1_ASAP7_75t_L g19125 ( 
.A(n_18994),
.B(n_6161),
.Y(n_19125)
);

NOR2x1_ASAP7_75t_L g19126 ( 
.A(n_19089),
.B(n_6161),
.Y(n_19126)
);

NOR3xp33_ASAP7_75t_L g19127 ( 
.A(n_19002),
.B(n_5403),
.C(n_5323),
.Y(n_19127)
);

NAND4xp25_ASAP7_75t_L g19128 ( 
.A(n_19003),
.B(n_7521),
.C(n_7526),
.D(n_7508),
.Y(n_19128)
);

INVx2_ASAP7_75t_L g19129 ( 
.A(n_19015),
.Y(n_19129)
);

NAND3xp33_ASAP7_75t_L g19130 ( 
.A(n_19007),
.B(n_5489),
.C(n_6806),
.Y(n_19130)
);

NOR3xp33_ASAP7_75t_L g19131 ( 
.A(n_19112),
.B(n_5403),
.C(n_5323),
.Y(n_19131)
);

INVx1_ASAP7_75t_L g19132 ( 
.A(n_19097),
.Y(n_19132)
);

NOR2x1_ASAP7_75t_L g19133 ( 
.A(n_19070),
.B(n_6161),
.Y(n_19133)
);

AND2x2_ASAP7_75t_L g19134 ( 
.A(n_19025),
.B(n_19026),
.Y(n_19134)
);

AND2x2_ASAP7_75t_L g19135 ( 
.A(n_18991),
.B(n_6658),
.Y(n_19135)
);

NOR2x1_ASAP7_75t_L g19136 ( 
.A(n_18998),
.B(n_6167),
.Y(n_19136)
);

NOR2x1_ASAP7_75t_L g19137 ( 
.A(n_18992),
.B(n_6167),
.Y(n_19137)
);

AO22x2_ASAP7_75t_L g19138 ( 
.A1(n_19046),
.A2(n_7106),
.B1(n_7110),
.B2(n_7057),
.Y(n_19138)
);

NAND3xp33_ASAP7_75t_L g19139 ( 
.A(n_19032),
.B(n_5489),
.C(n_6833),
.Y(n_19139)
);

NAND3xp33_ASAP7_75t_SL g19140 ( 
.A(n_19064),
.B(n_5564),
.C(n_5553),
.Y(n_19140)
);

NAND3xp33_ASAP7_75t_SL g19141 ( 
.A(n_19072),
.B(n_5564),
.C(n_5553),
.Y(n_19141)
);

NOR3xp33_ASAP7_75t_SL g19142 ( 
.A(n_19019),
.B(n_7134),
.C(n_7128),
.Y(n_19142)
);

AOI22xp5_ASAP7_75t_L g19143 ( 
.A1(n_18989),
.A2(n_6844),
.B1(n_6936),
.B2(n_6833),
.Y(n_19143)
);

NOR3xp33_ASAP7_75t_L g19144 ( 
.A(n_19092),
.B(n_5429),
.C(n_5411),
.Y(n_19144)
);

NAND4xp75_ASAP7_75t_L g19145 ( 
.A(n_19057),
.B(n_7390),
.C(n_7501),
.D(n_7336),
.Y(n_19145)
);

NAND4xp25_ASAP7_75t_L g19146 ( 
.A(n_19068),
.B(n_7532),
.C(n_7543),
.D(n_7526),
.Y(n_19146)
);

NAND2xp5_ASAP7_75t_L g19147 ( 
.A(n_19093),
.B(n_6658),
.Y(n_19147)
);

NAND2xp5_ASAP7_75t_L g19148 ( 
.A(n_19118),
.B(n_6693),
.Y(n_19148)
);

NAND4xp75_ASAP7_75t_L g19149 ( 
.A(n_19029),
.B(n_7390),
.C(n_7501),
.D(n_7336),
.Y(n_19149)
);

INVx1_ASAP7_75t_L g19150 ( 
.A(n_19012),
.Y(n_19150)
);

NAND2xp5_ASAP7_75t_L g19151 ( 
.A(n_19067),
.B(n_6693),
.Y(n_19151)
);

NAND2xp5_ASAP7_75t_L g19152 ( 
.A(n_19031),
.B(n_6693),
.Y(n_19152)
);

NAND3xp33_ASAP7_75t_L g19153 ( 
.A(n_19049),
.B(n_5489),
.C(n_6833),
.Y(n_19153)
);

NOR2xp33_ASAP7_75t_L g19154 ( 
.A(n_19055),
.B(n_19037),
.Y(n_19154)
);

NOR2xp33_ASAP7_75t_L g19155 ( 
.A(n_19048),
.B(n_5489),
.Y(n_19155)
);

NAND3xp33_ASAP7_75t_L g19156 ( 
.A(n_19079),
.B(n_6844),
.C(n_6833),
.Y(n_19156)
);

INVx1_ASAP7_75t_L g19157 ( 
.A(n_19041),
.Y(n_19157)
);

NAND4xp75_ASAP7_75t_L g19158 ( 
.A(n_19104),
.B(n_7390),
.C(n_7501),
.D(n_7336),
.Y(n_19158)
);

INVx1_ASAP7_75t_L g19159 ( 
.A(n_18988),
.Y(n_19159)
);

AOI22xp5_ASAP7_75t_L g19160 ( 
.A1(n_18986),
.A2(n_6844),
.B1(n_6936),
.B2(n_6833),
.Y(n_19160)
);

INVx1_ASAP7_75t_L g19161 ( 
.A(n_19113),
.Y(n_19161)
);

NOR3xp33_ASAP7_75t_L g19162 ( 
.A(n_19077),
.B(n_5429),
.C(n_5411),
.Y(n_19162)
);

NAND4xp75_ASAP7_75t_L g19163 ( 
.A(n_19043),
.B(n_7630),
.C(n_7390),
.D(n_7715),
.Y(n_19163)
);

NOR3xp33_ASAP7_75t_L g19164 ( 
.A(n_19086),
.B(n_5429),
.C(n_5411),
.Y(n_19164)
);

NAND4xp75_ASAP7_75t_L g19165 ( 
.A(n_19024),
.B(n_7630),
.C(n_7715),
.D(n_5873),
.Y(n_19165)
);

NAND3xp33_ASAP7_75t_L g19166 ( 
.A(n_19100),
.B(n_6844),
.C(n_6833),
.Y(n_19166)
);

NOR2xp33_ASAP7_75t_SL g19167 ( 
.A(n_19078),
.B(n_6157),
.Y(n_19167)
);

NAND4xp75_ASAP7_75t_L g19168 ( 
.A(n_19039),
.B(n_7630),
.C(n_7715),
.D(n_5873),
.Y(n_19168)
);

NAND4xp25_ASAP7_75t_L g19169 ( 
.A(n_19121),
.B(n_7543),
.C(n_7549),
.D(n_7532),
.Y(n_19169)
);

NOR3xp33_ASAP7_75t_L g19170 ( 
.A(n_19105),
.B(n_5429),
.C(n_5411),
.Y(n_19170)
);

NAND2xp5_ASAP7_75t_L g19171 ( 
.A(n_19063),
.B(n_6693),
.Y(n_19171)
);

NAND3xp33_ASAP7_75t_SL g19172 ( 
.A(n_19016),
.B(n_5564),
.C(n_5553),
.Y(n_19172)
);

NAND4xp75_ASAP7_75t_L g19173 ( 
.A(n_19090),
.B(n_7630),
.C(n_7715),
.D(n_5873),
.Y(n_19173)
);

INVx1_ASAP7_75t_L g19174 ( 
.A(n_19056),
.Y(n_19174)
);

NOR3xp33_ASAP7_75t_L g19175 ( 
.A(n_18990),
.B(n_5429),
.C(n_5411),
.Y(n_19175)
);

INVx1_ASAP7_75t_L g19176 ( 
.A(n_19051),
.Y(n_19176)
);

NOR2x1_ASAP7_75t_L g19177 ( 
.A(n_19011),
.B(n_6167),
.Y(n_19177)
);

NOR2x1_ASAP7_75t_L g19178 ( 
.A(n_19033),
.B(n_6167),
.Y(n_19178)
);

NOR2x1_ASAP7_75t_L g19179 ( 
.A(n_19117),
.B(n_6167),
.Y(n_19179)
);

HB1xp67_ASAP7_75t_L g19180 ( 
.A(n_19058),
.Y(n_19180)
);

NAND2xp5_ASAP7_75t_L g19181 ( 
.A(n_19023),
.B(n_6693),
.Y(n_19181)
);

INVxp67_ASAP7_75t_L g19182 ( 
.A(n_19071),
.Y(n_19182)
);

AND2x2_ASAP7_75t_L g19183 ( 
.A(n_19091),
.B(n_6693),
.Y(n_19183)
);

NOR4xp25_ASAP7_75t_L g19184 ( 
.A(n_19004),
.B(n_7106),
.C(n_7110),
.D(n_7057),
.Y(n_19184)
);

NAND3xp33_ASAP7_75t_SL g19185 ( 
.A(n_18983),
.B(n_5681),
.C(n_5564),
.Y(n_19185)
);

INVx1_ASAP7_75t_L g19186 ( 
.A(n_19027),
.Y(n_19186)
);

OR2x2_ASAP7_75t_L g19187 ( 
.A(n_19119),
.B(n_8790),
.Y(n_19187)
);

INVx1_ASAP7_75t_L g19188 ( 
.A(n_19108),
.Y(n_19188)
);

INVx1_ASAP7_75t_L g19189 ( 
.A(n_19087),
.Y(n_19189)
);

NAND3xp33_ASAP7_75t_L g19190 ( 
.A(n_19042),
.B(n_6936),
.C(n_6844),
.Y(n_19190)
);

NOR4xp25_ASAP7_75t_L g19191 ( 
.A(n_19081),
.B(n_7132),
.C(n_7158),
.D(n_7106),
.Y(n_19191)
);

NOR2x1_ASAP7_75t_L g19192 ( 
.A(n_19021),
.B(n_6248),
.Y(n_19192)
);

NOR3xp33_ASAP7_75t_L g19193 ( 
.A(n_18981),
.B(n_5443),
.C(n_5429),
.Y(n_19193)
);

NOR2x1_ASAP7_75t_L g19194 ( 
.A(n_19095),
.B(n_19060),
.Y(n_19194)
);

AOI211x1_ASAP7_75t_L g19195 ( 
.A1(n_18999),
.A2(n_7286),
.B(n_7145),
.C(n_7160),
.Y(n_19195)
);

INVx1_ASAP7_75t_L g19196 ( 
.A(n_19062),
.Y(n_19196)
);

NOR3xp33_ASAP7_75t_L g19197 ( 
.A(n_18982),
.B(n_5462),
.C(n_5443),
.Y(n_19197)
);

NOR4xp25_ASAP7_75t_L g19198 ( 
.A(n_19101),
.B(n_19109),
.C(n_19083),
.D(n_19001),
.Y(n_19198)
);

OAI222xp33_ASAP7_75t_L g19199 ( 
.A1(n_18997),
.A2(n_7290),
.B1(n_7225),
.B2(n_7303),
.C1(n_7262),
.C2(n_7254),
.Y(n_19199)
);

NAND3x1_ASAP7_75t_SL g19200 ( 
.A(n_18996),
.B(n_7605),
.C(n_7398),
.Y(n_19200)
);

NAND3xp33_ASAP7_75t_SL g19201 ( 
.A(n_19030),
.B(n_5687),
.C(n_5681),
.Y(n_19201)
);

NAND2x1p5_ASAP7_75t_L g19202 ( 
.A(n_19085),
.B(n_5443),
.Y(n_19202)
);

INVx1_ASAP7_75t_L g19203 ( 
.A(n_18984),
.Y(n_19203)
);

NOR4xp25_ASAP7_75t_L g19204 ( 
.A(n_19076),
.B(n_19047),
.C(n_18993),
.D(n_19005),
.Y(n_19204)
);

INVxp67_ASAP7_75t_SL g19205 ( 
.A(n_19050),
.Y(n_19205)
);

OA21x2_ASAP7_75t_L g19206 ( 
.A1(n_19099),
.A2(n_19103),
.B(n_19000),
.Y(n_19206)
);

NAND3xp33_ASAP7_75t_L g19207 ( 
.A(n_19034),
.B(n_6936),
.C(n_6844),
.Y(n_19207)
);

INVx1_ASAP7_75t_SL g19208 ( 
.A(n_19120),
.Y(n_19208)
);

INVx1_ASAP7_75t_L g19209 ( 
.A(n_19036),
.Y(n_19209)
);

NAND3xp33_ASAP7_75t_L g19210 ( 
.A(n_18995),
.B(n_6941),
.C(n_6936),
.Y(n_19210)
);

NAND2xp5_ASAP7_75t_L g19211 ( 
.A(n_19061),
.B(n_6701),
.Y(n_19211)
);

INVx1_ASAP7_75t_L g19212 ( 
.A(n_19059),
.Y(n_19212)
);

INVx1_ASAP7_75t_L g19213 ( 
.A(n_19013),
.Y(n_19213)
);

AND2x4_ASAP7_75t_L g19214 ( 
.A(n_19096),
.B(n_8279),
.Y(n_19214)
);

NOR2x1_ASAP7_75t_L g19215 ( 
.A(n_19094),
.B(n_6248),
.Y(n_19215)
);

INVx1_ASAP7_75t_L g19216 ( 
.A(n_19082),
.Y(n_19216)
);

INVx2_ASAP7_75t_L g19217 ( 
.A(n_19028),
.Y(n_19217)
);

NOR2xp67_ASAP7_75t_L g19218 ( 
.A(n_19115),
.B(n_5443),
.Y(n_19218)
);

NOR2x1_ASAP7_75t_L g19219 ( 
.A(n_19006),
.B(n_6248),
.Y(n_19219)
);

INVx1_ASAP7_75t_L g19220 ( 
.A(n_19088),
.Y(n_19220)
);

NAND4xp75_ASAP7_75t_L g19221 ( 
.A(n_19098),
.B(n_7715),
.C(n_5866),
.D(n_4871),
.Y(n_19221)
);

NAND2xp5_ASAP7_75t_L g19222 ( 
.A(n_19065),
.B(n_6701),
.Y(n_19222)
);

NAND4xp75_ASAP7_75t_L g19223 ( 
.A(n_19106),
.B(n_5866),
.C(n_4927),
.D(n_4932),
.Y(n_19223)
);

NOR2x1_ASAP7_75t_L g19224 ( 
.A(n_19008),
.B(n_6248),
.Y(n_19224)
);

NOR3xp33_ASAP7_75t_L g19225 ( 
.A(n_19084),
.B(n_5462),
.C(n_5443),
.Y(n_19225)
);

HB1xp67_ASAP7_75t_L g19226 ( 
.A(n_19066),
.Y(n_19226)
);

NAND3xp33_ASAP7_75t_SL g19227 ( 
.A(n_19018),
.B(n_5687),
.C(n_5681),
.Y(n_19227)
);

NOR3xp33_ASAP7_75t_L g19228 ( 
.A(n_19069),
.B(n_5462),
.C(n_5443),
.Y(n_19228)
);

NAND4xp25_ASAP7_75t_L g19229 ( 
.A(n_19107),
.B(n_7543),
.C(n_7549),
.D(n_7532),
.Y(n_19229)
);

NAND4xp25_ASAP7_75t_L g19230 ( 
.A(n_19110),
.B(n_7549),
.C(n_7575),
.D(n_7543),
.Y(n_19230)
);

INVx1_ASAP7_75t_L g19231 ( 
.A(n_18987),
.Y(n_19231)
);

AOI21xp5_ASAP7_75t_L g19232 ( 
.A1(n_18985),
.A2(n_19045),
.B(n_19010),
.Y(n_19232)
);

NAND3xp33_ASAP7_75t_SL g19233 ( 
.A(n_19053),
.B(n_5687),
.C(n_5681),
.Y(n_19233)
);

AO22x2_ASAP7_75t_L g19234 ( 
.A1(n_19073),
.A2(n_7158),
.B1(n_7218),
.B2(n_7132),
.Y(n_19234)
);

INVx1_ASAP7_75t_L g19235 ( 
.A(n_19116),
.Y(n_19235)
);

NOR2xp67_ASAP7_75t_SL g19236 ( 
.A(n_19074),
.B(n_19114),
.Y(n_19236)
);

NAND2xp5_ASAP7_75t_L g19237 ( 
.A(n_19111),
.B(n_6701),
.Y(n_19237)
);

AND3x4_ASAP7_75t_L g19238 ( 
.A(n_19035),
.B(n_6350),
.C(n_5890),
.Y(n_19238)
);

NAND4xp25_ASAP7_75t_L g19239 ( 
.A(n_19075),
.B(n_7575),
.C(n_7549),
.D(n_5881),
.Y(n_19239)
);

NAND3xp33_ASAP7_75t_L g19240 ( 
.A(n_19054),
.B(n_6941),
.C(n_6936),
.Y(n_19240)
);

NAND2xp5_ASAP7_75t_SL g19241 ( 
.A(n_19134),
.B(n_19040),
.Y(n_19241)
);

NAND2xp5_ASAP7_75t_SL g19242 ( 
.A(n_19129),
.B(n_19009),
.Y(n_19242)
);

NOR2x1_ASAP7_75t_L g19243 ( 
.A(n_19157),
.B(n_19080),
.Y(n_19243)
);

AOI322xp5_ASAP7_75t_L g19244 ( 
.A1(n_19155),
.A2(n_19038),
.A3(n_19014),
.B1(n_19052),
.B2(n_19102),
.C1(n_19044),
.C2(n_7280),
.Y(n_19244)
);

OAI211xp5_ASAP7_75t_L g19245 ( 
.A1(n_19154),
.A2(n_6342),
.B(n_6373),
.C(n_6248),
.Y(n_19245)
);

NAND4xp25_ASAP7_75t_L g19246 ( 
.A(n_19231),
.B(n_4475),
.C(n_4497),
.D(n_4474),
.Y(n_19246)
);

OAI21xp33_ASAP7_75t_L g19247 ( 
.A1(n_19167),
.A2(n_7158),
.B(n_7132),
.Y(n_19247)
);

OAI211xp5_ASAP7_75t_SL g19248 ( 
.A1(n_19182),
.A2(n_5462),
.B(n_5481),
.C(n_5472),
.Y(n_19248)
);

AOI22xp33_ASAP7_75t_L g19249 ( 
.A1(n_19123),
.A2(n_6948),
.B1(n_6951),
.B2(n_6941),
.Y(n_19249)
);

INVx1_ASAP7_75t_L g19250 ( 
.A(n_19186),
.Y(n_19250)
);

OAI211xp5_ASAP7_75t_SL g19251 ( 
.A1(n_19176),
.A2(n_5462),
.B(n_5481),
.C(n_5472),
.Y(n_19251)
);

NAND3xp33_ASAP7_75t_L g19252 ( 
.A(n_19174),
.B(n_6948),
.C(n_6941),
.Y(n_19252)
);

NOR4xp75_ASAP7_75t_SL g19253 ( 
.A(n_19171),
.B(n_7145),
.C(n_7160),
.D(n_7157),
.Y(n_19253)
);

OAI211xp5_ASAP7_75t_L g19254 ( 
.A1(n_19226),
.A2(n_6373),
.B(n_6381),
.C(n_6342),
.Y(n_19254)
);

AOI22xp5_ASAP7_75t_L g19255 ( 
.A1(n_19156),
.A2(n_6948),
.B1(n_6951),
.B2(n_6941),
.Y(n_19255)
);

AOI221x1_ASAP7_75t_SL g19256 ( 
.A1(n_19203),
.A2(n_6911),
.B1(n_7037),
.B2(n_6969),
.C(n_6916),
.Y(n_19256)
);

AND4x1_ASAP7_75t_L g19257 ( 
.A(n_19132),
.B(n_7157),
.C(n_7174),
.D(n_7160),
.Y(n_19257)
);

NOR2x1_ASAP7_75t_L g19258 ( 
.A(n_19159),
.B(n_6342),
.Y(n_19258)
);

AOI21xp5_ASAP7_75t_L g19259 ( 
.A1(n_19232),
.A2(n_7564),
.B(n_8279),
.Y(n_19259)
);

OAI22xp5_ASAP7_75t_L g19260 ( 
.A1(n_19130),
.A2(n_6948),
.B1(n_6951),
.B2(n_6941),
.Y(n_19260)
);

NAND4xp25_ASAP7_75t_L g19261 ( 
.A(n_19220),
.B(n_4475),
.C(n_4497),
.D(n_4474),
.Y(n_19261)
);

AOI221xp5_ASAP7_75t_L g19262 ( 
.A1(n_19204),
.A2(n_7431),
.B1(n_7437),
.B2(n_7073),
.C(n_7019),
.Y(n_19262)
);

NOR3xp33_ASAP7_75t_L g19263 ( 
.A(n_19161),
.B(n_5472),
.C(n_5462),
.Y(n_19263)
);

OAI21xp5_ASAP7_75t_L g19264 ( 
.A1(n_19126),
.A2(n_8597),
.B(n_8591),
.Y(n_19264)
);

NAND4xp25_ASAP7_75t_SL g19265 ( 
.A(n_19127),
.B(n_6885),
.C(n_6902),
.D(n_6887),
.Y(n_19265)
);

NAND3xp33_ASAP7_75t_L g19266 ( 
.A(n_19180),
.B(n_6948),
.C(n_6941),
.Y(n_19266)
);

NAND5xp2_ASAP7_75t_L g19267 ( 
.A(n_19196),
.B(n_5866),
.C(n_5864),
.D(n_5853),
.E(n_7398),
.Y(n_19267)
);

NOR3xp33_ASAP7_75t_L g19268 ( 
.A(n_19208),
.B(n_5481),
.C(n_5472),
.Y(n_19268)
);

OAI221xp5_ASAP7_75t_L g19269 ( 
.A1(n_19133),
.A2(n_5386),
.B1(n_5348),
.B2(n_4962),
.C(n_7575),
.Y(n_19269)
);

NOR2xp33_ASAP7_75t_L g19270 ( 
.A(n_19209),
.B(n_19217),
.Y(n_19270)
);

OR5x1_ASAP7_75t_L g19271 ( 
.A(n_19233),
.B(n_19128),
.C(n_19185),
.D(n_19141),
.E(n_19201),
.Y(n_19271)
);

NOR4xp25_ASAP7_75t_L g19272 ( 
.A(n_19212),
.B(n_7218),
.C(n_7224),
.D(n_7158),
.Y(n_19272)
);

NOR2xp33_ASAP7_75t_L g19273 ( 
.A(n_19216),
.B(n_4962),
.Y(n_19273)
);

NAND2xp5_ASAP7_75t_L g19274 ( 
.A(n_19150),
.B(n_6701),
.Y(n_19274)
);

OAI211xp5_ASAP7_75t_L g19275 ( 
.A1(n_19205),
.A2(n_6373),
.B(n_6381),
.C(n_6342),
.Y(n_19275)
);

NOR3xp33_ASAP7_75t_SL g19276 ( 
.A(n_19235),
.B(n_7174),
.C(n_7157),
.Y(n_19276)
);

AOI221xp5_ASAP7_75t_SL g19277 ( 
.A1(n_19188),
.A2(n_6951),
.B1(n_6989),
.B2(n_6948),
.C(n_6941),
.Y(n_19277)
);

NAND2xp5_ASAP7_75t_L g19278 ( 
.A(n_19122),
.B(n_6701),
.Y(n_19278)
);

AOI211xp5_ASAP7_75t_SL g19279 ( 
.A1(n_19213),
.A2(n_5481),
.B(n_5501),
.C(n_5472),
.Y(n_19279)
);

INVx1_ASAP7_75t_L g19280 ( 
.A(n_19206),
.Y(n_19280)
);

NAND4xp25_ASAP7_75t_SL g19281 ( 
.A(n_19124),
.B(n_6887),
.C(n_6902),
.D(n_6885),
.Y(n_19281)
);

NOR2xp33_ASAP7_75t_L g19282 ( 
.A(n_19189),
.B(n_4962),
.Y(n_19282)
);

NAND3xp33_ASAP7_75t_L g19283 ( 
.A(n_19236),
.B(n_6951),
.C(n_6948),
.Y(n_19283)
);

OAI211xp5_ASAP7_75t_SL g19284 ( 
.A1(n_19219),
.A2(n_5472),
.B(n_5501),
.C(n_5481),
.Y(n_19284)
);

O2A1O1Ixp5_ASAP7_75t_L g19285 ( 
.A1(n_19139),
.A2(n_7218),
.B(n_7224),
.C(n_7158),
.Y(n_19285)
);

AND2x4_ASAP7_75t_L g19286 ( 
.A(n_19218),
.B(n_6657),
.Y(n_19286)
);

AOI211x1_ASAP7_75t_SL g19287 ( 
.A1(n_19172),
.A2(n_7136),
.B(n_7304),
.C(n_7009),
.Y(n_19287)
);

OAI21xp5_ASAP7_75t_L g19288 ( 
.A1(n_19153),
.A2(n_8597),
.B(n_8591),
.Y(n_19288)
);

NAND4xp25_ASAP7_75t_L g19289 ( 
.A(n_19162),
.B(n_4475),
.C(n_4497),
.D(n_4474),
.Y(n_19289)
);

AOI211xp5_ASAP7_75t_L g19290 ( 
.A1(n_19198),
.A2(n_19131),
.B(n_19164),
.C(n_19227),
.Y(n_19290)
);

AO22x2_ASAP7_75t_L g19291 ( 
.A1(n_19238),
.A2(n_7224),
.B1(n_7280),
.B2(n_7218),
.Y(n_19291)
);

NAND4xp75_ASAP7_75t_L g19292 ( 
.A(n_19177),
.B(n_4710),
.C(n_6676),
.D(n_6634),
.Y(n_19292)
);

OAI321xp33_ASAP7_75t_L g19293 ( 
.A1(n_19211),
.A2(n_6951),
.A3(n_6989),
.B1(n_7019),
.B2(n_7009),
.C(n_6948),
.Y(n_19293)
);

AOI21xp5_ASAP7_75t_L g19294 ( 
.A1(n_19206),
.A2(n_7564),
.B(n_8279),
.Y(n_19294)
);

AND2x2_ASAP7_75t_L g19295 ( 
.A(n_19135),
.B(n_6701),
.Y(n_19295)
);

NAND5xp2_ASAP7_75t_L g19296 ( 
.A(n_19202),
.B(n_5864),
.C(n_5853),
.D(n_7605),
.E(n_7398),
.Y(n_19296)
);

OAI211xp5_ASAP7_75t_SL g19297 ( 
.A1(n_19194),
.A2(n_5481),
.B(n_5501),
.C(n_7610),
.Y(n_19297)
);

NAND3xp33_ASAP7_75t_SL g19298 ( 
.A(n_19197),
.B(n_5687),
.C(n_5681),
.Y(n_19298)
);

NAND2xp5_ASAP7_75t_SL g19299 ( 
.A(n_19125),
.B(n_6948),
.Y(n_19299)
);

XOR2xp5_ASAP7_75t_L g19300 ( 
.A(n_19215),
.B(n_6657),
.Y(n_19300)
);

NAND4xp25_ASAP7_75t_L g19301 ( 
.A(n_19136),
.B(n_4497),
.C(n_4518),
.D(n_4475),
.Y(n_19301)
);

INVx2_ASAP7_75t_SL g19302 ( 
.A(n_19137),
.Y(n_19302)
);

OAI21xp5_ASAP7_75t_L g19303 ( 
.A1(n_19207),
.A2(n_8301),
.B(n_8286),
.Y(n_19303)
);

NOR4xp25_ASAP7_75t_L g19304 ( 
.A(n_19140),
.B(n_7224),
.C(n_7280),
.D(n_7218),
.Y(n_19304)
);

NAND3xp33_ASAP7_75t_L g19305 ( 
.A(n_19144),
.B(n_6989),
.C(n_6951),
.Y(n_19305)
);

NAND4xp25_ASAP7_75t_L g19306 ( 
.A(n_19224),
.B(n_19228),
.C(n_19170),
.D(n_19179),
.Y(n_19306)
);

NAND4xp75_ASAP7_75t_L g19307 ( 
.A(n_19192),
.B(n_6676),
.C(n_6634),
.D(n_7174),
.Y(n_19307)
);

OAI221xp5_ASAP7_75t_L g19308 ( 
.A1(n_19222),
.A2(n_5386),
.B1(n_5348),
.B2(n_4962),
.C(n_7575),
.Y(n_19308)
);

NOR2xp33_ASAP7_75t_L g19309 ( 
.A(n_19152),
.B(n_4962),
.Y(n_19309)
);

NAND2xp5_ASAP7_75t_SL g19310 ( 
.A(n_19237),
.B(n_6989),
.Y(n_19310)
);

NAND4xp25_ASAP7_75t_L g19311 ( 
.A(n_19151),
.B(n_4497),
.C(n_4518),
.D(n_4475),
.Y(n_19311)
);

NAND2xp5_ASAP7_75t_L g19312 ( 
.A(n_19225),
.B(n_7997),
.Y(n_19312)
);

NOR3xp33_ASAP7_75t_L g19313 ( 
.A(n_19200),
.B(n_5501),
.C(n_4497),
.Y(n_19313)
);

AOI21xp5_ASAP7_75t_L g19314 ( 
.A1(n_19147),
.A2(n_7564),
.B(n_8286),
.Y(n_19314)
);

AOI221xp5_ASAP7_75t_L g19315 ( 
.A1(n_19184),
.A2(n_6989),
.B1(n_7437),
.B2(n_7431),
.C(n_7073),
.Y(n_19315)
);

AOI211xp5_ASAP7_75t_L g19316 ( 
.A1(n_19193),
.A2(n_8286),
.B(n_8301),
.C(n_8176),
.Y(n_19316)
);

NOR3xp33_ASAP7_75t_L g19317 ( 
.A(n_19148),
.B(n_5501),
.C(n_4518),
.Y(n_19317)
);

NOR2xp33_ASAP7_75t_L g19318 ( 
.A(n_19173),
.B(n_4962),
.Y(n_19318)
);

NAND2xp5_ASAP7_75t_L g19319 ( 
.A(n_19178),
.B(n_7997),
.Y(n_19319)
);

AOI211xp5_ASAP7_75t_L g19320 ( 
.A1(n_19190),
.A2(n_8301),
.B(n_8176),
.C(n_8137),
.Y(n_19320)
);

AND2x4_ASAP7_75t_L g19321 ( 
.A(n_19183),
.B(n_6682),
.Y(n_19321)
);

OAI211xp5_ASAP7_75t_SL g19322 ( 
.A1(n_19181),
.A2(n_5501),
.B(n_7610),
.C(n_7312),
.Y(n_19322)
);

AOI221xp5_ASAP7_75t_L g19323 ( 
.A1(n_19191),
.A2(n_7175),
.B1(n_7282),
.B2(n_7141),
.C(n_7094),
.Y(n_19323)
);

AOI211xp5_ASAP7_75t_L g19324 ( 
.A1(n_19240),
.A2(n_8140),
.B(n_8142),
.C(n_8137),
.Y(n_19324)
);

NAND4xp25_ASAP7_75t_L g19325 ( 
.A(n_19195),
.B(n_4518),
.C(n_4475),
.D(n_5876),
.Y(n_19325)
);

AOI22xp5_ASAP7_75t_SL g19326 ( 
.A1(n_19214),
.A2(n_4748),
.B1(n_4608),
.B2(n_4544),
.Y(n_19326)
);

OAI211xp5_ASAP7_75t_L g19327 ( 
.A1(n_19239),
.A2(n_6373),
.B(n_6381),
.C(n_6342),
.Y(n_19327)
);

AND2x2_ASAP7_75t_L g19328 ( 
.A(n_19142),
.B(n_8137),
.Y(n_19328)
);

NAND4xp25_ASAP7_75t_L g19329 ( 
.A(n_19175),
.B(n_4518),
.C(n_5881),
.D(n_5876),
.Y(n_19329)
);

NAND4xp75_ASAP7_75t_L g19330 ( 
.A(n_19143),
.B(n_6676),
.C(n_6634),
.D(n_7176),
.Y(n_19330)
);

OAI211xp5_ASAP7_75t_L g19331 ( 
.A1(n_19166),
.A2(n_6381),
.B(n_6393),
.C(n_6373),
.Y(n_19331)
);

AOI221xp5_ASAP7_75t_L g19332 ( 
.A1(n_19234),
.A2(n_7461),
.B1(n_7481),
.B2(n_7221),
.C(n_7147),
.Y(n_19332)
);

NAND5xp2_ASAP7_75t_L g19333 ( 
.A(n_19160),
.B(n_5864),
.C(n_5853),
.D(n_7605),
.E(n_7398),
.Y(n_19333)
);

NAND5xp2_ASAP7_75t_L g19334 ( 
.A(n_19158),
.B(n_7605),
.C(n_7398),
.D(n_6575),
.E(n_6676),
.Y(n_19334)
);

NAND3xp33_ASAP7_75t_SL g19335 ( 
.A(n_19187),
.B(n_5694),
.C(n_5687),
.Y(n_19335)
);

NAND3xp33_ASAP7_75t_L g19336 ( 
.A(n_19210),
.B(n_19230),
.C(n_19229),
.Y(n_19336)
);

AOI221xp5_ASAP7_75t_L g19337 ( 
.A1(n_19234),
.A2(n_6989),
.B1(n_7437),
.B2(n_7431),
.C(n_7073),
.Y(n_19337)
);

NOR2xp33_ASAP7_75t_L g19338 ( 
.A(n_19223),
.B(n_19149),
.Y(n_19338)
);

NAND3xp33_ASAP7_75t_L g19339 ( 
.A(n_19169),
.B(n_7009),
.C(n_6989),
.Y(n_19339)
);

OAI211xp5_ASAP7_75t_L g19340 ( 
.A1(n_19146),
.A2(n_6393),
.B(n_6461),
.C(n_6381),
.Y(n_19340)
);

NAND2xp5_ASAP7_75t_L g19341 ( 
.A(n_19145),
.B(n_19168),
.Y(n_19341)
);

INVx1_ASAP7_75t_L g19342 ( 
.A(n_19138),
.Y(n_19342)
);

NOR2x1_ASAP7_75t_L g19343 ( 
.A(n_19221),
.B(n_19165),
.Y(n_19343)
);

NAND4xp75_ASAP7_75t_L g19344 ( 
.A(n_19243),
.B(n_19138),
.C(n_19199),
.D(n_19163),
.Y(n_19344)
);

OR2x2_ASAP7_75t_L g19345 ( 
.A(n_19278),
.B(n_19214),
.Y(n_19345)
);

INVx1_ASAP7_75t_L g19346 ( 
.A(n_19280),
.Y(n_19346)
);

INVxp67_ASAP7_75t_L g19347 ( 
.A(n_19270),
.Y(n_19347)
);

INVx2_ASAP7_75t_L g19348 ( 
.A(n_19250),
.Y(n_19348)
);

NOR2xp33_ASAP7_75t_SL g19349 ( 
.A(n_19302),
.B(n_7398),
.Y(n_19349)
);

INVx1_ASAP7_75t_L g19350 ( 
.A(n_19341),
.Y(n_19350)
);

INVx1_ASAP7_75t_L g19351 ( 
.A(n_19282),
.Y(n_19351)
);

XOR2xp5_ASAP7_75t_L g19352 ( 
.A(n_19242),
.B(n_4819),
.Y(n_19352)
);

INVxp33_ASAP7_75t_L g19353 ( 
.A(n_19241),
.Y(n_19353)
);

AND2x4_ASAP7_75t_L g19354 ( 
.A(n_19321),
.B(n_19295),
.Y(n_19354)
);

NOR3xp33_ASAP7_75t_L g19355 ( 
.A(n_19290),
.B(n_4518),
.C(n_5694),
.Y(n_19355)
);

NAND4xp75_ASAP7_75t_L g19356 ( 
.A(n_19343),
.B(n_6634),
.C(n_7011),
.D(n_6998),
.Y(n_19356)
);

NAND2x1p5_ASAP7_75t_SL g19357 ( 
.A(n_19258),
.B(n_5783),
.Y(n_19357)
);

NAND2xp5_ASAP7_75t_L g19358 ( 
.A(n_19286),
.B(n_7997),
.Y(n_19358)
);

NAND2xp5_ASAP7_75t_L g19359 ( 
.A(n_19286),
.B(n_19300),
.Y(n_19359)
);

NAND2xp33_ASAP7_75t_L g19360 ( 
.A(n_19336),
.B(n_19342),
.Y(n_19360)
);

NOR4xp75_ASAP7_75t_L g19361 ( 
.A(n_19310),
.B(n_19247),
.C(n_19292),
.D(n_19274),
.Y(n_19361)
);

AND2x4_ASAP7_75t_L g19362 ( 
.A(n_19321),
.B(n_6682),
.Y(n_19362)
);

HB1xp67_ASAP7_75t_L g19363 ( 
.A(n_19338),
.Y(n_19363)
);

INVx2_ASAP7_75t_L g19364 ( 
.A(n_19271),
.Y(n_19364)
);

NAND4xp75_ASAP7_75t_L g19365 ( 
.A(n_19273),
.B(n_7011),
.C(n_7017),
.D(n_6998),
.Y(n_19365)
);

OR2x2_ASAP7_75t_L g19366 ( 
.A(n_19296),
.B(n_8790),
.Y(n_19366)
);

INVx2_ASAP7_75t_L g19367 ( 
.A(n_19291),
.Y(n_19367)
);

INVx1_ASAP7_75t_L g19368 ( 
.A(n_19306),
.Y(n_19368)
);

AOI22xp5_ASAP7_75t_L g19369 ( 
.A1(n_19283),
.A2(n_7019),
.B1(n_7073),
.B2(n_7009),
.Y(n_19369)
);

INVx1_ASAP7_75t_L g19370 ( 
.A(n_19309),
.Y(n_19370)
);

AOI22xp5_ASAP7_75t_L g19371 ( 
.A1(n_19252),
.A2(n_19318),
.B1(n_19268),
.B2(n_19313),
.Y(n_19371)
);

NAND2x1p5_ASAP7_75t_L g19372 ( 
.A(n_19299),
.B(n_5694),
.Y(n_19372)
);

INVx1_ASAP7_75t_L g19373 ( 
.A(n_19335),
.Y(n_19373)
);

INVx1_ASAP7_75t_L g19374 ( 
.A(n_19291),
.Y(n_19374)
);

INVxp33_ASAP7_75t_L g19375 ( 
.A(n_19263),
.Y(n_19375)
);

XOR2x2_ASAP7_75t_L g19376 ( 
.A(n_19307),
.B(n_5876),
.Y(n_19376)
);

NOR2xp33_ASAP7_75t_L g19377 ( 
.A(n_19311),
.B(n_4962),
.Y(n_19377)
);

XNOR2xp5_ASAP7_75t_L g19378 ( 
.A(n_19287),
.B(n_6682),
.Y(n_19378)
);

INVx2_ASAP7_75t_L g19379 ( 
.A(n_19285),
.Y(n_19379)
);

NOR2xp33_ASAP7_75t_L g19380 ( 
.A(n_19284),
.B(n_5348),
.Y(n_19380)
);

NAND4xp75_ASAP7_75t_L g19381 ( 
.A(n_19277),
.B(n_7011),
.C(n_7017),
.D(n_6998),
.Y(n_19381)
);

INVx1_ASAP7_75t_L g19382 ( 
.A(n_19317),
.Y(n_19382)
);

NOR4xp25_ASAP7_75t_L g19383 ( 
.A(n_19298),
.B(n_7224),
.C(n_7280),
.D(n_7218),
.Y(n_19383)
);

AND2x4_ASAP7_75t_L g19384 ( 
.A(n_19276),
.B(n_6692),
.Y(n_19384)
);

INVxp33_ASAP7_75t_SL g19385 ( 
.A(n_19328),
.Y(n_19385)
);

NAND4xp75_ASAP7_75t_L g19386 ( 
.A(n_19294),
.B(n_19319),
.C(n_19314),
.D(n_19262),
.Y(n_19386)
);

NOR2xp33_ASAP7_75t_L g19387 ( 
.A(n_19261),
.B(n_5348),
.Y(n_19387)
);

INVx2_ASAP7_75t_L g19388 ( 
.A(n_19330),
.Y(n_19388)
);

XNOR2xp5_ASAP7_75t_L g19389 ( 
.A(n_19325),
.B(n_6682),
.Y(n_19389)
);

AND2x2_ASAP7_75t_L g19390 ( 
.A(n_19244),
.B(n_7605),
.Y(n_19390)
);

NOR2x1_ASAP7_75t_L g19391 ( 
.A(n_19301),
.B(n_6393),
.Y(n_19391)
);

NOR2x1_ASAP7_75t_L g19392 ( 
.A(n_19289),
.B(n_6393),
.Y(n_19392)
);

OAI22xp5_ASAP7_75t_L g19393 ( 
.A1(n_19266),
.A2(n_7019),
.B1(n_7073),
.B2(n_7009),
.Y(n_19393)
);

NOR2x1_ASAP7_75t_SL g19394 ( 
.A(n_19327),
.B(n_19340),
.Y(n_19394)
);

NAND4xp75_ASAP7_75t_L g19395 ( 
.A(n_19312),
.B(n_7011),
.C(n_7017),
.D(n_6998),
.Y(n_19395)
);

INVx2_ASAP7_75t_L g19396 ( 
.A(n_19269),
.Y(n_19396)
);

NOR2xp67_ASAP7_75t_L g19397 ( 
.A(n_19246),
.B(n_5694),
.Y(n_19397)
);

AND2x4_ASAP7_75t_L g19398 ( 
.A(n_19339),
.B(n_19305),
.Y(n_19398)
);

OAI22xp5_ASAP7_75t_L g19399 ( 
.A1(n_19308),
.A2(n_7073),
.B1(n_7094),
.B2(n_7009),
.Y(n_19399)
);

NOR2xp67_ASAP7_75t_L g19400 ( 
.A(n_19334),
.B(n_19281),
.Y(n_19400)
);

INVx1_ASAP7_75t_L g19401 ( 
.A(n_19322),
.Y(n_19401)
);

OR2x2_ASAP7_75t_L g19402 ( 
.A(n_19329),
.B(n_8790),
.Y(n_19402)
);

AOI22xp5_ASAP7_75t_L g19403 ( 
.A1(n_19265),
.A2(n_7094),
.B1(n_7111),
.B2(n_7009),
.Y(n_19403)
);

AND2x4_ASAP7_75t_L g19404 ( 
.A(n_19326),
.B(n_6692),
.Y(n_19404)
);

INVx2_ASAP7_75t_L g19405 ( 
.A(n_19253),
.Y(n_19405)
);

OAI322xp33_ASAP7_75t_L g19406 ( 
.A1(n_19259),
.A2(n_19255),
.A3(n_19260),
.B1(n_19293),
.B2(n_19304),
.C1(n_19333),
.C2(n_19251),
.Y(n_19406)
);

OAI22xp5_ASAP7_75t_L g19407 ( 
.A1(n_19245),
.A2(n_7094),
.B1(n_7111),
.B2(n_7009),
.Y(n_19407)
);

INVx1_ASAP7_75t_L g19408 ( 
.A(n_19331),
.Y(n_19408)
);

XOR2xp5_ASAP7_75t_L g19409 ( 
.A(n_19303),
.B(n_4819),
.Y(n_19409)
);

INVx1_ASAP7_75t_L g19410 ( 
.A(n_19254),
.Y(n_19410)
);

INVx2_ASAP7_75t_L g19411 ( 
.A(n_19264),
.Y(n_19411)
);

INVx2_ASAP7_75t_L g19412 ( 
.A(n_19279),
.Y(n_19412)
);

OR2x2_ASAP7_75t_L g19413 ( 
.A(n_19267),
.B(n_8790),
.Y(n_19413)
);

NAND2xp5_ASAP7_75t_L g19414 ( 
.A(n_19256),
.B(n_8183),
.Y(n_19414)
);

INVxp67_ASAP7_75t_L g19415 ( 
.A(n_19275),
.Y(n_19415)
);

NAND4xp75_ASAP7_75t_L g19416 ( 
.A(n_19323),
.B(n_7032),
.C(n_7035),
.D(n_7017),
.Y(n_19416)
);

AOI22xp5_ASAP7_75t_L g19417 ( 
.A1(n_19297),
.A2(n_7094),
.B1(n_7111),
.B2(n_7009),
.Y(n_19417)
);

AOI221xp5_ASAP7_75t_SL g19418 ( 
.A1(n_19315),
.A2(n_7136),
.B1(n_7141),
.B2(n_7111),
.C(n_7094),
.Y(n_19418)
);

INVx1_ASAP7_75t_L g19419 ( 
.A(n_19248),
.Y(n_19419)
);

NAND4xp75_ASAP7_75t_L g19420 ( 
.A(n_19288),
.B(n_7035),
.C(n_7086),
.D(n_7032),
.Y(n_19420)
);

INVx2_ASAP7_75t_L g19421 ( 
.A(n_19272),
.Y(n_19421)
);

INVx2_ASAP7_75t_L g19422 ( 
.A(n_19257),
.Y(n_19422)
);

INVx2_ASAP7_75t_SL g19423 ( 
.A(n_19324),
.Y(n_19423)
);

INVx2_ASAP7_75t_L g19424 ( 
.A(n_19316),
.Y(n_19424)
);

INVx2_ASAP7_75t_SL g19425 ( 
.A(n_19320),
.Y(n_19425)
);

INVx1_ASAP7_75t_L g19426 ( 
.A(n_19249),
.Y(n_19426)
);

NOR2x1_ASAP7_75t_L g19427 ( 
.A(n_19332),
.B(n_6393),
.Y(n_19427)
);

AND2x4_ASAP7_75t_L g19428 ( 
.A(n_19337),
.B(n_6704),
.Y(n_19428)
);

INVx1_ASAP7_75t_L g19429 ( 
.A(n_19280),
.Y(n_19429)
);

NOR4xp75_ASAP7_75t_L g19430 ( 
.A(n_19242),
.B(n_7181),
.C(n_7253),
.D(n_7176),
.Y(n_19430)
);

NOR2x1p5_ASAP7_75t_L g19431 ( 
.A(n_19250),
.B(n_5876),
.Y(n_19431)
);

INVx1_ASAP7_75t_L g19432 ( 
.A(n_19280),
.Y(n_19432)
);

INVxp67_ASAP7_75t_L g19433 ( 
.A(n_19280),
.Y(n_19433)
);

INVx1_ASAP7_75t_L g19434 ( 
.A(n_19280),
.Y(n_19434)
);

AO22x2_ASAP7_75t_L g19435 ( 
.A1(n_19280),
.A2(n_7280),
.B1(n_7287),
.B2(n_7224),
.Y(n_19435)
);

NOR3xp33_ASAP7_75t_L g19436 ( 
.A(n_19433),
.B(n_5697),
.C(n_5694),
.Y(n_19436)
);

O2A1O1Ixp33_ASAP7_75t_L g19437 ( 
.A1(n_19346),
.A2(n_5799),
.B(n_5890),
.C(n_5881),
.Y(n_19437)
);

NAND3xp33_ASAP7_75t_L g19438 ( 
.A(n_19360),
.B(n_7111),
.C(n_7094),
.Y(n_19438)
);

AND4x1_ASAP7_75t_L g19439 ( 
.A(n_19350),
.B(n_7176),
.C(n_7253),
.D(n_7181),
.Y(n_19439)
);

NAND3xp33_ASAP7_75t_SL g19440 ( 
.A(n_19353),
.B(n_5697),
.C(n_5830),
.Y(n_19440)
);

OR2x2_ASAP7_75t_SL g19441 ( 
.A(n_19348),
.B(n_5348),
.Y(n_19441)
);

NOR2x1_ASAP7_75t_L g19442 ( 
.A(n_19429),
.B(n_6461),
.Y(n_19442)
);

NAND2xp5_ASAP7_75t_L g19443 ( 
.A(n_19432),
.B(n_6853),
.Y(n_19443)
);

NOR2x1_ASAP7_75t_L g19444 ( 
.A(n_19434),
.B(n_6461),
.Y(n_19444)
);

NOR4xp25_ASAP7_75t_L g19445 ( 
.A(n_19347),
.B(n_7287),
.C(n_7294),
.D(n_7280),
.Y(n_19445)
);

NOR4xp25_ASAP7_75t_L g19446 ( 
.A(n_19364),
.B(n_7294),
.C(n_7300),
.D(n_7287),
.Y(n_19446)
);

NOR2x1p5_ASAP7_75t_L g19447 ( 
.A(n_19359),
.B(n_19388),
.Y(n_19447)
);

AND2x4_ASAP7_75t_L g19448 ( 
.A(n_19361),
.B(n_6692),
.Y(n_19448)
);

AOI22xp33_ASAP7_75t_SL g19449 ( 
.A1(n_19363),
.A2(n_5386),
.B1(n_5348),
.B2(n_6575),
.Y(n_19449)
);

AOI211xp5_ASAP7_75t_L g19450 ( 
.A1(n_19368),
.A2(n_7868),
.B(n_7869),
.C(n_7860),
.Y(n_19450)
);

NOR3xp33_ASAP7_75t_SL g19451 ( 
.A(n_19344),
.B(n_7253),
.C(n_7181),
.Y(n_19451)
);

A2O1A1Ixp33_ASAP7_75t_L g19452 ( 
.A1(n_19400),
.A2(n_8142),
.B(n_8146),
.C(n_8140),
.Y(n_19452)
);

INVx1_ASAP7_75t_L g19453 ( 
.A(n_19352),
.Y(n_19453)
);

INVxp33_ASAP7_75t_L g19454 ( 
.A(n_19354),
.Y(n_19454)
);

NOR2x2_ASAP7_75t_L g19455 ( 
.A(n_19422),
.B(n_5799),
.Y(n_19455)
);

NAND2xp5_ASAP7_75t_L g19456 ( 
.A(n_19390),
.B(n_6853),
.Y(n_19456)
);

NOR4xp25_ASAP7_75t_L g19457 ( 
.A(n_19411),
.B(n_7294),
.C(n_7300),
.D(n_7287),
.Y(n_19457)
);

INVx2_ASAP7_75t_L g19458 ( 
.A(n_19357),
.Y(n_19458)
);

NAND4xp75_ASAP7_75t_L g19459 ( 
.A(n_19351),
.B(n_7035),
.C(n_7086),
.D(n_7032),
.Y(n_19459)
);

NAND4xp25_ASAP7_75t_SL g19460 ( 
.A(n_19371),
.B(n_7269),
.C(n_7273),
.D(n_7265),
.Y(n_19460)
);

NAND2xp5_ASAP7_75t_L g19461 ( 
.A(n_19405),
.B(n_6853),
.Y(n_19461)
);

NOR5xp2_ASAP7_75t_L g19462 ( 
.A(n_19415),
.B(n_7248),
.C(n_7251),
.D(n_7237),
.E(n_7232),
.Y(n_19462)
);

NAND5xp2_ASAP7_75t_L g19463 ( 
.A(n_19385),
.B(n_7605),
.C(n_6575),
.D(n_5386),
.E(n_5348),
.Y(n_19463)
);

OR2x6_ASAP7_75t_L g19464 ( 
.A(n_19370),
.B(n_5386),
.Y(n_19464)
);

NOR3xp33_ASAP7_75t_L g19465 ( 
.A(n_19373),
.B(n_5697),
.C(n_5830),
.Y(n_19465)
);

AND5x1_ASAP7_75t_L g19466 ( 
.A(n_19349),
.B(n_6575),
.C(n_8809),
.D(n_8790),
.E(n_8146),
.Y(n_19466)
);

INVx1_ASAP7_75t_L g19467 ( 
.A(n_19345),
.Y(n_19467)
);

INVx1_ASAP7_75t_L g19468 ( 
.A(n_19374),
.Y(n_19468)
);

NAND2xp5_ASAP7_75t_SL g19469 ( 
.A(n_19396),
.B(n_7111),
.Y(n_19469)
);

INVx1_ASAP7_75t_L g19470 ( 
.A(n_19421),
.Y(n_19470)
);

AND3x4_ASAP7_75t_L g19471 ( 
.A(n_19424),
.B(n_19412),
.C(n_19398),
.Y(n_19471)
);

AND4x1_ASAP7_75t_L g19472 ( 
.A(n_19426),
.B(n_7269),
.C(n_7273),
.D(n_7265),
.Y(n_19472)
);

NAND3xp33_ASAP7_75t_SL g19473 ( 
.A(n_19410),
.B(n_5697),
.C(n_5830),
.Y(n_19473)
);

NOR3x1_ASAP7_75t_L g19474 ( 
.A(n_19425),
.B(n_8011),
.C(n_8140),
.Y(n_19474)
);

INVx1_ASAP7_75t_SL g19475 ( 
.A(n_19408),
.Y(n_19475)
);

NAND2xp5_ASAP7_75t_L g19476 ( 
.A(n_19397),
.B(n_19384),
.Y(n_19476)
);

NOR3xp33_ASAP7_75t_SL g19477 ( 
.A(n_19386),
.B(n_7269),
.C(n_7265),
.Y(n_19477)
);

AND4x1_ASAP7_75t_L g19478 ( 
.A(n_19382),
.B(n_7275),
.C(n_7286),
.D(n_7273),
.Y(n_19478)
);

INVx2_ASAP7_75t_L g19479 ( 
.A(n_19372),
.Y(n_19479)
);

NOR3xp33_ASAP7_75t_L g19480 ( 
.A(n_19423),
.B(n_5697),
.C(n_5830),
.Y(n_19480)
);

NAND2xp5_ASAP7_75t_SL g19481 ( 
.A(n_19401),
.B(n_7111),
.Y(n_19481)
);

INVx2_ASAP7_75t_SL g19482 ( 
.A(n_19431),
.Y(n_19482)
);

OAI221xp5_ASAP7_75t_L g19483 ( 
.A1(n_19379),
.A2(n_5386),
.B1(n_5881),
.B2(n_6114),
.C(n_6017),
.Y(n_19483)
);

NAND2xp5_ASAP7_75t_L g19484 ( 
.A(n_19419),
.B(n_6853),
.Y(n_19484)
);

NAND4xp25_ASAP7_75t_L g19485 ( 
.A(n_19367),
.B(n_5899),
.C(n_5908),
.D(n_5890),
.Y(n_19485)
);

NAND5xp2_ASAP7_75t_L g19486 ( 
.A(n_19375),
.B(n_4581),
.C(n_4604),
.D(n_4592),
.E(n_4578),
.Y(n_19486)
);

NAND4xp25_ASAP7_75t_L g19487 ( 
.A(n_19355),
.B(n_5899),
.C(n_5908),
.D(n_5890),
.Y(n_19487)
);

NAND4xp25_ASAP7_75t_L g19488 ( 
.A(n_19377),
.B(n_5908),
.C(n_5934),
.D(n_5899),
.Y(n_19488)
);

AND4x1_ASAP7_75t_L g19489 ( 
.A(n_19387),
.B(n_7286),
.C(n_7302),
.D(n_7275),
.Y(n_19489)
);

INVx1_ASAP7_75t_SL g19490 ( 
.A(n_19378),
.Y(n_19490)
);

INVx1_ASAP7_75t_L g19491 ( 
.A(n_19394),
.Y(n_19491)
);

NOR2xp33_ASAP7_75t_L g19492 ( 
.A(n_19406),
.B(n_6640),
.Y(n_19492)
);

NAND4xp25_ASAP7_75t_SL g19493 ( 
.A(n_19418),
.B(n_7302),
.C(n_7357),
.D(n_7275),
.Y(n_19493)
);

AOI22xp5_ASAP7_75t_SL g19494 ( 
.A1(n_19389),
.A2(n_4748),
.B1(n_4608),
.B2(n_4552),
.Y(n_19494)
);

AND3x2_ASAP7_75t_L g19495 ( 
.A(n_19404),
.B(n_4581),
.C(n_4578),
.Y(n_19495)
);

NAND4xp25_ASAP7_75t_L g19496 ( 
.A(n_19362),
.B(n_5908),
.C(n_5934),
.D(n_5899),
.Y(n_19496)
);

NAND4xp25_ASAP7_75t_L g19497 ( 
.A(n_19391),
.B(n_6017),
.C(n_6087),
.D(n_5934),
.Y(n_19497)
);

NAND3xp33_ASAP7_75t_SL g19498 ( 
.A(n_19383),
.B(n_5862),
.C(n_5861),
.Y(n_19498)
);

NOR2xp67_ASAP7_75t_L g19499 ( 
.A(n_19428),
.B(n_5862),
.Y(n_19499)
);

AND2x4_ASAP7_75t_L g19500 ( 
.A(n_19392),
.B(n_6692),
.Y(n_19500)
);

NOR2x1_ASAP7_75t_L g19501 ( 
.A(n_19427),
.B(n_6461),
.Y(n_19501)
);

NOR2xp33_ASAP7_75t_L g19502 ( 
.A(n_19409),
.B(n_6640),
.Y(n_19502)
);

AND2x4_ASAP7_75t_L g19503 ( 
.A(n_19380),
.B(n_6704),
.Y(n_19503)
);

INVx2_ASAP7_75t_L g19504 ( 
.A(n_19376),
.Y(n_19504)
);

NOR3xp33_ASAP7_75t_L g19505 ( 
.A(n_19395),
.B(n_5862),
.C(n_5861),
.Y(n_19505)
);

NAND3xp33_ASAP7_75t_SL g19506 ( 
.A(n_19430),
.B(n_5862),
.C(n_5861),
.Y(n_19506)
);

AOI22xp5_ASAP7_75t_L g19507 ( 
.A1(n_19413),
.A2(n_7136),
.B1(n_7141),
.B2(n_7111),
.Y(n_19507)
);

INVx1_ASAP7_75t_L g19508 ( 
.A(n_19358),
.Y(n_19508)
);

NOR2x1_ASAP7_75t_L g19509 ( 
.A(n_19414),
.B(n_19366),
.Y(n_19509)
);

NOR5xp2_ASAP7_75t_L g19510 ( 
.A(n_19435),
.B(n_7248),
.C(n_7251),
.D(n_7237),
.E(n_7232),
.Y(n_19510)
);

NOR3xp33_ASAP7_75t_L g19511 ( 
.A(n_19402),
.B(n_5862),
.C(n_5861),
.Y(n_19511)
);

NAND3xp33_ASAP7_75t_SL g19512 ( 
.A(n_19399),
.B(n_5886),
.C(n_5861),
.Y(n_19512)
);

NAND3xp33_ASAP7_75t_L g19513 ( 
.A(n_19403),
.B(n_7136),
.C(n_7111),
.Y(n_19513)
);

AND5x1_ASAP7_75t_L g19514 ( 
.A(n_19417),
.B(n_8809),
.C(n_8790),
.D(n_8150),
.E(n_8168),
.Y(n_19514)
);

XNOR2xp5_ASAP7_75t_L g19515 ( 
.A(n_19356),
.B(n_5934),
.Y(n_19515)
);

NAND4xp25_ASAP7_75t_L g19516 ( 
.A(n_19369),
.B(n_6087),
.C(n_6114),
.D(n_6017),
.Y(n_19516)
);

NOR3xp33_ASAP7_75t_SL g19517 ( 
.A(n_19420),
.B(n_19416),
.C(n_19365),
.Y(n_19517)
);

AND2x4_ASAP7_75t_L g19518 ( 
.A(n_19435),
.B(n_6704),
.Y(n_19518)
);

NAND3xp33_ASAP7_75t_SL g19519 ( 
.A(n_19407),
.B(n_5914),
.C(n_5886),
.Y(n_19519)
);

NOR3xp33_ASAP7_75t_L g19520 ( 
.A(n_19381),
.B(n_19393),
.C(n_5914),
.Y(n_19520)
);

NOR4xp25_ASAP7_75t_L g19521 ( 
.A(n_19433),
.B(n_7294),
.C(n_7300),
.D(n_7287),
.Y(n_19521)
);

NOR3xp33_ASAP7_75t_L g19522 ( 
.A(n_19433),
.B(n_5914),
.C(n_5886),
.Y(n_19522)
);

NOR5xp2_ASAP7_75t_L g19523 ( 
.A(n_19433),
.B(n_7267),
.C(n_7268),
.D(n_7251),
.E(n_7248),
.Y(n_19523)
);

HB1xp67_ASAP7_75t_L g19524 ( 
.A(n_19468),
.Y(n_19524)
);

AOI221x1_ASAP7_75t_L g19525 ( 
.A1(n_19491),
.A2(n_7300),
.B1(n_7308),
.B2(n_7294),
.C(n_7287),
.Y(n_19525)
);

AOI21xp5_ASAP7_75t_SL g19526 ( 
.A1(n_19482),
.A2(n_5914),
.B(n_5886),
.Y(n_19526)
);

OAI22xp5_ASAP7_75t_L g19527 ( 
.A1(n_19454),
.A2(n_7141),
.B1(n_7147),
.B2(n_7136),
.Y(n_19527)
);

INVx1_ASAP7_75t_L g19528 ( 
.A(n_19448),
.Y(n_19528)
);

AND4x1_ASAP7_75t_L g19529 ( 
.A(n_19467),
.B(n_7357),
.C(n_7361),
.D(n_7302),
.Y(n_19529)
);

NOR3xp33_ASAP7_75t_L g19530 ( 
.A(n_19470),
.B(n_5914),
.C(n_5886),
.Y(n_19530)
);

OR2x2_ASAP7_75t_L g19531 ( 
.A(n_19443),
.B(n_8809),
.Y(n_19531)
);

NAND5xp2_ASAP7_75t_L g19532 ( 
.A(n_19492),
.B(n_4581),
.C(n_4604),
.D(n_4592),
.E(n_4578),
.Y(n_19532)
);

INVx1_ASAP7_75t_L g19533 ( 
.A(n_19448),
.Y(n_19533)
);

AOI211xp5_ASAP7_75t_L g19534 ( 
.A1(n_19475),
.A2(n_8146),
.B(n_8150),
.C(n_8142),
.Y(n_19534)
);

NAND3xp33_ASAP7_75t_SL g19535 ( 
.A(n_19490),
.B(n_5959),
.C(n_6461),
.Y(n_19535)
);

OAI311xp33_ASAP7_75t_L g19536 ( 
.A1(n_19476),
.A2(n_7610),
.A3(n_7294),
.B1(n_7312),
.C1(n_7308),
.Y(n_19536)
);

OAI22xp33_ASAP7_75t_L g19537 ( 
.A1(n_19461),
.A2(n_7136),
.B1(n_7147),
.B2(n_7141),
.Y(n_19537)
);

AO22x1_ASAP7_75t_L g19538 ( 
.A1(n_19471),
.A2(n_4748),
.B1(n_4608),
.B2(n_5431),
.Y(n_19538)
);

NAND5xp2_ASAP7_75t_L g19539 ( 
.A(n_19453),
.B(n_19517),
.C(n_19507),
.D(n_19451),
.E(n_19508),
.Y(n_19539)
);

INVx1_ASAP7_75t_L g19540 ( 
.A(n_19458),
.Y(n_19540)
);

NAND3xp33_ASAP7_75t_SL g19541 ( 
.A(n_19504),
.B(n_19479),
.C(n_19469),
.Y(n_19541)
);

NOR3x1_ASAP7_75t_L g19542 ( 
.A(n_19481),
.B(n_8011),
.C(n_8601),
.Y(n_19542)
);

NAND4xp25_ASAP7_75t_L g19543 ( 
.A(n_19509),
.B(n_6017),
.C(n_6114),
.D(n_6087),
.Y(n_19543)
);

OA211x2_ASAP7_75t_L g19544 ( 
.A1(n_19502),
.A2(n_7361),
.B(n_7362),
.C(n_7357),
.Y(n_19544)
);

NAND2xp5_ASAP7_75t_L g19545 ( 
.A(n_19500),
.B(n_19447),
.Y(n_19545)
);

AND4x1_ASAP7_75t_L g19546 ( 
.A(n_19438),
.B(n_7362),
.C(n_7375),
.D(n_7361),
.Y(n_19546)
);

OAI211xp5_ASAP7_75t_SL g19547 ( 
.A1(n_19484),
.A2(n_7308),
.B(n_7312),
.C(n_7300),
.Y(n_19547)
);

INVx1_ASAP7_75t_L g19548 ( 
.A(n_19499),
.Y(n_19548)
);

OAI211xp5_ASAP7_75t_L g19549 ( 
.A1(n_19511),
.A2(n_6474),
.B(n_6508),
.C(n_6481),
.Y(n_19549)
);

AOI22xp5_ASAP7_75t_L g19550 ( 
.A1(n_19500),
.A2(n_19503),
.B1(n_19520),
.B2(n_19456),
.Y(n_19550)
);

AO22x1_ASAP7_75t_L g19551 ( 
.A1(n_19442),
.A2(n_19444),
.B1(n_19501),
.B2(n_19503),
.Y(n_19551)
);

INVx1_ASAP7_75t_L g19552 ( 
.A(n_19441),
.Y(n_19552)
);

INVx1_ASAP7_75t_L g19553 ( 
.A(n_19515),
.Y(n_19553)
);

INVx1_ASAP7_75t_L g19554 ( 
.A(n_19518),
.Y(n_19554)
);

NAND2xp5_ASAP7_75t_SL g19555 ( 
.A(n_19522),
.B(n_7136),
.Y(n_19555)
);

NOR4xp25_ASAP7_75t_L g19556 ( 
.A(n_19498),
.B(n_7308),
.C(n_7312),
.D(n_7300),
.Y(n_19556)
);

OAI222xp33_ASAP7_75t_L g19557 ( 
.A1(n_19464),
.A2(n_7290),
.B1(n_7254),
.B2(n_7303),
.C1(n_7262),
.C2(n_7225),
.Y(n_19557)
);

OAI221xp5_ASAP7_75t_L g19558 ( 
.A1(n_19436),
.A2(n_6087),
.B1(n_6178),
.B2(n_6117),
.C(n_6114),
.Y(n_19558)
);

NAND2xp5_ASAP7_75t_L g19559 ( 
.A(n_19495),
.B(n_6911),
.Y(n_19559)
);

NAND5xp2_ASAP7_75t_L g19560 ( 
.A(n_19465),
.B(n_4604),
.C(n_4625),
.D(n_4622),
.E(n_4592),
.Y(n_19560)
);

OAI221xp5_ASAP7_75t_L g19561 ( 
.A1(n_19497),
.A2(n_6117),
.B1(n_6326),
.B2(n_6233),
.C(n_6178),
.Y(n_19561)
);

AOI22xp5_ASAP7_75t_L g19562 ( 
.A1(n_19480),
.A2(n_7431),
.B1(n_7437),
.B2(n_7350),
.Y(n_19562)
);

NOR3xp33_ASAP7_75t_L g19563 ( 
.A(n_19519),
.B(n_5959),
.C(n_6474),
.Y(n_19563)
);

NAND2xp5_ASAP7_75t_SL g19564 ( 
.A(n_19518),
.B(n_7136),
.Y(n_19564)
);

AOI22xp5_ASAP7_75t_L g19565 ( 
.A1(n_19488),
.A2(n_7304),
.B1(n_7515),
.B2(n_7282),
.Y(n_19565)
);

AO22x2_ASAP7_75t_L g19566 ( 
.A1(n_19512),
.A2(n_7312),
.B1(n_7313),
.B2(n_7308),
.Y(n_19566)
);

OAI211xp5_ASAP7_75t_L g19567 ( 
.A1(n_19487),
.A2(n_6474),
.B(n_6508),
.C(n_6481),
.Y(n_19567)
);

NAND2xp5_ASAP7_75t_L g19568 ( 
.A(n_19477),
.B(n_6911),
.Y(n_19568)
);

NAND3xp33_ASAP7_75t_SL g19569 ( 
.A(n_19446),
.B(n_5959),
.C(n_6474),
.Y(n_19569)
);

NOR2x1_ASAP7_75t_L g19570 ( 
.A(n_19506),
.B(n_19464),
.Y(n_19570)
);

AOI22xp5_ASAP7_75t_L g19571 ( 
.A1(n_19473),
.A2(n_7304),
.B1(n_7515),
.B2(n_7282),
.Y(n_19571)
);

AO22x2_ASAP7_75t_L g19572 ( 
.A1(n_19440),
.A2(n_7312),
.B1(n_7313),
.B2(n_7308),
.Y(n_19572)
);

XOR2xp5_ASAP7_75t_L g19573 ( 
.A(n_19493),
.B(n_4819),
.Y(n_19573)
);

OAI211xp5_ASAP7_75t_L g19574 ( 
.A1(n_19516),
.A2(n_6474),
.B(n_6508),
.C(n_6481),
.Y(n_19574)
);

NAND4xp25_ASAP7_75t_L g19575 ( 
.A(n_19463),
.B(n_6117),
.C(n_6233),
.D(n_6178),
.Y(n_19575)
);

AOI22xp33_ASAP7_75t_L g19576 ( 
.A1(n_19505),
.A2(n_7141),
.B1(n_7169),
.B2(n_7147),
.Y(n_19576)
);

AOI21xp5_ASAP7_75t_L g19577 ( 
.A1(n_19486),
.A2(n_5799),
.B(n_8011),
.Y(n_19577)
);

INVx1_ASAP7_75t_L g19578 ( 
.A(n_19513),
.Y(n_19578)
);

NOR2x1_ASAP7_75t_L g19579 ( 
.A(n_19496),
.B(n_6481),
.Y(n_19579)
);

INVx1_ASAP7_75t_SL g19580 ( 
.A(n_19455),
.Y(n_19580)
);

INVx1_ASAP7_75t_L g19581 ( 
.A(n_19489),
.Y(n_19581)
);

NOR3xp33_ASAP7_75t_L g19582 ( 
.A(n_19483),
.B(n_5959),
.C(n_6481),
.Y(n_19582)
);

NAND3xp33_ASAP7_75t_L g19583 ( 
.A(n_19449),
.B(n_5431),
.C(n_7141),
.Y(n_19583)
);

OAI211xp5_ASAP7_75t_L g19584 ( 
.A1(n_19521),
.A2(n_6508),
.B(n_6521),
.C(n_6517),
.Y(n_19584)
);

NAND3xp33_ASAP7_75t_L g19585 ( 
.A(n_19485),
.B(n_5431),
.C(n_7147),
.Y(n_19585)
);

NAND4xp25_ASAP7_75t_L g19586 ( 
.A(n_19437),
.B(n_6117),
.C(n_6233),
.D(n_6178),
.Y(n_19586)
);

NAND3xp33_ASAP7_75t_SL g19587 ( 
.A(n_19510),
.B(n_5959),
.C(n_6508),
.Y(n_19587)
);

AND5x1_ASAP7_75t_L g19588 ( 
.A(n_19450),
.B(n_19466),
.C(n_19445),
.D(n_19457),
.E(n_19514),
.Y(n_19588)
);

INVx2_ASAP7_75t_L g19589 ( 
.A(n_19459),
.Y(n_19589)
);

NAND4xp25_ASAP7_75t_L g19590 ( 
.A(n_19494),
.B(n_6326),
.C(n_6328),
.D(n_6233),
.Y(n_19590)
);

AND2x2_ASAP7_75t_L g19591 ( 
.A(n_19472),
.B(n_19478),
.Y(n_19591)
);

OAI22xp5_ASAP7_75t_L g19592 ( 
.A1(n_19452),
.A2(n_7169),
.B1(n_7175),
.B2(n_7147),
.Y(n_19592)
);

INVx1_ASAP7_75t_L g19593 ( 
.A(n_19439),
.Y(n_19593)
);

INVx1_ASAP7_75t_L g19594 ( 
.A(n_19474),
.Y(n_19594)
);

NAND4xp25_ASAP7_75t_L g19595 ( 
.A(n_19462),
.B(n_19523),
.C(n_19460),
.D(n_6328),
.Y(n_19595)
);

NAND5xp2_ASAP7_75t_L g19596 ( 
.A(n_19454),
.B(n_4622),
.C(n_4655),
.D(n_4631),
.E(n_4625),
.Y(n_19596)
);

OAI22xp5_ASAP7_75t_L g19597 ( 
.A1(n_19524),
.A2(n_7169),
.B1(n_7175),
.B2(n_7147),
.Y(n_19597)
);

BUFx2_ASAP7_75t_L g19598 ( 
.A(n_19528),
.Y(n_19598)
);

NOR2xp33_ASAP7_75t_L g19599 ( 
.A(n_19533),
.B(n_6640),
.Y(n_19599)
);

AND3x2_ASAP7_75t_L g19600 ( 
.A(n_19554),
.B(n_4625),
.C(n_4622),
.Y(n_19600)
);

AO22x2_ASAP7_75t_L g19601 ( 
.A1(n_19540),
.A2(n_7317),
.B1(n_7327),
.B2(n_7313),
.Y(n_19601)
);

OAI22xp5_ASAP7_75t_L g19602 ( 
.A1(n_19545),
.A2(n_7175),
.B1(n_7206),
.B2(n_7169),
.Y(n_19602)
);

AOI221xp5_ASAP7_75t_L g19603 ( 
.A1(n_19594),
.A2(n_7175),
.B1(n_7221),
.B2(n_7206),
.C(n_7169),
.Y(n_19603)
);

XOR2x1_ASAP7_75t_L g19604 ( 
.A(n_19553),
.B(n_4785),
.Y(n_19604)
);

AOI22xp5_ASAP7_75t_L g19605 ( 
.A1(n_19541),
.A2(n_7175),
.B1(n_7206),
.B2(n_7169),
.Y(n_19605)
);

NAND2xp5_ASAP7_75t_L g19606 ( 
.A(n_19591),
.B(n_19581),
.Y(n_19606)
);

OAI22xp5_ASAP7_75t_L g19607 ( 
.A1(n_19589),
.A2(n_7206),
.B1(n_7221),
.B2(n_7169),
.Y(n_19607)
);

HB1xp67_ASAP7_75t_L g19608 ( 
.A(n_19570),
.Y(n_19608)
);

OAI22xp5_ASAP7_75t_L g19609 ( 
.A1(n_19550),
.A2(n_7206),
.B1(n_7221),
.B2(n_7169),
.Y(n_19609)
);

INVxp67_ASAP7_75t_L g19610 ( 
.A(n_19539),
.Y(n_19610)
);

INVx3_ASAP7_75t_SL g19611 ( 
.A(n_19580),
.Y(n_19611)
);

NAND2xp5_ASAP7_75t_L g19612 ( 
.A(n_19593),
.B(n_6911),
.Y(n_19612)
);

INVx1_ASAP7_75t_SL g19613 ( 
.A(n_19552),
.Y(n_19613)
);

INVx2_ASAP7_75t_SL g19614 ( 
.A(n_19548),
.Y(n_19614)
);

INVx1_ASAP7_75t_L g19615 ( 
.A(n_19551),
.Y(n_19615)
);

NOR2xp67_ASAP7_75t_L g19616 ( 
.A(n_19578),
.B(n_6517),
.Y(n_19616)
);

OAI321xp33_ASAP7_75t_L g19617 ( 
.A1(n_19585),
.A2(n_7206),
.A3(n_7277),
.B1(n_7304),
.B2(n_7282),
.C(n_7221),
.Y(n_19617)
);

OAI22xp5_ASAP7_75t_L g19618 ( 
.A1(n_19573),
.A2(n_7221),
.B1(n_7277),
.B2(n_7206),
.Y(n_19618)
);

OAI21xp5_ASAP7_75t_L g19619 ( 
.A1(n_19579),
.A2(n_8168),
.B(n_8150),
.Y(n_19619)
);

NAND4xp25_ASAP7_75t_L g19620 ( 
.A(n_19532),
.B(n_6328),
.C(n_6334),
.D(n_6326),
.Y(n_19620)
);

OR2x2_ASAP7_75t_L g19621 ( 
.A(n_19568),
.B(n_8809),
.Y(n_19621)
);

AOI21xp33_ASAP7_75t_L g19622 ( 
.A1(n_19583),
.A2(n_5799),
.B(n_5431),
.Y(n_19622)
);

INVx2_ASAP7_75t_SL g19623 ( 
.A(n_19564),
.Y(n_19623)
);

AOI22xp5_ASAP7_75t_L g19624 ( 
.A1(n_19530),
.A2(n_7304),
.B1(n_7347),
.B2(n_7277),
.Y(n_19624)
);

NAND4xp25_ASAP7_75t_L g19625 ( 
.A(n_19575),
.B(n_6328),
.C(n_6334),
.D(n_6326),
.Y(n_19625)
);

NOR2xp33_ASAP7_75t_L g19626 ( 
.A(n_19559),
.B(n_6640),
.Y(n_19626)
);

NAND2xp5_ASAP7_75t_SL g19627 ( 
.A(n_19556),
.B(n_7277),
.Y(n_19627)
);

INVx1_ASAP7_75t_L g19628 ( 
.A(n_19595),
.Y(n_19628)
);

INVx2_ASAP7_75t_L g19629 ( 
.A(n_19566),
.Y(n_19629)
);

INVx2_ASAP7_75t_L g19630 ( 
.A(n_19566),
.Y(n_19630)
);

INVx1_ASAP7_75t_L g19631 ( 
.A(n_19569),
.Y(n_19631)
);

INVx2_ASAP7_75t_L g19632 ( 
.A(n_19572),
.Y(n_19632)
);

XNOR2xp5_ASAP7_75t_L g19633 ( 
.A(n_19590),
.B(n_6419),
.Y(n_19633)
);

NAND2xp5_ASAP7_75t_L g19634 ( 
.A(n_19555),
.B(n_6911),
.Y(n_19634)
);

HB1xp67_ASAP7_75t_L g19635 ( 
.A(n_19588),
.Y(n_19635)
);

HB1xp67_ASAP7_75t_L g19636 ( 
.A(n_19572),
.Y(n_19636)
);

NAND2xp33_ASAP7_75t_SL g19637 ( 
.A(n_19531),
.B(n_5314),
.Y(n_19637)
);

OA22x2_ASAP7_75t_L g19638 ( 
.A1(n_19567),
.A2(n_8173),
.B1(n_8175),
.B2(n_8168),
.Y(n_19638)
);

INVx2_ASAP7_75t_L g19639 ( 
.A(n_19561),
.Y(n_19639)
);

AND3x1_ASAP7_75t_L g19640 ( 
.A(n_19563),
.B(n_7375),
.C(n_7362),
.Y(n_19640)
);

AOI22xp5_ASAP7_75t_L g19641 ( 
.A1(n_19582),
.A2(n_7304),
.B1(n_7347),
.B2(n_7277),
.Y(n_19641)
);

INVx1_ASAP7_75t_L g19642 ( 
.A(n_19586),
.Y(n_19642)
);

NOR2x1_ASAP7_75t_L g19643 ( 
.A(n_19535),
.B(n_6517),
.Y(n_19643)
);

NOR3xp33_ASAP7_75t_L g19644 ( 
.A(n_19549),
.B(n_6521),
.C(n_6517),
.Y(n_19644)
);

XNOR2xp5_ASAP7_75t_L g19645 ( 
.A(n_19544),
.B(n_6435),
.Y(n_19645)
);

NAND2xp5_ASAP7_75t_L g19646 ( 
.A(n_19574),
.B(n_6916),
.Y(n_19646)
);

OAI22xp5_ASAP7_75t_SL g19647 ( 
.A1(n_19558),
.A2(n_6517),
.B1(n_6552),
.B2(n_6521),
.Y(n_19647)
);

NOR3xp33_ASAP7_75t_SL g19648 ( 
.A(n_19560),
.B(n_7378),
.C(n_7375),
.Y(n_19648)
);

AOI21xp5_ASAP7_75t_L g19649 ( 
.A1(n_19526),
.A2(n_6604),
.B(n_6576),
.Y(n_19649)
);

INVx4_ASAP7_75t_L g19650 ( 
.A(n_19596),
.Y(n_19650)
);

INVx1_ASAP7_75t_L g19651 ( 
.A(n_19547),
.Y(n_19651)
);

INVx1_ASAP7_75t_L g19652 ( 
.A(n_19584),
.Y(n_19652)
);

OAI22xp5_ASAP7_75t_L g19653 ( 
.A1(n_19576),
.A2(n_7304),
.B1(n_7347),
.B2(n_7277),
.Y(n_19653)
);

OAI211xp5_ASAP7_75t_SL g19654 ( 
.A1(n_19577),
.A2(n_19565),
.B(n_19571),
.C(n_19527),
.Y(n_19654)
);

NAND4xp25_ASAP7_75t_L g19655 ( 
.A(n_19543),
.B(n_6336),
.C(n_6340),
.D(n_6334),
.Y(n_19655)
);

INVx1_ASAP7_75t_L g19656 ( 
.A(n_19525),
.Y(n_19656)
);

OA22x2_ASAP7_75t_L g19657 ( 
.A1(n_19562),
.A2(n_8175),
.B1(n_8176),
.B2(n_8173),
.Y(n_19657)
);

INVx1_ASAP7_75t_L g19658 ( 
.A(n_19608),
.Y(n_19658)
);

NAND2xp5_ASAP7_75t_SL g19659 ( 
.A(n_19615),
.B(n_19537),
.Y(n_19659)
);

AND2x4_ASAP7_75t_L g19660 ( 
.A(n_19598),
.B(n_19546),
.Y(n_19660)
);

INVx2_ASAP7_75t_L g19661 ( 
.A(n_19614),
.Y(n_19661)
);

INVx1_ASAP7_75t_L g19662 ( 
.A(n_19635),
.Y(n_19662)
);

INVx1_ASAP7_75t_L g19663 ( 
.A(n_19606),
.Y(n_19663)
);

AND3x4_ASAP7_75t_L g19664 ( 
.A(n_19639),
.B(n_19529),
.C(n_19536),
.Y(n_19664)
);

OR3x1_ASAP7_75t_L g19665 ( 
.A(n_19628),
.B(n_19587),
.C(n_19538),
.Y(n_19665)
);

INVx1_ASAP7_75t_L g19666 ( 
.A(n_19636),
.Y(n_19666)
);

AOI22x1_ASAP7_75t_L g19667 ( 
.A1(n_19613),
.A2(n_19592),
.B1(n_19557),
.B2(n_19542),
.Y(n_19667)
);

NAND2xp5_ASAP7_75t_L g19668 ( 
.A(n_19604),
.B(n_19534),
.Y(n_19668)
);

INVx1_ASAP7_75t_L g19669 ( 
.A(n_19656),
.Y(n_19669)
);

INVx1_ASAP7_75t_L g19670 ( 
.A(n_19610),
.Y(n_19670)
);

INVx4_ASAP7_75t_L g19671 ( 
.A(n_19611),
.Y(n_19671)
);

INVx1_ASAP7_75t_L g19672 ( 
.A(n_19651),
.Y(n_19672)
);

OAI22x1_ASAP7_75t_L g19673 ( 
.A1(n_19642),
.A2(n_19623),
.B1(n_19631),
.B2(n_19652),
.Y(n_19673)
);

INVxp67_ASAP7_75t_L g19674 ( 
.A(n_19629),
.Y(n_19674)
);

OAI22xp5_ASAP7_75t_L g19675 ( 
.A1(n_19599),
.A2(n_7304),
.B1(n_7347),
.B2(n_7277),
.Y(n_19675)
);

NAND2xp5_ASAP7_75t_L g19676 ( 
.A(n_19650),
.B(n_6916),
.Y(n_19676)
);

INVx1_ASAP7_75t_L g19677 ( 
.A(n_19630),
.Y(n_19677)
);

INVx1_ASAP7_75t_L g19678 ( 
.A(n_19632),
.Y(n_19678)
);

INVx1_ASAP7_75t_L g19679 ( 
.A(n_19637),
.Y(n_19679)
);

INVxp67_ASAP7_75t_L g19680 ( 
.A(n_19626),
.Y(n_19680)
);

XOR2xp5_ASAP7_75t_L g19681 ( 
.A(n_19633),
.B(n_4819),
.Y(n_19681)
);

XOR2xp5_ASAP7_75t_L g19682 ( 
.A(n_19612),
.B(n_4819),
.Y(n_19682)
);

XOR2xp5_ASAP7_75t_L g19683 ( 
.A(n_19645),
.B(n_4819),
.Y(n_19683)
);

INVx1_ASAP7_75t_L g19684 ( 
.A(n_19654),
.Y(n_19684)
);

INVx3_ASAP7_75t_SL g19685 ( 
.A(n_19621),
.Y(n_19685)
);

INVx1_ASAP7_75t_L g19686 ( 
.A(n_19643),
.Y(n_19686)
);

INVx1_ASAP7_75t_L g19687 ( 
.A(n_19634),
.Y(n_19687)
);

INVx1_ASAP7_75t_L g19688 ( 
.A(n_19627),
.Y(n_19688)
);

AOI22xp5_ASAP7_75t_L g19689 ( 
.A1(n_19625),
.A2(n_7304),
.B1(n_7347),
.B2(n_7277),
.Y(n_19689)
);

INVx2_ASAP7_75t_L g19690 ( 
.A(n_19646),
.Y(n_19690)
);

AO22x2_ASAP7_75t_L g19691 ( 
.A1(n_19649),
.A2(n_7317),
.B1(n_7333),
.B2(n_7313),
.Y(n_19691)
);

XNOR2xp5_ASAP7_75t_L g19692 ( 
.A(n_19648),
.B(n_19620),
.Y(n_19692)
);

INVx1_ASAP7_75t_L g19693 ( 
.A(n_19616),
.Y(n_19693)
);

INVx1_ASAP7_75t_L g19694 ( 
.A(n_19640),
.Y(n_19694)
);

INVx1_ASAP7_75t_L g19695 ( 
.A(n_19617),
.Y(n_19695)
);

INVx1_ASAP7_75t_L g19696 ( 
.A(n_19655),
.Y(n_19696)
);

INVx2_ASAP7_75t_L g19697 ( 
.A(n_19600),
.Y(n_19697)
);

AOI22x1_ASAP7_75t_L g19698 ( 
.A1(n_19622),
.A2(n_6552),
.B1(n_6556),
.B2(n_6521),
.Y(n_19698)
);

AND2x4_ASAP7_75t_L g19699 ( 
.A(n_19605),
.B(n_6704),
.Y(n_19699)
);

INVx1_ASAP7_75t_L g19700 ( 
.A(n_19647),
.Y(n_19700)
);

OAI22xp5_ASAP7_75t_SL g19701 ( 
.A1(n_19658),
.A2(n_19641),
.B1(n_19602),
.B2(n_19609),
.Y(n_19701)
);

NAND5xp2_ASAP7_75t_L g19702 ( 
.A(n_19662),
.B(n_19644),
.C(n_19619),
.D(n_19603),
.E(n_19624),
.Y(n_19702)
);

INVx1_ASAP7_75t_L g19703 ( 
.A(n_19666),
.Y(n_19703)
);

OAI22xp5_ASAP7_75t_SL g19704 ( 
.A1(n_19671),
.A2(n_19607),
.B1(n_19597),
.B2(n_19618),
.Y(n_19704)
);

INVx1_ASAP7_75t_L g19705 ( 
.A(n_19663),
.Y(n_19705)
);

OAI31xp67_ASAP7_75t_L g19706 ( 
.A1(n_19661),
.A2(n_19638),
.A3(n_19601),
.B(n_19653),
.Y(n_19706)
);

AND3x1_ASAP7_75t_L g19707 ( 
.A(n_19677),
.B(n_19601),
.C(n_19657),
.Y(n_19707)
);

INVx1_ASAP7_75t_L g19708 ( 
.A(n_19670),
.Y(n_19708)
);

INVx1_ASAP7_75t_L g19709 ( 
.A(n_19669),
.Y(n_19709)
);

OAI22xp5_ASAP7_75t_SL g19710 ( 
.A1(n_19674),
.A2(n_6521),
.B1(n_6556),
.B2(n_6552),
.Y(n_19710)
);

NAND4xp75_ASAP7_75t_L g19711 ( 
.A(n_19678),
.B(n_7378),
.C(n_5325),
.D(n_7190),
.Y(n_19711)
);

HB1xp67_ASAP7_75t_L g19712 ( 
.A(n_19665),
.Y(n_19712)
);

INVx2_ASAP7_75t_L g19713 ( 
.A(n_19667),
.Y(n_19713)
);

AND3x1_ASAP7_75t_L g19714 ( 
.A(n_19684),
.B(n_4818),
.C(n_4614),
.Y(n_19714)
);

INVx1_ASAP7_75t_SL g19715 ( 
.A(n_19660),
.Y(n_19715)
);

XNOR2xp5_ASAP7_75t_L g19716 ( 
.A(n_19673),
.B(n_6334),
.Y(n_19716)
);

INVx1_ASAP7_75t_L g19717 ( 
.A(n_19692),
.Y(n_19717)
);

OA21x2_ASAP7_75t_L g19718 ( 
.A1(n_19688),
.A2(n_8175),
.B(n_8173),
.Y(n_19718)
);

INVx1_ASAP7_75t_SL g19719 ( 
.A(n_19685),
.Y(n_19719)
);

OAI22xp5_ASAP7_75t_L g19720 ( 
.A1(n_19664),
.A2(n_19676),
.B1(n_19672),
.B2(n_19694),
.Y(n_19720)
);

INVx3_ASAP7_75t_L g19721 ( 
.A(n_19697),
.Y(n_19721)
);

OAI21x1_ASAP7_75t_L g19722 ( 
.A1(n_19679),
.A2(n_7944),
.B(n_7968),
.Y(n_19722)
);

NAND3xp33_ASAP7_75t_SL g19723 ( 
.A(n_19687),
.B(n_6556),
.C(n_6552),
.Y(n_19723)
);

OAI21x1_ASAP7_75t_SL g19724 ( 
.A1(n_19668),
.A2(n_7378),
.B(n_6744),
.Y(n_19724)
);

AND2x2_ASAP7_75t_L g19725 ( 
.A(n_19690),
.B(n_6640),
.Y(n_19725)
);

BUFx2_ASAP7_75t_L g19726 ( 
.A(n_19695),
.Y(n_19726)
);

OAI22xp5_ASAP7_75t_L g19727 ( 
.A1(n_19683),
.A2(n_7347),
.B1(n_7350),
.B2(n_7277),
.Y(n_19727)
);

AOI21xp5_ASAP7_75t_L g19728 ( 
.A1(n_19659),
.A2(n_6604),
.B(n_5799),
.Y(n_19728)
);

INVx2_ASAP7_75t_L g19729 ( 
.A(n_19693),
.Y(n_19729)
);

INVx1_ASAP7_75t_L g19730 ( 
.A(n_19686),
.Y(n_19730)
);

AOI22xp5_ASAP7_75t_L g19731 ( 
.A1(n_19680),
.A2(n_7350),
.B1(n_7366),
.B2(n_7347),
.Y(n_19731)
);

INVx1_ASAP7_75t_L g19732 ( 
.A(n_19696),
.Y(n_19732)
);

AO22x2_ASAP7_75t_L g19733 ( 
.A1(n_19703),
.A2(n_19700),
.B1(n_19681),
.B2(n_19682),
.Y(n_19733)
);

NAND4xp25_ASAP7_75t_L g19734 ( 
.A(n_19719),
.B(n_19699),
.C(n_19689),
.D(n_19675),
.Y(n_19734)
);

INVx1_ASAP7_75t_L g19735 ( 
.A(n_19716),
.Y(n_19735)
);

INVxp67_ASAP7_75t_L g19736 ( 
.A(n_19712),
.Y(n_19736)
);

NOR3xp33_ASAP7_75t_L g19737 ( 
.A(n_19721),
.B(n_19698),
.C(n_19691),
.Y(n_19737)
);

INVx3_ASAP7_75t_SL g19738 ( 
.A(n_19715),
.Y(n_19738)
);

OAI222xp33_ASAP7_75t_L g19739 ( 
.A1(n_19709),
.A2(n_19691),
.B1(n_5799),
.B2(n_6556),
.C1(n_6595),
.C2(n_6562),
.Y(n_19739)
);

NOR3xp33_ASAP7_75t_L g19740 ( 
.A(n_19720),
.B(n_6556),
.C(n_6552),
.Y(n_19740)
);

AOI22xp5_ASAP7_75t_L g19741 ( 
.A1(n_19705),
.A2(n_19708),
.B1(n_19730),
.B2(n_19713),
.Y(n_19741)
);

OAI321xp33_ASAP7_75t_L g19742 ( 
.A1(n_19717),
.A2(n_7371),
.A3(n_7350),
.B1(n_7431),
.B2(n_7366),
.C(n_7347),
.Y(n_19742)
);

XOR2xp5_ASAP7_75t_L g19743 ( 
.A(n_19726),
.B(n_4819),
.Y(n_19743)
);

NAND2xp5_ASAP7_75t_L g19744 ( 
.A(n_19729),
.B(n_19732),
.Y(n_19744)
);

AOI22xp5_ASAP7_75t_L g19745 ( 
.A1(n_19707),
.A2(n_7350),
.B1(n_7366),
.B2(n_7347),
.Y(n_19745)
);

INVx1_ASAP7_75t_L g19746 ( 
.A(n_19701),
.Y(n_19746)
);

INVx1_ASAP7_75t_L g19747 ( 
.A(n_19704),
.Y(n_19747)
);

NAND3x1_ASAP7_75t_L g19748 ( 
.A(n_19725),
.B(n_4818),
.C(n_4614),
.Y(n_19748)
);

AOI221xp5_ASAP7_75t_L g19749 ( 
.A1(n_19702),
.A2(n_7371),
.B1(n_7431),
.B2(n_7366),
.C(n_7350),
.Y(n_19749)
);

INVx1_ASAP7_75t_L g19750 ( 
.A(n_19706),
.Y(n_19750)
);

NOR3xp33_ASAP7_75t_L g19751 ( 
.A(n_19723),
.B(n_6595),
.C(n_6562),
.Y(n_19751)
);

OAI221xp5_ASAP7_75t_SL g19752 ( 
.A1(n_19728),
.A2(n_6350),
.B1(n_6400),
.B2(n_6340),
.C(n_6336),
.Y(n_19752)
);

NAND4xp75_ASAP7_75t_L g19753 ( 
.A(n_19714),
.B(n_5135),
.C(n_5142),
.D(n_5133),
.Y(n_19753)
);

INVx4_ASAP7_75t_L g19754 ( 
.A(n_19738),
.Y(n_19754)
);

AOI22xp5_ASAP7_75t_L g19755 ( 
.A1(n_19736),
.A2(n_19710),
.B1(n_19727),
.B2(n_19731),
.Y(n_19755)
);

OAI22xp5_ASAP7_75t_SL g19756 ( 
.A1(n_19746),
.A2(n_19724),
.B1(n_19718),
.B2(n_19711),
.Y(n_19756)
);

O2A1O1Ixp33_ASAP7_75t_L g19757 ( 
.A1(n_19744),
.A2(n_19718),
.B(n_19722),
.C(n_6340),
.Y(n_19757)
);

AOI22x1_ASAP7_75t_L g19758 ( 
.A1(n_19747),
.A2(n_6595),
.B1(n_6597),
.B2(n_6562),
.Y(n_19758)
);

INVx1_ASAP7_75t_L g19759 ( 
.A(n_19741),
.Y(n_19759)
);

INVx2_ASAP7_75t_L g19760 ( 
.A(n_19733),
.Y(n_19760)
);

XNOR2x1_ASAP7_75t_L g19761 ( 
.A(n_19750),
.B(n_6336),
.Y(n_19761)
);

INVx2_ASAP7_75t_L g19762 ( 
.A(n_19733),
.Y(n_19762)
);

INVx1_ASAP7_75t_L g19763 ( 
.A(n_19743),
.Y(n_19763)
);

INVx1_ASAP7_75t_L g19764 ( 
.A(n_19735),
.Y(n_19764)
);

AOI21xp5_ASAP7_75t_L g19765 ( 
.A1(n_19734),
.A2(n_6854),
.B(n_6807),
.Y(n_19765)
);

OAI22xp5_ASAP7_75t_L g19766 ( 
.A1(n_19737),
.A2(n_7366),
.B1(n_7371),
.B2(n_7350),
.Y(n_19766)
);

XNOR2x1_ASAP7_75t_L g19767 ( 
.A(n_19753),
.B(n_6336),
.Y(n_19767)
);

XNOR2xp5_ASAP7_75t_L g19768 ( 
.A(n_19740),
.B(n_6340),
.Y(n_19768)
);

AOI22x1_ASAP7_75t_L g19769 ( 
.A1(n_19751),
.A2(n_6597),
.B1(n_6595),
.B2(n_6562),
.Y(n_19769)
);

NAND2xp5_ASAP7_75t_L g19770 ( 
.A(n_19754),
.B(n_19745),
.Y(n_19770)
);

NOR3xp33_ASAP7_75t_L g19771 ( 
.A(n_19759),
.B(n_19752),
.C(n_19739),
.Y(n_19771)
);

OAI322xp33_ASAP7_75t_L g19772 ( 
.A1(n_19760),
.A2(n_19748),
.A3(n_19742),
.B1(n_19749),
.B2(n_6597),
.C1(n_6595),
.C2(n_7366),
.Y(n_19772)
);

NOR4xp25_ASAP7_75t_L g19773 ( 
.A(n_19762),
.B(n_7317),
.C(n_7327),
.D(n_7313),
.Y(n_19773)
);

INVx1_ASAP7_75t_L g19774 ( 
.A(n_19761),
.Y(n_19774)
);

NAND3x1_ASAP7_75t_L g19775 ( 
.A(n_19764),
.B(n_4818),
.C(n_4614),
.Y(n_19775)
);

OR2x6_ASAP7_75t_L g19776 ( 
.A(n_19763),
.B(n_6350),
.Y(n_19776)
);

NAND2xp5_ASAP7_75t_L g19777 ( 
.A(n_19755),
.B(n_6640),
.Y(n_19777)
);

INVx1_ASAP7_75t_L g19778 ( 
.A(n_19756),
.Y(n_19778)
);

XNOR2xp5_ASAP7_75t_L g19779 ( 
.A(n_19768),
.B(n_6350),
.Y(n_19779)
);

AOI22xp5_ASAP7_75t_L g19780 ( 
.A1(n_19778),
.A2(n_19767),
.B1(n_19765),
.B2(n_19766),
.Y(n_19780)
);

OAI21xp5_ASAP7_75t_L g19781 ( 
.A1(n_19770),
.A2(n_19757),
.B(n_19769),
.Y(n_19781)
);

OAI22xp5_ASAP7_75t_L g19782 ( 
.A1(n_19774),
.A2(n_19758),
.B1(n_7366),
.B2(n_7371),
.Y(n_19782)
);

OAI21xp5_ASAP7_75t_L g19783 ( 
.A1(n_19771),
.A2(n_7987),
.B(n_7968),
.Y(n_19783)
);

AO21x2_ASAP7_75t_L g19784 ( 
.A1(n_19777),
.A2(n_7944),
.B(n_7968),
.Y(n_19784)
);

OAI22xp5_ASAP7_75t_L g19785 ( 
.A1(n_19779),
.A2(n_19775),
.B1(n_19772),
.B2(n_19776),
.Y(n_19785)
);

AOI221x1_ASAP7_75t_L g19786 ( 
.A1(n_19773),
.A2(n_7317),
.B1(n_7333),
.B2(n_7327),
.C(n_7313),
.Y(n_19786)
);

INVx2_ASAP7_75t_L g19787 ( 
.A(n_19776),
.Y(n_19787)
);

INVx1_ASAP7_75t_L g19788 ( 
.A(n_19787),
.Y(n_19788)
);

AOI21xp33_ASAP7_75t_L g19789 ( 
.A1(n_19781),
.A2(n_6419),
.B(n_6400),
.Y(n_19789)
);

OAI22xp5_ASAP7_75t_L g19790 ( 
.A1(n_19780),
.A2(n_19785),
.B1(n_19782),
.B2(n_19786),
.Y(n_19790)
);

AOI21xp5_ASAP7_75t_L g19791 ( 
.A1(n_19784),
.A2(n_6854),
.B(n_6807),
.Y(n_19791)
);

INVx1_ASAP7_75t_L g19792 ( 
.A(n_19783),
.Y(n_19792)
);

OAI22xp5_ASAP7_75t_SL g19793 ( 
.A1(n_19780),
.A2(n_6597),
.B1(n_6419),
.B2(n_6435),
.Y(n_19793)
);

XNOR2xp5_ASAP7_75t_L g19794 ( 
.A(n_19788),
.B(n_6400),
.Y(n_19794)
);

OR2x6_ASAP7_75t_L g19795 ( 
.A(n_19790),
.B(n_6400),
.Y(n_19795)
);

AOI22xp33_ASAP7_75t_L g19796 ( 
.A1(n_19792),
.A2(n_7371),
.B1(n_7431),
.B2(n_7350),
.Y(n_19796)
);

AOI21xp5_ASAP7_75t_L g19797 ( 
.A1(n_19789),
.A2(n_6854),
.B(n_6807),
.Y(n_19797)
);

XNOR2x1_ASAP7_75t_L g19798 ( 
.A(n_19791),
.B(n_6419),
.Y(n_19798)
);

AOI32xp33_ASAP7_75t_L g19799 ( 
.A1(n_19798),
.A2(n_19793),
.A3(n_6597),
.B1(n_6459),
.B2(n_6528),
.Y(n_19799)
);

BUFx3_ASAP7_75t_L g19800 ( 
.A(n_19794),
.Y(n_19800)
);

AOI22xp33_ASAP7_75t_L g19801 ( 
.A1(n_19795),
.A2(n_7371),
.B1(n_7431),
.B2(n_7350),
.Y(n_19801)
);

XOR2xp5_ASAP7_75t_L g19802 ( 
.A(n_19800),
.B(n_19797),
.Y(n_19802)
);

OR2x2_ASAP7_75t_L g19803 ( 
.A(n_19801),
.B(n_19795),
.Y(n_19803)
);

INVx1_ASAP7_75t_L g19804 ( 
.A(n_19799),
.Y(n_19804)
);

OAI22xp5_ASAP7_75t_L g19805 ( 
.A1(n_19802),
.A2(n_19796),
.B1(n_6456),
.B2(n_6459),
.Y(n_19805)
);

AOI22xp5_ASAP7_75t_L g19806 ( 
.A1(n_19804),
.A2(n_4748),
.B1(n_4608),
.B2(n_4544),
.Y(n_19806)
);

OAI21xp5_ASAP7_75t_L g19807 ( 
.A1(n_19803),
.A2(n_7987),
.B(n_7931),
.Y(n_19807)
);

OAI221xp5_ASAP7_75t_R g19808 ( 
.A1(n_19805),
.A2(n_6854),
.B1(n_7483),
.B2(n_7722),
.C(n_4748),
.Y(n_19808)
);

AOI22xp5_ASAP7_75t_L g19809 ( 
.A1(n_19808),
.A2(n_19806),
.B1(n_19807),
.B2(n_4748),
.Y(n_19809)
);

AOI211xp5_ASAP7_75t_L g19810 ( 
.A1(n_19809),
.A2(n_6435),
.B(n_6459),
.C(n_6456),
.Y(n_19810)
);


endmodule