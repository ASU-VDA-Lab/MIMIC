module fake_jpeg_18752_n_86 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_14),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_15),
.B1(n_19),
.B2(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_32),
.B1(n_11),
.B2(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_27),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_23),
.B1(n_20),
.B2(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_14),
.C(n_35),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_49),
.B1(n_8),
.B2(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_53),
.B(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_69),
.C(n_64),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_59),
.B1(n_55),
.B2(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_72),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_12),
.Y(n_77)
);

OA21x2_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_58),
.B(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_75),
.B(n_76),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_58),
.C(n_10),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_77),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_4),
.B(n_5),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_78),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_81),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_6),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_6),
.Y(n_86)
);


endmodule