module real_jpeg_6720_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_2),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_2),
.B(n_67),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_2),
.B(n_105),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_2),
.B(n_51),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_2),
.B(n_250),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_2),
.B(n_269),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_2),
.B(n_402),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_3),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_3),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_60),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_4),
.B(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_5),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_5),
.Y(n_310)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_7),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_7),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_7),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_7),
.B(n_400),
.Y(n_399)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_9),
.B(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_9),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_10),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_10),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_10),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_10),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_10),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_13),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_13),
.B(n_165),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_13),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_13),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_13),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_14),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_14),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_14),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_80),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_15),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_15),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_15),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_15),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_15),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_15),
.B(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_16),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_17),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_17),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_17),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_17),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_17),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_17),
.B(n_250),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_195),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_194),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_143),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_21),
.B(n_143),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_21),
.Y(n_442)
);

FAx1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_90),
.CI(n_118),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_61),
.C(n_74),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_23),
.A2(n_24),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.C(n_48),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_25),
.A2(n_26),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_32),
.C(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_42),
.C(n_45),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_32),
.A2(n_33),
.B1(n_45),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_35),
.B(n_93),
.C(n_96),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_35),
.A2(n_36),
.B1(n_96),
.B2(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_40),
.Y(n_307)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_40),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_41),
.B(n_48),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_42),
.A2(n_43),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_45),
.Y(n_171)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_47),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_47),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_50),
.B(n_55),
.C(n_59),
.Y(n_140)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_54),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_74),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_68),
.C(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_68),
.A2(n_69),
.B1(n_88),
.B2(n_89),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_75),
.C(n_88),
.Y(n_74)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_72),
.Y(n_226)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_76),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_84),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_77),
.B(n_81),
.CI(n_84),
.CON(n_152),
.SN(n_152)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_80),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_86),
.Y(n_246)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_110),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_97),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_108),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_100),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_103),
.B1(n_108),
.B2(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_107),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_114),
.Y(n_319)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_137),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_135),
.B2(n_136),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_144),
.B(n_147),
.Y(n_438)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_149),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_172),
.C(n_174),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_150),
.A2(n_151),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_168),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_152),
.B(n_420),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g443 ( 
.A(n_152),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_153),
.B(n_168),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_164),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_154),
.B(n_164),
.Y(n_396)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_158),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_172),
.B(n_174),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.C(n_191),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_175),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_184),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_176),
.B(n_387),
.Y(n_386)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_178),
.A2(n_179),
.B1(n_184),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_183),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_184),
.Y(n_388)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_187),
.B(n_191),
.Y(n_417)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_190),
.Y(n_316)
);

INVx6_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_436),
.B(n_440),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_424),
.B(n_435),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_406),
.B(n_423),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_380),
.B(n_405),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_300),
.B(n_379),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_285),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_201),
.B(n_285),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_240),
.B2(n_284),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_202),
.B(n_241),
.C(n_270),
.Y(n_404)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_218),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_204),
.B(n_219),
.C(n_239),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.C(n_217),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_205),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_215),
.B(n_217),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_228),
.B1(n_238),
.B2(n_239),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_223),
.B(n_227),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_223),
.Y(n_227)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_227),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_227),
.B(n_385),
.C(n_390),
.Y(n_413)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_403)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_270),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_253),
.C(n_264),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_247),
.C(n_252),
.Y(n_283)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_251),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_254),
.B1(n_264),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_262),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_255),
.A2(n_256),
.B1(n_262),
.B2(n_263),
.Y(n_372)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_258),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_259),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

XOR2x1_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_281),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_271),
.B(n_282),
.C(n_283),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_272),
.B(n_276),
.C(n_279),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_276),
.Y(n_280)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_298),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_286),
.B(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_289),
.B(n_298),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_290),
.B(n_291),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_292),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_296),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_374),
.B(n_378),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_359),
.B(n_373),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_339),
.B(n_358),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_326),
.B(n_338),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_308),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_320),
.B2(n_321),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_317),
.C(n_320),
.Y(n_357)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_325),
.Y(n_343)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_333),
.B(n_337),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_329),
.Y(n_337)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_357),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_357),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_343),
.C(n_361),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_354),
.C(n_356),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx11_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_349)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_362),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_366),
.B2(n_367),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_369),
.C(n_370),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_376),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_404),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_404),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_392),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_384),
.C(n_392),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_389),
.B2(n_391),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_389),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_395),
.C(n_397),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_403),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_401),
.C(n_403),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_408),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_419),
.C(n_421),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_419),
.B1(n_421),
.B2(n_422),
.Y(n_410)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_411),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_414),
.B2(n_418),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_415),
.C(n_416),
.Y(n_426)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_414),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_419),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_434),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_434),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_428),
.C(n_431),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_429),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_432),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_439),
.Y(n_440)
);


endmodule