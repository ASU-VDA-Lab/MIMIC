module fake_jpeg_30275_n_469 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_47),
.Y(n_143)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_50),
.B(n_56),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_53),
.Y(n_133)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_7),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_63),
.Y(n_106)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_73),
.Y(n_113)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_9),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_25),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_15),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_88),
.Y(n_136)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_17),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_33),
.Y(n_114)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_17),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_25),
.B1(n_93),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_124),
.B1(n_125),
.B2(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_46),
.B1(n_45),
.B2(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_102),
.A2(n_141),
.B1(n_70),
.B2(n_82),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_38),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_144),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_46),
.B1(n_27),
.B2(n_17),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_84),
.B1(n_53),
.B2(n_17),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_126),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_49),
.A2(n_45),
.B1(n_42),
.B2(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_54),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_59),
.A2(n_20),
.B1(n_35),
.B2(n_38),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_88),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_60),
.A2(n_85),
.B1(n_90),
.B2(n_89),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_77),
.A2(n_88),
.B1(n_83),
.B2(n_47),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_77),
.B1(n_53),
.B2(n_111),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_32),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_143),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_66),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_62),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_153),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_163),
.Y(n_197)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_147),
.B1(n_98),
.B2(n_127),
.Y(n_208)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_27),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_162),
.A2(n_40),
.A3(n_44),
.B1(n_41),
.B2(n_30),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_97),
.A2(n_27),
.B(n_23),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_167),
.A2(n_27),
.B(n_64),
.C(n_81),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_174),
.Y(n_205)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_173),
.A2(n_175),
.B1(n_181),
.B2(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_113),
.B(n_40),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_74),
.C(n_87),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_184),
.C(n_187),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_124),
.B1(n_134),
.B2(n_125),
.Y(n_194)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_121),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_183),
.Y(n_198)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_32),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_57),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_41),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_100),
.B(n_91),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_111),
.A2(n_48),
.B1(n_34),
.B2(n_26),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_120),
.Y(n_210)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_26),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_193),
.Y(n_213)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_34),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_208),
.B1(n_209),
.B2(n_215),
.Y(n_244)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_116),
.A3(n_140),
.B1(n_146),
.B2(n_110),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_231),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_135),
.B1(n_147),
.B2(n_127),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_219),
.B(n_149),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_140),
.C(n_100),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_228),
.C(n_187),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_142),
.B1(n_69),
.B2(n_80),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_167),
.A2(n_68),
.B1(n_71),
.B2(n_98),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_223),
.B1(n_224),
.B2(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_164),
.B(n_44),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_154),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_163),
.A2(n_119),
.B1(n_137),
.B2(n_131),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_153),
.A2(n_151),
.B1(n_184),
.B2(n_161),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_146),
.C(n_95),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_186),
.A2(n_137),
.B1(n_99),
.B2(n_23),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_190),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_157),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_238),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_182),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_148),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_200),
.C(n_229),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_184),
.B1(n_153),
.B2(n_151),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_241),
.A2(n_243),
.B1(n_265),
.B2(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_246),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_162),
.B1(n_178),
.B2(n_170),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_202),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_187),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_150),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_251),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_220),
.B(n_219),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_171),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_149),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_196),
.B(n_203),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_264),
.B(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_95),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_220),
.B(n_200),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_172),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_199),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_192),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_257),
.B(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_189),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_222),
.B(n_168),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_194),
.B(n_160),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_219),
.A2(n_181),
.B(n_152),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_196),
.A2(n_175),
.B1(n_159),
.B2(n_154),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_271),
.C(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_280),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_231),
.B(n_210),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_272),
.A2(n_286),
.B(n_234),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_276),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_201),
.C(n_205),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_232),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_205),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_284),
.C(n_245),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_208),
.B1(n_217),
.B2(n_215),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_244),
.B1(n_258),
.B2(n_243),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_204),
.C(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_292),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_294),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_291),
.A2(n_251),
.B1(n_255),
.B2(n_260),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_199),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_265),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_285),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_305),
.A2(n_309),
.B1(n_313),
.B2(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_308),
.B(n_280),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_244),
.B1(n_249),
.B2(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_311),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_279),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_249),
.B1(n_264),
.B2(n_234),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_314),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_320),
.B1(n_322),
.B2(n_324),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_325),
.B(n_273),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_255),
.C(n_251),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_327),
.C(n_328),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_277),
.A2(n_243),
.B1(n_241),
.B2(n_239),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_255),
.B1(n_253),
.B2(n_245),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_284),
.A2(n_278),
.B1(n_287),
.B2(n_297),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_286),
.A2(n_246),
.B(n_242),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_323),
.A2(n_227),
.B(n_206),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_295),
.A2(n_238),
.B1(n_236),
.B2(n_235),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_253),
.B(n_240),
.Y(n_325)
);

BUFx24_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_326),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_239),
.C(n_248),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_281),
.C(n_278),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_339),
.C(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_293),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_347),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_344),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_273),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_336),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_297),
.C(n_271),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_267),
.B1(n_283),
.B2(n_270),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_343),
.B1(n_355),
.B2(n_326),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_270),
.B1(n_272),
.B2(n_241),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_304),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_293),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_356),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_275),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_298),
.B(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_275),
.C(n_274),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_274),
.C(n_247),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_323),
.C(n_311),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_328),
.B(n_261),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_319),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_321),
.A2(n_259),
.B1(n_254),
.B2(n_233),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_300),
.Y(n_360)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_331),
.B(n_325),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_366),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_298),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_305),
.B1(n_309),
.B2(n_322),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_370),
.B1(n_377),
.B2(n_355),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_348),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_372),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_317),
.B1(n_313),
.B2(n_326),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_303),
.Y(n_371)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_306),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_347),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_374),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_339),
.C(n_329),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_307),
.B1(n_299),
.B2(n_207),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_335),
.A2(n_211),
.B1(n_204),
.B2(n_230),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_335),
.A2(n_211),
.B1(n_225),
.B2(n_230),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_212),
.B1(n_31),
.B2(n_3),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_385),
.C(n_389),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_332),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_397),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_388),
.A2(n_378),
.B1(n_381),
.B2(n_370),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_332),
.C(n_346),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_352),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_395),
.C(n_399),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_354),
.B(n_341),
.Y(n_393)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_393),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_375),
.C(n_374),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_396),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_356),
.Y(n_397)
);

NOR3xp33_ASAP7_75t_SL g398 ( 
.A(n_366),
.B(n_337),
.C(n_342),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_SL g416 ( 
.A(n_398),
.B(n_372),
.C(n_377),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_350),
.C(n_31),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_31),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_395),
.C(n_399),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_358),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_409),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_385),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_383),
.A2(n_362),
.B(n_371),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_412),
.A2(n_416),
.B(n_392),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_364),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_414),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_391),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_418),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_363),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_431),
.Y(n_438)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_388),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_425),
.C(n_427),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_402),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_367),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_389),
.C(n_392),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_0),
.C(n_1),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_398),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_363),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_433),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_9),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_405),
.A2(n_11),
.B(n_14),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_434),
.B(n_5),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_422),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_440),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_429),
.A2(n_414),
.B1(n_419),
.B2(n_417),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_439),
.A2(n_443),
.B1(n_446),
.B2(n_437),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_421),
.A2(n_416),
.B1(n_405),
.B2(n_58),
.Y(n_440)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_444),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_5),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_426),
.A2(n_11),
.B(n_13),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_446),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_0),
.C(n_1),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_424),
.Y(n_448)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_448),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_449),
.A2(n_451),
.B(n_3),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_430),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_435),
.A2(n_421),
.B1(n_425),
.B2(n_420),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_454),
.B1(n_4),
.B2(n_12),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_459),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_449),
.A2(n_4),
.B(n_11),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_461),
.B(n_455),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_453),
.A2(n_4),
.B(n_12),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_4),
.C(n_12),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_450),
.B(n_452),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_464),
.B1(n_12),
.B2(n_13),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_462),
.A2(n_457),
.B(n_448),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_466),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_13),
.C(n_14),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_13),
.Y(n_469)
);


endmodule