module fake_jpeg_30972_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_0),
.B(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_18),
.C(n_17),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_31),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_29),
.B(n_26),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.C(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_38),
.B(n_36),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_35),
.B(n_25),
.Y(n_41)
);


endmodule