module fake_jpeg_17601_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_9),
.B(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_27),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_10),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_10),
.B(n_1),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_18),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_17),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_13),
.C(n_19),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_27),
.B1(n_15),
.B2(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_52),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_51),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_24),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_26),
.B(n_11),
.C(n_17),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_33),
.C(n_30),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_71),
.C(n_49),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_47),
.B(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_68),
.B1(n_36),
.B2(n_40),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_40),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_53),
.B(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_33),
.C(n_31),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_52),
.C(n_20),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_23),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_71),
.C(n_67),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_18),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_21),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_87),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_73),
.C(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_94),
.C(n_95),
.Y(n_101)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_96),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_23),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_13),
.C(n_36),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_83),
.B1(n_82),
.B2(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_101),
.B1(n_96),
.B2(n_3),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_92),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.C(n_105),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_96),
.B1(n_91),
.B2(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_106),
.Y(n_111)
);


endmodule