module fake_jpeg_30038_n_46 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_21),
.B(n_1),
.C(n_2),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_0),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_5),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_35),
.B(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_36),
.C(n_32),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_28),
.C(n_9),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_5),
.B(n_6),
.Y(n_43)
);

NOR2xp67_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_6),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_7),
.B(n_8),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_42),
.Y(n_46)
);


endmodule