module fake_jpeg_27170_n_262 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_13),
.B1(n_20),
.B2(n_19),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_58),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_59),
.B1(n_33),
.B2(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_28),
.B1(n_33),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_44),
.B1(n_33),
.B2(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_77),
.B1(n_39),
.B2(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_72),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_62),
.B1(n_59),
.B2(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_41),
.B1(n_24),
.B2(n_25),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_82),
.Y(n_83)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_49),
.B1(n_47),
.B2(n_51),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_93),
.B1(n_95),
.B2(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_87),
.B1(n_98),
.B2(n_40),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_72),
.B1(n_80),
.B2(n_75),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_49),
.A3(n_58),
.B1(n_30),
.B2(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_59),
.C(n_26),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_97),
.C(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_42),
.B1(n_37),
.B2(n_53),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_70),
.C(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_53),
.B1(n_42),
.B2(n_56),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_18),
.B(n_63),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_107),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_119),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_76),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_18),
.B(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_71),
.B(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_56),
.B1(n_71),
.B2(n_48),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_35),
.B1(n_40),
.B2(n_21),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_91),
.B1(n_96),
.B2(n_99),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_35),
.B1(n_21),
.B2(n_34),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_31),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_118),
.B1(n_102),
.B2(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_129),
.C(n_22),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_99),
.C(n_96),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_135),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_101),
.B1(n_116),
.B2(n_115),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_26),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_138),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_34),
.B(n_26),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_112),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_17),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_15),
.B1(n_23),
.B2(n_16),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_12),
.B1(n_23),
.B2(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_15),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_150),
.B(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_148),
.B1(n_142),
.B2(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_15),
.B1(n_23),
.B2(n_16),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_0),
.B(n_3),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_137),
.B(n_121),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_26),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_12),
.B1(n_23),
.B2(n_16),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_132),
.B1(n_131),
.B2(n_127),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_0),
.B(n_3),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

OAI22x1_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_128),
.B1(n_135),
.B2(n_136),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_14),
.B1(n_12),
.B2(n_22),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_178),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_142),
.B1(n_134),
.B2(n_34),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_14),
.B1(n_12),
.B2(n_15),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_29),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_29),
.C(n_22),
.D(n_14),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_159),
.A3(n_145),
.B1(n_157),
.B2(n_147),
.C1(n_165),
.C2(n_152),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_166),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_161),
.C(n_158),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_183),
.C(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_144),
.B1(n_154),
.B2(n_156),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_186),
.B1(n_167),
.B2(n_190),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_169),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_22),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_175),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_176),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_174),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_22),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_194),
.C(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_185),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_197),
.B1(n_196),
.B2(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_199),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_222),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_207),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_29),
.C(n_5),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_204),
.B(n_5),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_238),
.B(n_10),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_29),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_4),
.C(n_7),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_225),
.B1(n_223),
.B2(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_225),
.B(n_5),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_4),
.B(n_7),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_7),
.C(n_8),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_248),
.B(n_250),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_8),
.C(n_9),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_9),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_258),
.B(n_256),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_259),
.B(n_9),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_10),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_10),
.Y(n_262)
);


endmodule