module real_aes_17538_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1914;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_1899;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_1343;
wire n_465;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1931;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1633 ( .A1(n_0), .A2(n_113), .B1(n_1625), .B2(n_1628), .Y(n_1633) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1), .Y(n_1124) );
INVx1_ASAP7_75t_L g897 ( .A(n_2), .Y(n_897) );
AO22x1_ASAP7_75t_L g922 ( .A1(n_2), .A2(n_248), .B1(n_525), .B2(n_608), .Y(n_922) );
INVx1_ASAP7_75t_L g388 ( .A(n_3), .Y(n_388) );
AND2x2_ASAP7_75t_L g459 ( .A(n_3), .B(n_271), .Y(n_459) );
AND2x2_ASAP7_75t_L g476 ( .A(n_3), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_3), .B(n_398), .Y(n_695) );
INVx1_ASAP7_75t_L g906 ( .A(n_4), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_4), .A2(n_146), .B1(n_478), .B2(n_492), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g1210 ( .A1(n_5), .A2(n_338), .B1(n_466), .B2(n_1167), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_5), .A2(n_6), .B1(n_497), .B2(n_1225), .C(n_1227), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1215 ( .A1(n_6), .A2(n_9), .B1(n_641), .B2(n_1025), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g1166 ( .A1(n_7), .A2(n_335), .B1(n_1013), .B2(n_1167), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_7), .A2(n_281), .B1(n_832), .B2(n_1140), .C(n_1184), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_8), .A2(n_218), .B1(n_646), .B2(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_8), .A2(n_203), .B1(n_610), .B2(n_1043), .Y(n_1142) );
A2O1A1Ixp33_ASAP7_75t_L g1238 ( .A1(n_9), .A2(n_1061), .B(n_1239), .C(n_1245), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1934 ( .A1(n_10), .A2(n_238), .B1(n_437), .B2(n_1288), .Y(n_1934) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_11), .A2(n_241), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_11), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_12), .A2(n_330), .B1(n_517), .B2(n_797), .C(n_1353), .Y(n_1352) );
AOI22xp33_ASAP7_75t_SL g1369 ( .A1(n_12), .A2(n_351), .B1(n_582), .B2(n_732), .Y(n_1369) );
INVxp67_ASAP7_75t_SL g587 ( .A(n_13), .Y(n_587) );
AND4x1_ASAP7_75t_L g657 ( .A(n_13), .B(n_589), .C(n_594), .D(n_627), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_14), .A2(n_311), .B1(n_578), .B2(n_1264), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_14), .A2(n_103), .B1(n_492), .B2(n_516), .C(n_606), .Y(n_1268) );
INVx2_ASAP7_75t_L g419 ( .A(n_15), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g1317 ( .A1(n_16), .A2(n_305), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
OAI221xp5_ASAP7_75t_L g1329 ( .A1(n_16), .A2(n_305), .B1(n_474), .B2(n_506), .C(n_1330), .Y(n_1329) );
XNOR2x1_ASAP7_75t_L g1297 ( .A(n_17), .B(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1918 ( .A(n_18), .Y(n_1918) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_19), .A2(n_246), .B1(n_732), .B2(n_1261), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_19), .A2(n_161), .B1(n_1270), .B2(n_1272), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_20), .A2(n_328), .B1(n_1187), .B2(n_1231), .Y(n_1527) );
INVx1_ASAP7_75t_L g1549 ( .A(n_20), .Y(n_1549) );
INVx1_ASAP7_75t_L g992 ( .A(n_21), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_22), .A2(n_285), .B1(n_1046), .B2(n_1186), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_22), .A2(n_282), .B1(n_724), .B2(n_859), .Y(n_1373) );
INVx1_ASAP7_75t_L g1916 ( .A(n_23), .Y(n_1916) );
AOI22xp33_ASAP7_75t_L g1928 ( .A1(n_23), .A2(n_83), .B1(n_1044), .B2(n_1105), .Y(n_1928) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_24), .A2(n_185), .B1(n_533), .B2(n_593), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_24), .A2(n_523), .B(n_596), .C(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g1531 ( .A(n_25), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_26), .A2(n_149), .B1(n_646), .B2(n_1080), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_26), .A2(n_313), .B1(n_1044), .B2(n_1105), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_27), .A2(n_110), .B1(n_608), .B2(n_610), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_27), .A2(n_38), .B1(n_644), .B2(n_646), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_28), .Y(n_1291) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_29), .Y(n_383) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_29), .B(n_381), .Y(n_1619) );
INVx1_ASAP7_75t_L g1328 ( .A(n_30), .Y(n_1328) );
OAI211xp5_ASAP7_75t_SL g1580 ( .A1(n_31), .A2(n_523), .B(n_1581), .C(n_1585), .Y(n_1580) );
OAI22xp5_ASAP7_75t_L g1590 ( .A1(n_31), .A2(n_293), .B1(n_437), .B2(n_1303), .Y(n_1590) );
OAI22xp5_ASAP7_75t_SL g959 ( .A1(n_32), .A2(n_314), .B1(n_960), .B2(n_961), .Y(n_959) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_32), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_33), .Y(n_1000) );
INVx1_ASAP7_75t_L g422 ( .A(n_34), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_34), .A2(n_472), .B(n_480), .C(n_499), .Y(n_471) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_35), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_36), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_37), .A2(n_351), .B1(n_828), .B2(n_1186), .Y(n_1358) );
AOI22xp5_ASAP7_75t_L g1370 ( .A1(n_37), .A2(n_330), .B1(n_732), .B2(n_1371), .Y(n_1370) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_38), .A2(n_360), .B1(n_492), .B2(n_625), .C(n_626), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g1438 ( .A(n_39), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_40), .A2(n_60), .B1(n_647), .B2(n_651), .Y(n_792) );
INVx1_ASAP7_75t_L g805 ( .A(n_40), .Y(n_805) );
AOI21xp33_ASAP7_75t_L g1390 ( .A1(n_41), .A2(n_517), .B(n_1041), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_41), .A2(n_341), .B1(n_732), .B2(n_870), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_42), .A2(n_82), .B1(n_1618), .B2(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g705 ( .A(n_43), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_44), .A2(n_59), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_44), .A2(n_183), .B1(n_650), .B2(n_732), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_45), .A2(n_132), .B1(n_606), .B2(n_625), .C(n_1395), .Y(n_1523) );
INVx1_ASAP7_75t_L g1550 ( .A(n_45), .Y(n_1550) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_46), .A2(n_115), .B1(n_1130), .B2(n_1132), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_46), .A2(n_220), .B1(n_1184), .B2(n_1241), .C(n_1242), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1568 ( .A(n_47), .B(n_449), .Y(n_1568) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_48), .A2(n_331), .B1(n_492), .B2(n_516), .C(n_517), .Y(n_515) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_48), .Y(n_545) );
INVx1_ASAP7_75t_L g1403 ( .A(n_49), .Y(n_1403) );
INVx1_ASAP7_75t_L g1844 ( .A(n_50), .Y(n_1844) );
INVx1_ASAP7_75t_L g464 ( .A(n_51), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_51), .A2(n_232), .B1(n_520), .B2(n_523), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_52), .A2(n_369), .B1(n_433), .B2(n_783), .C(n_784), .Y(n_782) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_52), .A2(n_138), .B1(n_796), .B2(n_797), .C(n_804), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_53), .Y(n_1428) );
OAI211xp5_ASAP7_75t_SL g1453 ( .A1(n_54), .A2(n_1280), .B(n_1454), .C(n_1457), .Y(n_1453) );
INVx1_ASAP7_75t_L g1503 ( .A(n_54), .Y(n_1503) );
CKINVDCx5p33_ASAP7_75t_R g1434 ( .A(n_55), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_56), .A2(n_304), .B1(n_855), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1050 ( .A(n_56), .Y(n_1050) );
OAI21xp5_ASAP7_75t_L g1362 ( .A1(n_57), .A2(n_1303), .B(n_1363), .Y(n_1362) );
NAND5xp2_ASAP7_75t_L g820 ( .A(n_58), .B(n_821), .C(n_850), .D(n_866), .E(n_873), .Y(n_820) );
INVx1_ASAP7_75t_L g882 ( .A(n_58), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_59), .A2(n_197), .B1(n_719), .B2(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g799 ( .A(n_60), .Y(n_799) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_61), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_61), .A2(n_157), .B1(n_577), .B2(n_578), .Y(n_576) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_62), .Y(n_395) );
INVx1_ASAP7_75t_L g597 ( .A(n_63), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_63), .A2(n_119), .B1(n_630), .B2(n_635), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g1127 ( .A1(n_64), .A2(n_65), .B1(n_724), .B2(n_1023), .Y(n_1127) );
INVx1_ASAP7_75t_L g1146 ( .A(n_64), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g1139 ( .A1(n_65), .A2(n_158), .B1(n_601), .B2(n_606), .C(n_1140), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1644 ( .A1(n_66), .A2(n_133), .B1(n_1618), .B2(n_1632), .Y(n_1644) );
INVx1_ASAP7_75t_L g1400 ( .A(n_67), .Y(n_1400) );
OAI22xp33_ASAP7_75t_L g1414 ( .A1(n_67), .A2(n_332), .B1(n_868), .B2(n_1086), .Y(n_1414) );
AOI22xp5_ASAP7_75t_L g1651 ( .A1(n_68), .A2(n_275), .B1(n_1618), .B2(n_1632), .Y(n_1651) );
INVx1_ASAP7_75t_L g1008 ( .A(n_69), .Y(n_1008) );
INVx1_ASAP7_75t_L g1254 ( .A(n_70), .Y(n_1254) );
OAI222xp33_ASAP7_75t_L g1278 ( .A1(n_70), .A2(n_373), .B1(n_614), .B2(n_1093), .C1(n_1279), .C2(n_1284), .Y(n_1278) );
INVx1_ASAP7_75t_L g1327 ( .A(n_71), .Y(n_1327) );
INVx1_ASAP7_75t_L g1462 ( .A(n_72), .Y(n_1462) );
OAI211xp5_ASAP7_75t_L g1490 ( .A1(n_72), .A2(n_1491), .B(n_1493), .C(n_1495), .Y(n_1490) );
XOR2x2_ASAP7_75t_L g1415 ( .A(n_73), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1536 ( .A(n_74), .Y(n_1536) );
OAI332xp33_ASAP7_75t_SL g1539 ( .A1(n_74), .A2(n_630), .A3(n_861), .B1(n_1540), .B2(n_1546), .B3(n_1547), .C1(n_1553), .C2(n_1557), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g1277 ( .A(n_75), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1582 ( .A1(n_76), .A2(n_134), .B1(n_497), .B2(n_1226), .C(n_1583), .Y(n_1582) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_76), .A2(n_267), .B1(n_1025), .B2(n_1135), .Y(n_1598) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_77), .A2(n_194), .B1(n_478), .B2(n_492), .C(n_517), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_77), .A2(n_255), .B1(n_732), .B2(n_857), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_78), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_79), .A2(n_255), .B1(n_608), .B2(n_828), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_79), .A2(n_194), .B1(n_732), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_80), .A2(n_179), .B1(n_1019), .B2(n_1129), .Y(n_1170) );
AOI21xp33_ASAP7_75t_L g1193 ( .A1(n_80), .A2(n_601), .B(n_626), .Y(n_1193) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_81), .A2(n_359), .B1(n_601), .B2(n_603), .C(n_606), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_81), .A2(n_320), .B1(n_650), .B2(n_652), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1342 ( .A1(n_82), .A2(n_1343), .B1(n_1344), .B2(n_1375), .Y(n_1342) );
INVxp67_ASAP7_75t_SL g1375 ( .A(n_82), .Y(n_1375) );
INVx1_ASAP7_75t_L g1906 ( .A(n_83), .Y(n_1906) );
OAI22xp33_ASAP7_75t_L g1876 ( .A1(n_84), .A2(n_324), .B1(n_390), .B2(n_1877), .Y(n_1876) );
OAI22xp33_ASAP7_75t_L g1879 ( .A1(n_84), .A2(n_324), .B1(n_1484), .B2(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1207 ( .A(n_85), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_86), .A2(n_274), .B1(n_1187), .B2(n_1231), .Y(n_1524) );
INVx1_ASAP7_75t_L g1556 ( .A(n_86), .Y(n_1556) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_87), .A2(n_356), .B1(n_671), .B2(n_674), .C(n_678), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_87), .A2(n_316), .B1(n_727), .B2(n_728), .C(n_730), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_88), .A2(n_116), .B1(n_1046), .B2(n_1105), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_88), .A2(n_252), .B1(n_1022), .B2(n_1025), .Y(n_1413) );
AOI22xp33_ASAP7_75t_SL g1012 ( .A1(n_89), .A2(n_200), .B1(n_727), .B2(n_1013), .Y(n_1012) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_89), .Y(n_1056) );
OAI211xp5_ASAP7_75t_SL g773 ( .A1(n_90), .A2(n_741), .B(n_748), .C(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g810 ( .A(n_90), .Y(n_810) );
INVx1_ASAP7_75t_L g1533 ( .A(n_91), .Y(n_1533) );
INVx1_ASAP7_75t_L g1350 ( .A(n_92), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1173 ( .A(n_93), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_94), .Y(n_841) );
OAI21xp5_ASAP7_75t_SL g1198 ( .A1(n_95), .A2(n_533), .B(n_1199), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_96), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_96), .A2(n_366), .B1(n_734), .B2(n_737), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_97), .A2(n_264), .B1(n_1618), .B2(n_1632), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g1431 ( .A(n_98), .Y(n_1431) );
AOI22xp33_ASAP7_75t_SL g1169 ( .A1(n_99), .A2(n_281), .B1(n_641), .B2(n_1023), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_99), .A2(n_335), .B1(n_610), .B2(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1351 ( .A(n_100), .Y(n_1351) );
OR2x2_ASAP7_75t_L g448 ( .A(n_101), .B(n_449), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_102), .A2(n_230), .B1(n_502), .B2(n_506), .C(n_511), .Y(n_501) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_102), .A2(n_544), .A3(n_552), .B1(n_555), .B2(n_563), .C1(n_569), .C2(n_580), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_103), .A2(n_152), .B1(n_578), .B2(n_1261), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1637 ( .A1(n_104), .A2(n_270), .B1(n_1625), .B2(n_1628), .Y(n_1637) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_105), .A2(n_182), .B1(n_525), .B2(n_965), .Y(n_964) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_105), .Y(n_988) );
INVx1_ASAP7_75t_L g1301 ( .A(n_106), .Y(n_1301) );
AOI22xp33_ASAP7_75t_SL g1310 ( .A1(n_107), .A2(n_308), .B1(n_853), .B2(n_990), .Y(n_1310) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_107), .A2(n_114), .B1(n_496), .B2(n_832), .C(n_1041), .Y(n_1323) );
INVx1_ASAP7_75t_L g1064 ( .A(n_108), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1638 ( .A1(n_108), .A2(n_124), .B1(n_1618), .B2(n_1639), .Y(n_1638) );
AO22x1_ASAP7_75t_L g1624 ( .A1(n_109), .A2(n_277), .B1(n_1625), .B2(n_1628), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_110), .A2(n_360), .B1(n_644), .B2(n_646), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g1287 ( .A1(n_111), .A2(n_1288), .B(n_1289), .Y(n_1287) );
INVx1_ASAP7_75t_L g1304 ( .A(n_112), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_114), .A2(n_212), .B1(n_577), .B2(n_727), .Y(n_1316) );
AOI22xp33_ASAP7_75t_SL g1230 ( .A1(n_115), .A2(n_155), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_116), .A2(n_279), .B1(n_432), .B2(n_1013), .Y(n_1410) );
INVx1_ASAP7_75t_L g1915 ( .A(n_117), .Y(n_1915) );
AOI221xp5_ASAP7_75t_L g1923 ( .A1(n_117), .A2(n_243), .B1(n_516), .B2(n_626), .C(n_1140), .Y(n_1923) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_118), .Y(n_1181) );
INVx1_ASAP7_75t_L g598 ( .A(n_119), .Y(n_598) );
OAI211xp5_ASAP7_75t_L g834 ( .A1(n_120), .A2(n_835), .B(n_837), .C(n_839), .Y(n_834) );
INVx1_ASAP7_75t_L g878 ( .A(n_120), .Y(n_878) );
INVx1_ASAP7_75t_L g1122 ( .A(n_121), .Y(n_1122) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_121), .A2(n_160), .B1(n_506), .B2(n_613), .C(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g512 ( .A(n_122), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_123), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_123), .A2(n_142), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_125), .A2(n_251), .B1(n_525), .B2(n_827), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_125), .A2(n_276), .B1(n_641), .B2(n_723), .Y(n_984) );
INVx1_ASAP7_75t_L g1574 ( .A(n_126), .Y(n_1574) );
INVx1_ASAP7_75t_L g950 ( .A(n_127), .Y(n_950) );
INVx1_ASAP7_75t_L g1125 ( .A(n_128), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_129), .A2(n_291), .B1(n_613), .B2(n_614), .C(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g656 ( .A(n_129), .Y(n_656) );
INVx1_ASAP7_75t_L g381 ( .A(n_130), .Y(n_381) );
INVx1_ASAP7_75t_L g1849 ( .A(n_131), .Y(n_1849) );
INVx1_ASAP7_75t_L g1562 ( .A(n_132), .Y(n_1562) );
AOI22xp33_ASAP7_75t_L g1596 ( .A1(n_134), .A2(n_284), .B1(n_432), .B2(n_1135), .Y(n_1596) );
INVx1_ASAP7_75t_L g1586 ( .A(n_135), .Y(n_1586) );
OAI22xp33_ASAP7_75t_L g1600 ( .A1(n_135), .A2(n_206), .B1(n_630), .B2(n_868), .Y(n_1600) );
AO221x2_ASAP7_75t_L g1703 ( .A1(n_136), .A2(n_358), .B1(n_1625), .B2(n_1628), .C(n_1704), .Y(n_1703) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_137), .A2(n_207), .B1(n_855), .B2(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1054 ( .A(n_137), .Y(n_1054) );
INVx1_ASAP7_75t_L g789 ( .A(n_138), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g1903 ( .A1(n_139), .A2(n_325), .B1(n_630), .B2(n_635), .Y(n_1903) );
INVx1_ASAP7_75t_L g1930 ( .A(n_139), .Y(n_1930) );
OAI222xp33_ASAP7_75t_L g912 ( .A1(n_140), .A2(n_355), .B1(n_744), .B2(n_746), .C1(n_913), .C2(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g925 ( .A(n_140), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g1427 ( .A(n_141), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_142), .Y(n_1175) );
INVx1_ASAP7_75t_L g1387 ( .A(n_143), .Y(n_1387) );
OAI211xp5_ASAP7_75t_L g1392 ( .A1(n_144), .A2(n_1102), .B(n_1393), .C(n_1399), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_144), .A2(n_286), .B1(n_437), .B2(n_1303), .Y(n_1404) );
INVx1_ASAP7_75t_L g1835 ( .A(n_145), .Y(n_1835) );
INVx1_ASAP7_75t_L g902 ( .A(n_146), .Y(n_902) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_147), .A2(n_954), .B(n_955), .C(n_956), .Y(n_953) );
INVxp33_ASAP7_75t_SL g976 ( .A(n_147), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_148), .A2(n_192), .B1(n_752), .B2(n_755), .Y(n_751) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_148), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_149), .A2(n_258), .B1(n_516), .B2(n_626), .C(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1907 ( .A(n_150), .Y(n_1907) );
AOI221xp5_ASAP7_75t_L g1926 ( .A1(n_150), .A2(n_302), .B1(n_516), .B2(n_1241), .C(n_1927), .Y(n_1926) );
INVx1_ASAP7_75t_L g1356 ( .A(n_151), .Y(n_1356) );
INVx1_ASAP7_75t_L g1282 ( .A(n_152), .Y(n_1282) );
INVxp67_ASAP7_75t_SL g1389 ( .A(n_153), .Y(n_1389) );
AOI22xp33_ASAP7_75t_SL g1412 ( .A1(n_153), .A2(n_298), .B1(n_582), .B2(n_732), .Y(n_1412) );
INVx1_ASAP7_75t_L g1004 ( .A(n_154), .Y(n_1004) );
OAI222xp33_ASAP7_75t_L g1048 ( .A1(n_154), .A2(n_228), .B1(n_472), .B2(n_614), .C1(n_1049), .C2(n_1055), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_155), .A2(n_220), .B1(n_1130), .B2(n_1213), .Y(n_1212) );
XOR2x2_ASAP7_75t_L g1068 ( .A(n_156), .B(n_1069), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_157), .A2(n_240), .B1(n_492), .B2(n_496), .C(n_497), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_158), .A2(n_164), .B1(n_1025), .B2(n_1135), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_159), .A2(n_282), .B1(n_796), .B2(n_832), .C(n_1229), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_159), .A2(n_285), .B1(n_432), .B2(n_724), .Y(n_1368) );
INVx1_ASAP7_75t_L g1121 ( .A(n_160), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1259 ( .A1(n_161), .A2(n_247), .B1(n_732), .B2(n_1022), .Y(n_1259) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_162), .A2(n_372), .B1(n_752), .B2(n_755), .Y(n_772) );
INVxp33_ASAP7_75t_SL g814 ( .A(n_162), .Y(n_814) );
AO22x1_ASAP7_75t_L g1648 ( .A1(n_163), .A2(n_363), .B1(n_1625), .B2(n_1628), .Y(n_1648) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_164), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_165), .Y(n_775) );
OA21x2_ASAP7_75t_L g1299 ( .A1(n_166), .A2(n_449), .B(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g779 ( .A(n_167), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_167), .A2(n_265), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_168), .A2(n_193), .B1(n_1025), .B2(n_1077), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_168), .A2(n_213), .B1(n_497), .B2(n_1040), .C(n_1107), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_169), .A2(n_321), .B1(n_580), .B2(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1111 ( .A(n_169), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_170), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_171), .A2(n_183), .B1(n_669), .B2(n_690), .C(n_691), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_171), .A2(n_356), .B1(n_723), .B2(n_724), .C(n_725), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g1475 ( .A1(n_172), .A2(n_326), .B1(n_1476), .B2(n_1477), .Y(n_1475) );
OAI22xp33_ASAP7_75t_L g1483 ( .A1(n_172), .A2(n_326), .B1(n_1484), .B2(n_1487), .Y(n_1483) );
INVx1_ASAP7_75t_L g1346 ( .A(n_173), .Y(n_1346) );
INVx1_ASAP7_75t_L g1029 ( .A(n_174), .Y(n_1029) );
OAI211xp5_ASAP7_75t_L g1864 ( .A1(n_175), .A2(n_1865), .B(n_1866), .C(n_1867), .Y(n_1864) );
INVx1_ASAP7_75t_L g1885 ( .A(n_175), .Y(n_1885) );
INVx1_ASAP7_75t_L g1292 ( .A(n_176), .Y(n_1292) );
AO22x1_ASAP7_75t_L g1164 ( .A1(n_177), .A2(n_219), .B1(n_1129), .B2(n_1130), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_177), .B(n_1098), .Y(n_1189) );
INVx1_ASAP7_75t_L g872 ( .A(n_178), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g1185 ( .A1(n_179), .A2(n_219), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
INVx1_ASAP7_75t_L g1868 ( .A(n_180), .Y(n_1868) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_181), .Y(n_1089) );
INVx1_ASAP7_75t_L g983 ( .A(n_182), .Y(n_983) );
AO22x1_ASAP7_75t_L g1617 ( .A1(n_184), .A2(n_365), .B1(n_1618), .B2(n_1622), .Y(n_1617) );
OA22x2_ASAP7_75t_L g1569 ( .A1(n_186), .A2(n_1570), .B1(n_1601), .B2(n_1602), .Y(n_1569) );
CKINVDCx16_ASAP7_75t_R g1601 ( .A(n_186), .Y(n_1601) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_187), .A2(n_364), .B1(n_533), .B2(n_593), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_188), .A2(n_312), .B1(n_533), .B2(n_593), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_189), .Y(n_958) );
OAI211xp5_ASAP7_75t_L g1385 ( .A1(n_190), .A2(n_613), .B(n_1386), .C(n_1388), .Y(n_1385) );
INVx1_ASAP7_75t_L g1408 ( .A(n_190), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1872 ( .A1(n_191), .A2(n_310), .B1(n_1873), .B2(n_1874), .Y(n_1872) );
OAI22xp33_ASAP7_75t_L g1886 ( .A1(n_191), .A2(n_310), .B1(n_1887), .B2(n_1888), .Y(n_1886) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_192), .Y(n_700) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_193), .Y(n_1095) );
INVx1_ASAP7_75t_L g899 ( .A(n_195), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_195), .A2(n_283), .B1(n_608), .B2(n_828), .Y(n_933) );
INVx1_ASAP7_75t_L g1589 ( .A(n_196), .Y(n_1589) );
INVx1_ASAP7_75t_L g692 ( .A(n_197), .Y(n_692) );
INVx1_ASAP7_75t_L g1847 ( .A(n_198), .Y(n_1847) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_199), .A2(n_294), .B1(n_1466), .B2(n_1470), .Y(n_1465) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_199), .A2(n_294), .B1(n_1505), .B2(n_1508), .Y(n_1504) );
AOI221xp5_ASAP7_75t_L g1036 ( .A1(n_200), .A2(n_241), .B1(n_606), .B2(n_1037), .C(n_1040), .Y(n_1036) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_201), .Y(n_957) );
INVx1_ASAP7_75t_L g968 ( .A(n_202), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g1128 ( .A1(n_203), .A2(n_295), .B1(n_1129), .B2(n_1130), .Y(n_1128) );
INVx1_ASAP7_75t_L g1309 ( .A(n_204), .Y(n_1309) );
AOI221xp5_ASAP7_75t_L g1336 ( .A1(n_204), .A2(n_242), .B1(n_1107), .B2(n_1229), .C(n_1242), .Y(n_1336) );
OAI211xp5_ASAP7_75t_L g822 ( .A1(n_205), .A2(n_823), .B(n_825), .C(n_833), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_205), .B(n_437), .Y(n_849) );
INVx1_ASAP7_75t_L g1587 ( .A(n_206), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_207), .A2(n_304), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
INVx1_ASAP7_75t_L g1828 ( .A(n_208), .Y(n_1828) );
INVx1_ASAP7_75t_L g1074 ( .A(n_209), .Y(n_1074) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_209), .A2(n_337), .B1(n_506), .B2(n_1093), .C(n_1094), .Y(n_1092) );
INVx2_ASAP7_75t_L g1621 ( .A(n_210), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_210), .B(n_319), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_210), .B(n_1627), .Y(n_1629) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_211), .Y(n_542) );
INVx1_ASAP7_75t_L g1335 ( .A(n_212), .Y(n_1335) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_213), .A2(n_315), .B1(n_641), .B2(n_723), .Y(n_1084) );
XNOR2xp5_ASAP7_75t_L g1382 ( .A(n_214), .B(n_1383), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_215), .A2(n_307), .B1(n_437), .B2(n_533), .Y(n_1220) );
OAI211xp5_ASAP7_75t_L g1222 ( .A1(n_215), .A2(n_523), .B(n_1223), .C(n_1233), .Y(n_1222) );
XOR2x2_ASAP7_75t_L g1517 ( .A(n_216), .B(n_1518), .Y(n_1517) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_217), .Y(n_1180) );
AOI221xp5_ASAP7_75t_L g1148 ( .A1(n_218), .A2(n_295), .B1(n_492), .B2(n_517), .C(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g940 ( .A(n_221), .Y(n_940) );
INVx1_ASAP7_75t_L g1028 ( .A(n_222), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_223), .A2(n_301), .B1(n_827), .B2(n_828), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_223), .A2(n_318), .B1(n_724), .B2(n_859), .Y(n_858) );
AOI21xp33_ASAP7_75t_L g1577 ( .A1(n_224), .A2(n_1529), .B(n_1578), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_224), .A2(n_342), .B1(n_732), .B2(n_870), .Y(n_1597) );
INVx1_ASAP7_75t_L g1911 ( .A(n_225), .Y(n_1911) );
OAI211xp5_ASAP7_75t_L g1572 ( .A1(n_226), .A2(n_613), .B(n_1573), .C(n_1575), .Y(n_1572) );
INVx1_ASAP7_75t_L g1594 ( .A(n_226), .Y(n_1594) );
INVx1_ASAP7_75t_L g1315 ( .A(n_227), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_227), .A2(n_292), .B1(n_828), .B2(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1005 ( .A(n_228), .Y(n_1005) );
INVx1_ASAP7_75t_L g1257 ( .A(n_229), .Y(n_1257) );
OAI211xp5_ASAP7_75t_L g1266 ( .A1(n_229), .A2(n_1102), .B(n_1267), .C(n_1274), .Y(n_1266) );
INVx1_ASAP7_75t_L g408 ( .A(n_230), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_231), .Y(n_901) );
INVx1_ASAP7_75t_L g435 ( .A(n_232), .Y(n_435) );
INVx1_ASAP7_75t_L g1836 ( .A(n_233), .Y(n_1836) );
INVx1_ASAP7_75t_L g583 ( .A(n_234), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_235), .Y(n_844) );
INVx2_ASAP7_75t_L g421 ( .A(n_236), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_236), .B(n_419), .Y(n_456) );
INVx1_ASAP7_75t_L g568 ( .A(n_236), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_237), .Y(n_1275) );
OAI211xp5_ASAP7_75t_L g1924 ( .A1(n_238), .A2(n_1102), .B(n_1925), .C(n_1929), .Y(n_1924) );
INVx1_ASAP7_75t_L g910 ( .A(n_239), .Y(n_910) );
NAND2xp33_ASAP7_75t_SL g934 ( .A(n_239), .B(n_478), .Y(n_934) );
INVx1_ASAP7_75t_L g560 ( .A(n_240), .Y(n_560) );
INVx1_ASAP7_75t_L g1314 ( .A(n_242), .Y(n_1314) );
INVx1_ASAP7_75t_L g1912 ( .A(n_243), .Y(n_1912) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_244), .A2(n_327), .B1(n_835), .B2(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g876 ( .A(n_244), .Y(n_876) );
INVx1_ASAP7_75t_L g490 ( .A(n_245), .Y(n_490) );
INVx1_ASAP7_75t_L g1281 ( .A(n_246), .Y(n_1281) );
INVx1_ASAP7_75t_L g1285 ( .A(n_247), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g911 ( .A1(n_248), .A2(n_651), .B(n_725), .Y(n_911) );
INVx1_ASAP7_75t_L g936 ( .A(n_249), .Y(n_936) );
BUFx3_ASAP7_75t_L g413 ( .A(n_250), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_251), .A2(n_296), .B1(n_723), .B2(n_990), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1394 ( .A1(n_252), .A2(n_279), .B1(n_606), .B2(n_1226), .C(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1538 ( .A(n_253), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1662 ( .A1(n_254), .A2(n_259), .B1(n_1625), .B2(n_1628), .Y(n_1662) );
XOR2xp5_ASAP7_75t_L g1823 ( .A(n_254), .B(n_1824), .Y(n_1823) );
AOI22xp33_ASAP7_75t_L g1893 ( .A1(n_254), .A2(n_1894), .B1(n_1897), .B2(n_1935), .Y(n_1893) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_256), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g1901 ( .A1(n_257), .A2(n_261), .B1(n_979), .B2(n_1902), .Y(n_1901) );
OAI221xp5_ASAP7_75t_L g1921 ( .A1(n_257), .A2(n_261), .B1(n_613), .B2(n_614), .C(n_1922), .Y(n_1921) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_258), .A2(n_313), .B1(n_572), .B2(n_646), .Y(n_1082) );
INVx1_ASAP7_75t_L g892 ( .A(n_260), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_260), .B(n_752), .Y(n_894) );
AOI21xp33_ASAP7_75t_L g971 ( .A1(n_262), .A2(n_517), .B(n_797), .Y(n_971) );
INVx1_ASAP7_75t_L g982 ( .A(n_262), .Y(n_982) );
INVx1_ASAP7_75t_L g1831 ( .A(n_263), .Y(n_1831) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_265), .A2(n_572), .B(n_730), .Y(n_791) );
XOR2x2_ASAP7_75t_L g945 ( .A(n_266), .B(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_267), .A2(n_284), .B1(n_1046), .B2(n_1105), .Y(n_1579) );
OAI22xp33_ASAP7_75t_L g1216 ( .A1(n_268), .A2(n_288), .B1(n_580), .B2(n_630), .Y(n_1216) );
INVx1_ASAP7_75t_L g1234 ( .A(n_268), .Y(n_1234) );
CKINVDCx5p33_ASAP7_75t_R g1422 ( .A(n_269), .Y(n_1422) );
BUFx3_ASAP7_75t_L g398 ( .A(n_271), .Y(n_398) );
INVx1_ASAP7_75t_L g477 ( .A(n_271), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g1706 ( .A(n_272), .Y(n_1706) );
AOI22xp5_ASAP7_75t_L g1650 ( .A1(n_273), .A2(n_289), .B1(n_1625), .B2(n_1628), .Y(n_1650) );
INVx1_ASAP7_75t_L g1543 ( .A(n_274), .Y(n_1543) );
NAND2xp5_ASAP7_75t_SL g963 ( .A(n_276), .B(n_797), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_278), .A2(n_342), .B1(n_1046), .B2(n_1398), .Y(n_1584) );
AOI22xp33_ASAP7_75t_SL g1599 ( .A1(n_278), .A2(n_353), .B1(n_582), .B2(n_1130), .Y(n_1599) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_280), .Y(n_781) );
INVx1_ASAP7_75t_L g908 ( .A(n_283), .Y(n_908) );
INVx1_ASAP7_75t_L g1208 ( .A(n_287), .Y(n_1208) );
INVx1_ASAP7_75t_L g1235 ( .A(n_288), .Y(n_1235) );
INVx1_ASAP7_75t_L g483 ( .A(n_290), .Y(n_483) );
INVx1_ASAP7_75t_L g654 ( .A(n_291), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g1311 ( .A(n_292), .B(n_1016), .Y(n_1311) );
NAND2xp5_ASAP7_75t_SL g966 ( .A(n_296), .B(n_496), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g1643 ( .A1(n_297), .A2(n_368), .B1(n_1625), .B2(n_1628), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_298), .A2(n_341), .B1(n_1046), .B2(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g763 ( .A(n_299), .Y(n_763) );
AO22x1_ASAP7_75t_L g1647 ( .A1(n_299), .A2(n_306), .B1(n_1618), .B2(n_1632), .Y(n_1647) );
XNOR2x2_ASAP7_75t_L g1202 ( .A(n_300), .B(n_1203), .Y(n_1202) );
AOI22xp33_ASAP7_75t_SL g852 ( .A1(n_301), .A2(n_374), .B1(n_724), .B2(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1919 ( .A(n_302), .Y(n_1919) );
INVx1_ASAP7_75t_L g429 ( .A(n_303), .Y(n_429) );
INVx1_ASAP7_75t_L g443 ( .A(n_303), .Y(n_443) );
INVx1_ASAP7_75t_L g1332 ( .A(n_308), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_309), .Y(n_1117) );
INVx1_ASAP7_75t_L g1286 ( .A(n_311), .Y(n_1286) );
OAI211xp5_ASAP7_75t_L g1137 ( .A1(n_312), .A2(n_1102), .B(n_1138), .C(n_1143), .Y(n_1137) );
OAI21xp33_ASAP7_75t_L g974 ( .A1(n_314), .A2(n_868), .B(n_975), .Y(n_974) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_315), .Y(n_1096) );
INVx1_ASAP7_75t_L g693 ( .A(n_316), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_317), .Y(n_891) );
AOI221xp5_ASAP7_75t_SL g831 ( .A1(n_318), .A2(n_374), .B1(n_478), .B2(n_605), .C(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_319), .B(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1627 ( .A(n_319), .Y(n_1627) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_320), .Y(n_623) );
INVx1_ASAP7_75t_L g1112 ( .A(n_321), .Y(n_1112) );
INVx1_ASAP7_75t_L g1534 ( .A(n_322), .Y(n_1534) );
INVx1_ASAP7_75t_L g1361 ( .A(n_323), .Y(n_1361) );
INVx1_ASAP7_75t_L g1931 ( .A(n_325), .Y(n_1931) );
INVx1_ASAP7_75t_L g865 ( .A(n_327), .Y(n_865) );
INVx1_ASAP7_75t_L g1558 ( .A(n_328), .Y(n_1558) );
XNOR2xp5_ASAP7_75t_L g764 ( .A(n_329), .B(n_765), .Y(n_764) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_331), .Y(n_573) );
INVx1_ASAP7_75t_L g1401 ( .A(n_332), .Y(n_1401) );
INVx1_ASAP7_75t_L g1360 ( .A(n_333), .Y(n_1360) );
CKINVDCx16_ASAP7_75t_R g914 ( .A(n_334), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_336), .Y(n_1437) );
INVx1_ASAP7_75t_L g1073 ( .A(n_337), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_338), .B(n_1244), .Y(n_1243) );
OAI21xp33_ASAP7_75t_L g1026 ( .A1(n_339), .A2(n_533), .B(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g767 ( .A(n_340), .Y(n_767) );
INVx1_ASAP7_75t_L g787 ( .A(n_343), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g1424 ( .A(n_344), .Y(n_1424) );
INVx1_ASAP7_75t_L g1869 ( .A(n_345), .Y(n_1869) );
OAI211xp5_ASAP7_75t_L g1881 ( .A1(n_345), .A2(n_1551), .B(n_1882), .C(n_1883), .Y(n_1881) );
XNOR2xp5_ASAP7_75t_L g1898 ( .A(n_346), .B(n_1899), .Y(n_1898) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_347), .Y(n_1201) );
OAI211xp5_ASAP7_75t_L g1521 ( .A1(n_348), .A2(n_472), .B(n_499), .C(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1565 ( .A(n_348), .Y(n_1565) );
AOI221xp5_ASAP7_75t_L g1528 ( .A1(n_349), .A2(n_371), .B1(n_1226), .B2(n_1242), .C(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1541 ( .A(n_349), .Y(n_1541) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_350), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_350), .A2(n_359), .B1(n_641), .B2(n_642), .Y(n_640) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_352), .Y(n_394) );
INVxp67_ASAP7_75t_SL g1576 ( .A(n_353), .Y(n_1576) );
INVx1_ASAP7_75t_L g1842 ( .A(n_354), .Y(n_1842) );
NOR2xp33_ASAP7_75t_R g927 ( .A(n_355), .B(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g887 ( .A(n_357), .Y(n_887) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_361), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_361), .A2(n_362), .B1(n_744), .B2(n_746), .C(n_748), .Y(n_743) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_362), .A2(n_366), .B1(n_681), .B2(n_686), .C(n_687), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g1101 ( .A1(n_364), .A2(n_1102), .B(n_1103), .C(n_1110), .Y(n_1101) );
XOR2x2_ASAP7_75t_L g1114 ( .A(n_365), .B(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g416 ( .A(n_367), .Y(n_416) );
INVx1_ASAP7_75t_L g447 ( .A(n_367), .Y(n_447) );
INVx2_ASAP7_75t_L g530 ( .A(n_367), .Y(n_530) );
INVx1_ASAP7_75t_L g800 ( .A(n_369), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g1933 ( .A(n_370), .Y(n_1933) );
INVxp67_ASAP7_75t_SL g1554 ( .A(n_371), .Y(n_1554) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_372), .Y(n_770) );
INVx1_ASAP7_75t_L g1253 ( .A(n_373), .Y(n_1253) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_399), .B(n_1608), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_384), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g1892 ( .A(n_378), .B(n_387), .Y(n_1892) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g1896 ( .A(n_380), .B(n_383), .Y(n_1896) );
INVx1_ASAP7_75t_L g1938 ( .A(n_380), .Y(n_1938) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1941 ( .A(n_383), .B(n_1938), .Y(n_1941) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g1480 ( .A(n_387), .B(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g498 ( .A(n_388), .B(n_398), .Y(n_498) );
AND2x4_ASAP7_75t_L g518 ( .A(n_388), .B(n_397), .Y(n_518) );
INVx1_ASAP7_75t_L g1476 ( .A(n_389), .Y(n_1476) );
AND2x4_ASAP7_75t_SL g1891 ( .A(n_389), .B(n_1892), .Y(n_1891) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_396), .Y(n_390) );
INVxp67_ASAP7_75t_L g1244 ( .A(n_391), .Y(n_1244) );
OR2x6_ASAP7_75t_L g1468 ( .A(n_391), .B(n_1469), .Y(n_1468) );
BUFx4f_ASAP7_75t_L g1854 ( .A(n_391), .Y(n_1854) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g482 ( .A(n_392), .Y(n_482) );
BUFx4f_ASAP7_75t_L g836 ( .A(n_392), .Y(n_836) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g461 ( .A(n_394), .Y(n_461) );
AND2x2_ASAP7_75t_L g479 ( .A(n_394), .B(n_395), .Y(n_479) );
INVx2_ASAP7_75t_L g489 ( .A(n_394), .Y(n_489) );
AND2x2_ASAP7_75t_L g494 ( .A(n_394), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g537 ( .A(n_394), .Y(n_537) );
NAND2x1_ASAP7_75t_L g677 ( .A(n_394), .B(n_395), .Y(n_677) );
INVx1_ASAP7_75t_L g462 ( .A(n_395), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_395), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g495 ( .A(n_395), .Y(n_495) );
BUFx2_ASAP7_75t_L g509 ( .A(n_395), .Y(n_509) );
AND2x2_ASAP7_75t_L g526 ( .A(n_395), .B(n_489), .Y(n_526) );
OR2x2_ASAP7_75t_L g673 ( .A(n_395), .B(n_461), .Y(n_673) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g1456 ( .A(n_397), .Y(n_1456) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g1460 ( .A(n_398), .Y(n_1460) );
AND2x4_ASAP7_75t_L g1464 ( .A(n_398), .B(n_536), .Y(n_1464) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_1153), .B2(n_1607), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_658), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_584), .B2(n_585), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
XNOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_583), .Y(n_404) );
NOR2x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_469), .Y(n_405) );
NAND5xp2_ASAP7_75t_L g406 ( .A(n_407), .B(n_430), .C(n_434), .D(n_448), .E(n_463), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_422), .B2(n_423), .Y(n_407) );
AO22x1_ASAP7_75t_L g1003 ( .A1(n_409), .A2(n_423), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_409), .A2(n_423), .B1(n_1175), .B2(n_1176), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_409), .A2(n_423), .B1(n_1207), .B2(n_1208), .Y(n_1206) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
AND2x2_ASAP7_75t_L g655 ( .A(n_410), .B(n_414), .Y(n_655) );
AND2x6_ASAP7_75t_L g745 ( .A(n_410), .B(n_417), .Y(n_745) );
AND2x4_ASAP7_75t_SL g863 ( .A(n_410), .B(n_414), .Y(n_863) );
NAND2x1_ASAP7_75t_L g979 ( .A(n_410), .B(n_414), .Y(n_979) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_412), .B(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g647 ( .A(n_412), .B(n_427), .Y(n_647) );
BUFx2_ASAP7_75t_L g1499 ( .A(n_412), .Y(n_1499) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g433 ( .A(n_413), .B(n_428), .Y(n_433) );
INVx2_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_413), .B(n_429), .Y(n_453) );
OR2x2_ASAP7_75t_L g559 ( .A(n_413), .B(n_442), .Y(n_559) );
AND2x4_ASAP7_75t_L g423 ( .A(n_414), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g431 ( .A(n_414), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_SL g864 ( .A(n_414), .B(n_424), .Y(n_864) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
OR2x2_ASAP7_75t_L g457 ( .A(n_415), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g698 ( .A(n_415), .Y(n_698) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g567 ( .A(n_416), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_416), .B(n_476), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_417), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g747 ( .A(n_417), .B(n_426), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_417), .Y(n_750) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
NAND3x1_ASAP7_75t_L g566 ( .A(n_418), .B(n_567), .C(n_568), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g725 ( .A(n_418), .B(n_568), .Y(n_725) );
OR2x4_ASAP7_75t_L g1486 ( .A(n_418), .B(n_559), .Y(n_1486) );
INVx1_ASAP7_75t_L g1489 ( .A(n_418), .Y(n_1489) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_418), .B(n_433), .Y(n_1494) );
OR2x6_ASAP7_75t_L g1509 ( .A(n_418), .B(n_575), .Y(n_1509) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_419), .B(n_421), .Y(n_554) );
BUFx3_ASAP7_75t_L g638 ( .A(n_419), .Y(n_638) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND3x4_ASAP7_75t_L g637 ( .A(n_421), .B(n_638), .C(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g903 ( .A(n_421), .B(n_638), .Y(n_903) );
HB1xp67_ASAP7_75t_L g1512 ( .A(n_421), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_423), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
AOI221x1_ASAP7_75t_L g977 ( .A1(n_423), .A2(n_950), .B1(n_957), .B2(n_978), .C(n_980), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_423), .A2(n_978), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_423), .A2(n_978), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_423), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_423), .A2(n_978), .B1(n_1531), .B2(n_1565), .Y(n_1564) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g541 ( .A(n_429), .Y(n_541) );
AND4x1_ASAP7_75t_L g627 ( .A(n_430), .B(n_628), .C(n_636), .D(n_653), .Y(n_627) );
AND5x1_ASAP7_75t_L g946 ( .A(n_430), .B(n_947), .C(n_977), .D(n_991), .E(n_994), .Y(n_946) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_430), .Y(n_1087) );
NAND4xp75_ASAP7_75t_L g1115 ( .A(n_430), .B(n_1116), .C(n_1119), .D(n_1136), .Y(n_1115) );
AND4x1_ASAP7_75t_L g1251 ( .A(n_430), .B(n_1252), .C(n_1256), .D(n_1258), .Y(n_1251) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_431), .A2(n_841), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_862) );
INVx3_ASAP7_75t_L g1009 ( .A(n_431), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_431), .Y(n_1217) );
NOR3xp33_ASAP7_75t_SL g1305 ( .A(n_431), .B(n_1306), .C(n_1317), .Y(n_1305) );
AOI211xp5_ASAP7_75t_L g1364 ( .A1(n_431), .A2(n_436), .B(n_1356), .C(n_1365), .Y(n_1364) );
NOR3xp33_ASAP7_75t_L g1591 ( .A(n_431), .B(n_1592), .C(n_1600), .Y(n_1591) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_432), .Y(n_1167) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g579 ( .A(n_433), .Y(n_579) );
BUFx2_ASAP7_75t_L g642 ( .A(n_433), .Y(n_642) );
BUFx3_ASAP7_75t_L g723 ( .A(n_433), .Y(n_723) );
AND2x2_ASAP7_75t_L g738 ( .A(n_433), .B(n_736), .Y(n_738) );
BUFx2_ASAP7_75t_L g853 ( .A(n_433), .Y(n_853) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_433), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_436), .B(n_1173), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_436), .A2(n_1301), .B1(n_1302), .B2(n_1304), .Y(n_1300) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx5_ASAP7_75t_L g996 ( .A(n_437), .Y(n_996) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_444), .Y(n_437) );
OR2x2_ASAP7_75t_L g593 ( .A(n_438), .B(n_444), .Y(n_593) );
INVx2_ASAP7_75t_L g742 ( .A(n_438), .Y(n_742) );
INVx8_ASAP7_75t_L g467 ( .A(n_439), .Y(n_467) );
BUFx3_ASAP7_75t_L g641 ( .A(n_439), .Y(n_641) );
BUFx3_ASAP7_75t_L g651 ( .A(n_439), .Y(n_651) );
AND2x2_ASAP7_75t_L g735 ( .A(n_439), .B(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_439), .Y(n_990) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x4_ASAP7_75t_L g548 ( .A(n_440), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g549 ( .A(n_443), .Y(n_549) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g534 ( .A(n_445), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g686 ( .A(n_445), .B(n_535), .Y(n_686) );
INVx1_ASAP7_75t_L g715 ( .A(n_445), .Y(n_715) );
INVx1_ASAP7_75t_L g1481 ( .A(n_445), .Y(n_1481) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g455 ( .A(n_446), .Y(n_455) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx8_ASAP7_75t_L g590 ( .A(n_449), .Y(n_590) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_457), .Y(n_449) );
INVx1_ASAP7_75t_L g877 ( .A(n_450), .Y(n_877) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
BUFx3_ASAP7_75t_L g780 ( .A(n_451), .Y(n_780) );
INVx1_ASAP7_75t_L g1545 ( .A(n_451), .Y(n_1545) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_452), .Y(n_551) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g575 ( .A(n_453), .Y(n_575) );
INVx1_ASAP7_75t_L g468 ( .A(n_454), .Y(n_468) );
OR2x2_ASAP7_75t_L g538 ( .A(n_454), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g634 ( .A(n_454), .Y(n_634) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OR2x2_ASAP7_75t_L g553 ( .A(n_455), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_455), .B(n_498), .Y(n_679) );
INVx1_ASAP7_75t_L g808 ( .A(n_455), .Y(n_808) );
HB1xp67_ASAP7_75t_L g1514 ( .A(n_455), .Y(n_1514) );
INVx1_ASAP7_75t_L g736 ( .A(n_456), .Y(n_736) );
INVx1_ASAP7_75t_L g754 ( .A(n_456), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_457), .B(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g699 ( .A(n_458), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
AND2x6_ASAP7_75t_L g500 ( .A(n_459), .B(n_478), .Y(n_500) );
INVx1_ASAP7_75t_L g510 ( .A(n_459), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_459), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_459), .B(n_530), .Y(n_683) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_459), .B(n_840), .Y(n_1197) );
AND2x2_ASAP7_75t_L g522 ( .A(n_460), .B(n_476), .Y(n_522) );
INVx3_ASAP7_75t_L g609 ( .A(n_460), .Y(n_609) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_460), .Y(n_827) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_461), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_465), .A2(n_581), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_465), .A2(n_581), .B1(n_1180), .B2(n_1181), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_465), .A2(n_581), .B1(n_1275), .B2(n_1277), .Y(n_1289) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_465), .A2(n_1327), .B1(n_1328), .B2(n_1339), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_465), .A2(n_869), .B1(n_1360), .B2(n_1361), .Y(n_1363) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
AND2x4_ASAP7_75t_L g875 ( .A(n_466), .B(n_468), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_466), .A2(n_859), .B1(n_891), .B2(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g577 ( .A(n_467), .Y(n_577) );
INVx8_ASAP7_75t_L g724 ( .A(n_467), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_467), .Y(n_783) );
INVx3_ASAP7_75t_L g1022 ( .A(n_467), .Y(n_1022) );
AND2x4_ASAP7_75t_L g581 ( .A(n_468), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_531), .Y(n_469) );
OAI31xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_501), .A3(n_519), .B(n_527), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g613 ( .A(n_473), .Y(n_613) );
INVx2_ASAP7_75t_L g1093 ( .A(n_473), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_473), .A2(n_507), .B1(n_1207), .B2(n_1208), .Y(n_1245) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g951 ( .A(n_475), .Y(n_951) );
AND2x4_ASAP7_75t_SL g475 ( .A(n_476), .B(n_478), .Y(n_475) );
AND2x4_ASAP7_75t_L g504 ( .A(n_476), .B(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g524 ( .A(n_476), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g762 ( .A(n_476), .B(n_505), .Y(n_762) );
AND2x2_ASAP7_75t_L g824 ( .A(n_476), .B(n_704), .Y(n_824) );
BUFx2_ASAP7_75t_L g846 ( .A(n_476), .Y(n_846) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_477), .Y(n_1469) );
BUFx3_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
BUFx3_ASAP7_75t_L g516 ( .A(n_478), .Y(n_516) );
INVx1_ASAP7_75t_L g602 ( .A(n_478), .Y(n_602) );
BUFx3_ASAP7_75t_L g796 ( .A(n_478), .Y(n_796) );
BUFx6f_ASAP7_75t_L g1226 ( .A(n_478), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_478), .B(n_1456), .Y(n_1455) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g1039 ( .A(n_479), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B1(n_484), .B2(n_490), .C(n_491), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_481), .A2(n_512), .B1(n_513), .B2(n_514), .C(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g669 ( .A(n_481), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_481), .A2(n_621), .B1(n_1146), .B2(n_1147), .C(n_1148), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_481), .A2(n_620), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
OAI221xp5_ASAP7_75t_SL g1922 ( .A1(n_481), .A2(n_620), .B1(n_1911), .B2(n_1918), .C(n_1923), .Y(n_1922) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g618 ( .A(n_482), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_482), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_798) );
OAI22x1_ASAP7_75t_SL g804 ( .A1(n_482), .A2(n_781), .B1(n_801), .B2(n_805), .Y(n_804) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_482), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_483), .A2(n_545), .B1(n_546), .B2(n_550), .Y(n_544) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g622 ( .A(n_486), .Y(n_622) );
INVx2_ASAP7_75t_L g801 ( .A(n_486), .Y(n_801) );
INVx4_ASAP7_75t_L g961 ( .A(n_486), .Y(n_961) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_486), .Y(n_1061) );
INVx1_ASAP7_75t_L g1334 ( .A(n_486), .Y(n_1334) );
INVx8_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g513 ( .A(n_487), .Y(n_513) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_487), .B(n_1460), .Y(n_1474) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_490), .A2(n_570), .B1(n_573), .B2(n_574), .C(n_576), .Y(n_569) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g605 ( .A(n_493), .Y(n_605) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
BUFx3_ASAP7_75t_L g797 ( .A(n_494), .Y(n_797) );
AND2x4_ASAP7_75t_L g1478 ( .A(n_494), .B(n_1469), .Y(n_1478) );
HB1xp67_ASAP7_75t_SL g1927 ( .A(n_497), .Y(n_1927) );
INVx4_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g606 ( .A(n_498), .Y(n_606) );
AND2x4_ASAP7_75t_L g806 ( .A(n_498), .B(n_807), .Y(n_806) );
INVx4_ASAP7_75t_L g832 ( .A(n_498), .Y(n_832) );
NAND4xp25_ASAP7_75t_L g962 ( .A(n_498), .B(n_963), .C(n_964), .D(n_966), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_498), .B(n_807), .Y(n_1451) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_500), .A2(n_600), .B(n_607), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_500), .A2(n_1036), .B(n_1042), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g1103 ( .A1(n_500), .A2(n_1104), .B(n_1106), .Y(n_1103) );
AOI21xp5_ASAP7_75t_SL g1138 ( .A1(n_500), .A2(n_1139), .B(n_1142), .Y(n_1138) );
AOI221xp5_ASAP7_75t_SL g1182 ( .A1(n_500), .A2(n_524), .B1(n_1173), .B2(n_1183), .C(n_1185), .Y(n_1182) );
AOI21xp5_ASAP7_75t_L g1223 ( .A1(n_500), .A2(n_1224), .B(n_1230), .Y(n_1223) );
AOI21xp5_ASAP7_75t_L g1267 ( .A1(n_500), .A2(n_1268), .B(n_1269), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_500), .A2(n_824), .B1(n_1304), .B2(n_1323), .C(n_1324), .Y(n_1322) );
AOI221xp5_ASAP7_75t_L g1355 ( .A1(n_500), .A2(n_824), .B1(n_1356), .B2(n_1357), .C(n_1358), .Y(n_1355) );
AOI21xp5_ASAP7_75t_L g1393 ( .A1(n_500), .A2(n_1394), .B(n_1397), .Y(n_1393) );
AOI21xp5_ASAP7_75t_L g1581 ( .A1(n_500), .A2(n_1582), .B(n_1584), .Y(n_1581) );
AOI21xp5_ASAP7_75t_L g1925 ( .A1(n_500), .A2(n_1926), .B(n_1928), .Y(n_1925) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_503), .A2(n_521), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_503), .A2(n_1033), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_503), .A2(n_521), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_503), .A2(n_1033), .B1(n_1586), .B2(n_1587), .Y(n_1585) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_504), .A2(n_1028), .B1(n_1029), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_504), .A2(n_521), .B1(n_1124), .B2(n_1125), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_504), .A2(n_521), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
INVx1_ASAP7_75t_L g1237 ( .A(n_504), .Y(n_1237) );
HB1xp67_ASAP7_75t_L g1276 ( .A(n_504), .Y(n_1276) );
AOI22xp5_ASAP7_75t_L g1326 ( .A1(n_504), .A2(n_521), .B1(n_1327), .B2(n_1328), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_504), .A2(n_521), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_504), .A2(n_824), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_505), .Y(n_1041) );
INVx2_ASAP7_75t_L g1100 ( .A(n_505), .Y(n_1100) );
INVx1_ASAP7_75t_L g1530 ( .A(n_505), .Y(n_1530) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g615 ( .A(n_507), .Y(n_615) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g685 ( .A(n_509), .Y(n_685) );
BUFx2_ASAP7_75t_L g840 ( .A(n_509), .Y(n_840) );
AND2x4_ASAP7_75t_L g1459 ( .A(n_509), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g845 ( .A(n_510), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_512), .A2(n_556), .B1(n_560), .B2(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g690 ( .A(n_513), .Y(n_690) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g626 ( .A(n_518), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_518), .A2(n_675), .B1(n_1050), .B2(n_1051), .C(n_1054), .Y(n_1049) );
INVx2_ASAP7_75t_L g1242 ( .A(n_518), .Y(n_1242) );
INVx1_ASAP7_75t_L g1578 ( .A(n_518), .Y(n_1578) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_521), .B(n_1536), .Y(n_1535) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g714 ( .A(n_522), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1034 ( .A(n_522), .Y(n_1034) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_R g1047 ( .A(n_524), .B(n_1008), .Y(n_1047) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_524), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_525), .Y(n_1187) );
INVx1_ASAP7_75t_L g1273 ( .A(n_525), .Y(n_1273) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g611 ( .A(n_526), .Y(n_611) );
BUFx3_ASAP7_75t_L g828 ( .A(n_526), .Y(n_828) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_526), .Y(n_1046) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_527), .A2(n_595), .B(n_612), .Y(n_594) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_528), .B(n_756), .Y(n_942) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_528), .Y(n_1063) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g694 ( .A(n_529), .B(n_695), .Y(n_694) );
OR2x6_ASAP7_75t_L g861 ( .A(n_529), .B(n_725), .Y(n_861) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g639 ( .A(n_530), .Y(n_639) );
AOI21xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_542), .B(n_543), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g1537 ( .A1(n_532), .A2(n_1538), .B(n_1539), .Y(n_1537) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g1288 ( .A(n_533), .Y(n_1288) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
INVx2_ASAP7_75t_SL g812 ( .A(n_534), .Y(n_812) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_534), .B(n_538), .Y(n_1303) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g874 ( .A(n_538), .Y(n_874) );
INVx3_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
INVx4_ASAP7_75t_L g1552 ( .A(n_539), .Y(n_1552) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g749 ( .A(n_540), .Y(n_749) );
BUFx3_ASAP7_75t_L g1433 ( .A(n_540), .Y(n_1433) );
BUFx2_ASAP7_75t_L g1502 ( .A(n_541), .Y(n_1502) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g645 ( .A(n_547), .Y(n_645) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_547), .Y(n_855) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_547), .Y(n_857) );
INVx2_ASAP7_75t_L g1372 ( .A(n_547), .Y(n_1372) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_547), .B(n_1489), .Y(n_1488) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
BUFx8_ASAP7_75t_L g582 ( .A(n_548), .Y(n_582) );
INVx2_ASAP7_75t_L g720 ( .A(n_548), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_550), .A2(n_905), .B1(n_982), .B2(n_983), .C(n_984), .Y(n_981) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g898 ( .A(n_551), .Y(n_898) );
INVx3_ASAP7_75t_L g907 ( .A(n_551), .Y(n_907) );
CKINVDCx8_ASAP7_75t_R g1843 ( .A(n_551), .Y(n_1843) );
OAI22xp5_ASAP7_75t_SL g980 ( .A1(n_552), .A2(n_981), .B1(n_985), .B2(n_987), .Y(n_980) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx4f_ASAP7_75t_L g1307 ( .A(n_553), .Y(n_1307) );
BUFx4f_ASAP7_75t_L g1420 ( .A(n_553), .Y(n_1420) );
BUFx8_ASAP7_75t_L g1546 ( .A(n_553), .Y(n_1546) );
BUFx2_ASAP7_75t_L g730 ( .A(n_554), .Y(n_730) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_558), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_896) );
HB1xp67_ASAP7_75t_L g1423 ( .A(n_558), .Y(n_1423) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g632 ( .A(n_559), .Y(n_632) );
OR2x4_ASAP7_75t_L g1507 ( .A(n_559), .B(n_1489), .Y(n_1507) );
BUFx3_ASAP7_75t_L g1548 ( .A(n_559), .Y(n_1548) );
BUFx3_ASAP7_75t_L g1559 ( .A(n_559), .Y(n_1559) );
OAI22xp33_ASAP7_75t_L g1905 ( .A1(n_561), .A2(n_907), .B1(n_1906), .B2(n_1907), .Y(n_1905) );
OAI22xp33_ASAP7_75t_L g1917 ( .A1(n_561), .A2(n_1909), .B1(n_1918), .B2(n_1919), .Y(n_1917) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g790 ( .A(n_562), .Y(n_790) );
INVx2_ASAP7_75t_L g1425 ( .A(n_562), .Y(n_1425) );
OAI33xp33_ASAP7_75t_L g1904 ( .A1(n_563), .A2(n_1546), .A3(n_1905), .B1(n_1908), .B2(n_1913), .B3(n_1917), .Y(n_1904) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI33xp33_ASAP7_75t_L g636 ( .A1(n_564), .A2(n_637), .A3(n_640), .B1(n_643), .B2(n_648), .B3(n_649), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g1168 ( .A(n_564), .B(n_1169), .C(n_1170), .Y(n_1168) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_565), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_565), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_565), .Y(n_1214) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g986 ( .A(n_566), .Y(n_986) );
INVx1_ASAP7_75t_L g1261 ( .A(n_570), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1908 ( .A1(n_570), .A2(n_1909), .B1(n_1911), .B2(n_1912), .Y(n_1908) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_571), .A2(n_780), .B1(n_968), .B2(n_988), .C(n_989), .Y(n_987) );
INVx8_ASAP7_75t_L g1213 ( .A(n_571), .Y(n_1213) );
INVx5_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g729 ( .A(n_572), .Y(n_729) );
INVx2_ASAP7_75t_SL g905 ( .A(n_572), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g1312 ( .A1(n_574), .A2(n_1313), .B1(n_1314), .B2(n_1315), .C(n_1316), .Y(n_1312) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g1839 ( .A(n_575), .Y(n_1839) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g652 ( .A(n_579), .Y(n_652) );
INVx2_ASAP7_75t_L g727 ( .A(n_579), .Y(n_727) );
INVx2_ASAP7_75t_L g859 ( .A(n_579), .Y(n_859) );
INVxp67_ASAP7_75t_L g1339 ( .A(n_580), .Y(n_1339) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g635 ( .A(n_581), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_581), .A2(n_875), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_581), .B(n_1533), .Y(n_1567) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_582), .Y(n_1129) );
INVx3_ASAP7_75t_L g1542 ( .A(n_582), .Y(n_1542) );
INVx2_ASAP7_75t_SL g1914 ( .A(n_582), .Y(n_1914) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_657), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g588 ( .A(n_589), .B(n_594), .C(n_627), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
AOI211x1_ASAP7_75t_L g999 ( .A1(n_590), .A2(n_1000), .B(n_1001), .C(n_1026), .Y(n_999) );
AOI21xp33_ASAP7_75t_SL g1088 ( .A1(n_590), .A2(n_1089), .B(n_1090), .Y(n_1088) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_590), .A2(n_1117), .B(n_1118), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_590), .B(n_1201), .Y(n_1200) );
AOI21xp5_ASAP7_75t_L g1218 ( .A1(n_590), .A2(n_1219), .B(n_1220), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_590), .B(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_590), .B(n_1346), .Y(n_1345) );
AOI21xp33_ASAP7_75t_L g1402 ( .A1(n_590), .A2(n_1403), .B(n_1404), .Y(n_1402) );
AOI21xp5_ASAP7_75t_L g1588 ( .A1(n_590), .A2(n_1589), .B(n_1590), .Y(n_1588) );
AOI21xp33_ASAP7_75t_L g1932 ( .A1(n_590), .A2(n_1933), .B(n_1934), .Y(n_1932) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_593), .B(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g625 ( .A(n_602), .Y(n_625) );
INVx1_ASAP7_75t_L g1149 ( .A(n_602), .Y(n_1149) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g1141 ( .A(n_605), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1241 ( .A(n_605), .Y(n_1241) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g965 ( .A(n_609), .Y(n_965) );
INVx2_ASAP7_75t_L g1043 ( .A(n_609), .Y(n_1043) );
INVx1_ASAP7_75t_L g1105 ( .A(n_609), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1186 ( .A(n_609), .Y(n_1186) );
INVx2_ASAP7_75t_L g1231 ( .A(n_609), .Y(n_1231) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g704 ( .A(n_611), .Y(n_704) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_620), .B2(n_623), .C(n_624), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g1448 ( .A1(n_617), .A2(n_1280), .B1(n_1428), .B2(n_1434), .Y(n_1448) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g668 ( .A(n_621), .Y(n_668) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g1283 ( .A(n_626), .Y(n_1283) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_630), .B(n_713), .Y(n_993) );
OR2x6_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_631), .B(n_633), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1910 ( .A(n_631), .Y(n_1910) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g1830 ( .A(n_632), .Y(n_1830) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g869 ( .A(n_634), .B(n_870), .Y(n_869) );
AOI33xp33_ASAP7_75t_L g851 ( .A1(n_637), .A2(n_852), .A3(n_854), .B1(n_856), .B2(n_858), .B3(n_860), .Y(n_851) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_637), .Y(n_1011) );
AOI33xp33_ASAP7_75t_L g1075 ( .A1(n_637), .A2(n_1076), .A3(n_1079), .B1(n_1082), .B2(n_1083), .B3(n_1084), .Y(n_1075) );
AOI33xp33_ASAP7_75t_L g1367 ( .A1(n_637), .A2(n_1368), .A3(n_1369), .B1(n_1370), .B2(n_1373), .B3(n_1374), .Y(n_1367) );
AOI33xp33_ASAP7_75t_L g1409 ( .A1(n_637), .A2(n_1374), .A3(n_1410), .B1(n_1411), .B2(n_1412), .B3(n_1413), .Y(n_1409) );
AOI33xp33_ASAP7_75t_L g1595 ( .A1(n_637), .A2(n_1374), .A3(n_1596), .B1(n_1597), .B2(n_1598), .B3(n_1599), .Y(n_1595) );
INVx3_ASAP7_75t_L g1498 ( .A(n_638), .Y(n_1498) );
INVx1_ASAP7_75t_L g758 ( .A(n_639), .Y(n_758) );
OAI31xp33_ASAP7_75t_SL g771 ( .A1(n_639), .A2(n_772), .A3(n_773), .B(n_777), .Y(n_771) );
OAI31xp33_ASAP7_75t_L g893 ( .A1(n_639), .A2(n_894), .A3(n_895), .B(n_912), .Y(n_893) );
INVx2_ASAP7_75t_SL g1113 ( .A(n_639), .Y(n_1113) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_641), .Y(n_1014) );
INVx1_ASAP7_75t_L g1078 ( .A(n_641), .Y(n_1078) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_641), .Y(n_1135) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_645), .A2(n_907), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g721 ( .A(n_647), .Y(n_721) );
BUFx12f_ASAP7_75t_L g732 ( .A(n_647), .Y(n_732) );
AND2x4_ASAP7_75t_L g756 ( .A(n_647), .B(n_754), .Y(n_756) );
INVx5_ASAP7_75t_L g1017 ( .A(n_647), .Y(n_1017) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_647), .Y(n_1130) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g1318 ( .A(n_655), .Y(n_1318) );
AO22x2_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_1067), .B1(n_1151), .B2(n_1152), .Y(n_658) );
XOR2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_816), .Y(n_659) );
XNOR2x1_ASAP7_75t_L g1152 ( .A(n_660), .B(n_816), .Y(n_1152) );
BUFx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_764), .Y(n_662) );
XNOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_763), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_716), .Y(n_664) );
NAND3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_696), .C(n_710), .Y(n_665) );
AOI211xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_670), .B(n_680), .C(n_689), .Y(n_666) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_672), .A2(n_675), .B1(n_692), .B2(n_693), .C(n_694), .Y(n_691) );
BUFx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g932 ( .A(n_673), .Y(n_932) );
BUFx2_ASAP7_75t_L g960 ( .A(n_673), .Y(n_960) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_673), .Y(n_1053) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
BUFx4f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x6_ASAP7_75t_L g687 ( .A(n_676), .B(n_688), .Y(n_687) );
INVx4_ASAP7_75t_L g838 ( .A(n_676), .Y(n_838) );
BUFx4f_ASAP7_75t_L g848 ( .A(n_676), .Y(n_848) );
BUFx4f_ASAP7_75t_L g1859 ( .A(n_676), .Y(n_1859) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx3_ASAP7_75t_L g708 ( .A(n_677), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g929 ( .A1(n_678), .A2(n_687), .B(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g811 ( .A(n_681), .Y(n_811) );
INVx2_ASAP7_75t_SL g926 ( .A(n_681), .Y(n_926) );
NAND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g688 ( .A(n_682), .Y(n_688) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g924 ( .A(n_686), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_687), .Y(n_815) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_694), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_694), .B(n_921), .Y(n_920) );
INVx4_ASAP7_75t_L g1440 ( .A(n_694), .Y(n_1440) );
INVx2_ASAP7_75t_L g1852 ( .A(n_694), .Y(n_1852) );
AOI222xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B1(n_701), .B2(n_705), .C1(n_706), .C2(n_709), .Y(n_696) );
AOI21xp33_ASAP7_75t_SL g813 ( .A1(n_697), .A2(n_814), .B(n_815), .Y(n_813) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g809 ( .A1(n_701), .A2(n_775), .B1(n_787), .B2(n_810), .C1(n_811), .C2(n_812), .Y(n_809) );
INVx1_ASAP7_75t_L g938 ( .A(n_701), .Y(n_938) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g707 ( .A(n_703), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g928 ( .A(n_703), .B(n_708), .Y(n_928) );
AOI211xp5_ASAP7_75t_L g739 ( .A1(n_705), .A2(n_740), .B(n_743), .C(n_751), .Y(n_739) );
AOI222xp33_ASAP7_75t_L g794 ( .A1(n_706), .A2(n_776), .B1(n_795), .B2(n_802), .C1(n_803), .C2(n_806), .Y(n_794) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g970 ( .A(n_708), .Y(n_970) );
BUFx2_ASAP7_75t_SL g1280 ( .A(n_708), .Y(n_1280) );
BUFx3_ASAP7_75t_L g1865 ( .A(n_708), .Y(n_1865) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_714), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_714), .A2(n_761), .B1(n_891), .B2(n_892), .Y(n_890) );
AND2x4_ASAP7_75t_L g761 ( .A(n_715), .B(n_762), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_739), .B(n_757), .C(n_759), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .B1(n_726), .B2(n_731), .C(n_733), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OR2x6_ASAP7_75t_SL g752 ( .A(n_720), .B(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g870 ( .A(n_720), .Y(n_870) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_720), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1133 ( .A(n_720), .Y(n_1133) );
BUFx2_ASAP7_75t_L g1264 ( .A(n_724), .Y(n_1264) );
INVx3_ASAP7_75t_L g785 ( .A(n_725), .Y(n_785) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_729), .A2(n_779), .B1(n_780), .B2(n_781), .C(n_782), .Y(n_778) );
OAI221xp5_ASAP7_75t_L g900 ( .A1(n_729), .A2(n_749), .B1(n_901), .B2(n_902), .C(n_903), .Y(n_900) );
OAI22xp33_ASAP7_75t_SL g1834 ( .A1(n_729), .A2(n_1835), .B1(n_1836), .B2(n_1837), .Y(n_1834) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_732), .Y(n_1019) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_735), .A2(n_738), .B1(n_767), .B2(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx4_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_745), .A2(n_747), .B1(n_775), .B2(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g895 ( .A1(n_748), .A2(n_896), .B1(n_900), .B2(n_904), .C(n_909), .Y(n_895) );
OR2x6_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g1561 ( .A(n_749), .Y(n_1561) );
INVx1_ASAP7_75t_L g1833 ( .A(n_749), .Y(n_1833) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_754), .Y(n_916) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_757), .Y(n_973) );
INVx1_ASAP7_75t_L g1247 ( .A(n_757), .Y(n_1247) );
BUFx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI21x1_ASAP7_75t_L g821 ( .A1(n_758), .A2(n_822), .B(n_849), .Y(n_821) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_758), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_761), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g871 ( .A(n_761), .Y(n_871) );
AOI211x1_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B(n_768), .C(n_793), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_771), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_786), .C(n_788), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_780), .A2(n_1554), .B1(n_1555), .B2(n_1556), .Y(n_1553) );
INVx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_791), .C(n_792), .Y(n_788) );
OAI21xp5_ASAP7_75t_SL g909 ( .A1(n_790), .A2(n_910), .B(n_911), .Y(n_909) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_809), .C(n_813), .Y(n_793) );
INVx1_ASAP7_75t_L g1396 ( .A(n_797), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g1583 ( .A(n_797), .Y(n_1583) );
INVx2_ASAP7_75t_L g1860 ( .A(n_806), .Y(n_1860) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AO22x2_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_997), .B1(n_1065), .B2(n_1066), .Y(n_816) );
INVx1_ASAP7_75t_L g1065 ( .A(n_817), .Y(n_1065) );
XNOR2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_945), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_886), .B1(n_943), .B2(n_944), .Y(n_818) );
INVx1_ASAP7_75t_L g944 ( .A(n_819), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_879), .C(n_883), .Y(n_819) );
INVx1_ASAP7_75t_L g880 ( .A(n_821), .Y(n_880) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_825) );
INVx3_ASAP7_75t_L g1192 ( .A(n_827), .Y(n_1192) );
BUFx6f_ASAP7_75t_L g1271 ( .A(n_827), .Y(n_1271) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_833) );
INVx2_ASAP7_75t_SL g1443 ( .A(n_835), .Y(n_1443) );
INVx3_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx4_ASAP7_75t_L g954 ( .A(n_836), .Y(n_954) );
BUFx6f_ASAP7_75t_L g1058 ( .A(n_836), .Y(n_1058) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g955 ( .A(n_838), .Y(n_955) );
INVx1_ASAP7_75t_L g1857 ( .A(n_838), .Y(n_1857) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_841), .B1(n_842), .B2(n_844), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_840), .A2(n_842), .B1(n_957), .B2(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AOI222xp33_ASAP7_75t_L g873 ( .A1(n_844), .A2(n_874), .B1(n_875), .B2(n_876), .C1(n_877), .C2(n_878), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_845), .A2(n_846), .B1(n_953), .B2(n_959), .Y(n_952) );
OAI211xp5_ASAP7_75t_L g1388 ( .A1(n_848), .A2(n_1389), .B(n_1390), .C(n_1391), .Y(n_1388) );
OAI211xp5_ASAP7_75t_L g1575 ( .A1(n_848), .A2(n_1576), .B(n_1577), .C(n_1579), .Y(n_1575) );
INVx1_ASAP7_75t_L g881 ( .A(n_850), .Y(n_881) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_862), .Y(n_850) );
INVx2_ASAP7_75t_L g1555 ( .A(n_855), .Y(n_1555) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_SL g1374 ( .A(n_861), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_863), .A2(n_864), .B1(n_1350), .B2(n_1351), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_863), .A2(n_864), .B1(n_1387), .B2(n_1408), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_863), .A2(n_864), .B1(n_1574), .B2(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1319 ( .A(n_864), .Y(n_1319) );
INVx1_ASAP7_75t_L g885 ( .A(n_866), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_872), .Y(n_866) );
NAND2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_871), .Y(n_867) );
INVx2_ASAP7_75t_SL g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g1313 ( .A(n_870), .Y(n_1313) );
INVx1_ASAP7_75t_L g884 ( .A(n_873), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_874), .A2(n_877), .B1(n_958), .B2(n_976), .Y(n_975) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B(n_882), .Y(n_879) );
OAI21xp33_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_884), .B(n_885), .Y(n_883) );
INVx1_ASAP7_75t_L g943 ( .A(n_886), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_917), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g1436 ( .A1(n_898), .A2(n_1423), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
OAI211xp5_ASAP7_75t_L g930 ( .A1(n_901), .A2(n_931), .B(n_933), .C(n_934), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_904) );
OAI211xp5_ASAP7_75t_L g1308 ( .A1(n_905), .A2(n_1309), .B(n_1310), .C(n_1311), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1913 ( .A1(n_907), .A2(n_1914), .B1(n_1915), .B2(n_1916), .Y(n_1913) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_914), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_935), .C(n_939), .Y(n_917) );
NOR3xp33_ASAP7_75t_SL g918 ( .A(n_919), .B(n_927), .C(n_929), .Y(n_918) );
OAI21xp5_ASAP7_75t_SL g919 ( .A1(n_920), .A2(n_922), .B(n_923), .Y(n_919) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_948), .A2(n_973), .B(n_974), .Y(n_947) );
NAND4xp25_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .C(n_962), .D(n_967), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g1195 ( .A(n_951), .Y(n_1195) );
AOI222xp33_ASAP7_75t_L g1349 ( .A1(n_951), .A2(n_1197), .B1(n_1350), .B2(n_1351), .C1(n_1352), .C2(n_1354), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_960), .A2(n_969), .B1(n_1427), .B2(n_1431), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_960), .A2(n_1424), .B1(n_1438), .B2(n_1444), .Y(n_1447) );
INVx2_ASAP7_75t_L g1445 ( .A(n_961), .Y(n_1445) );
OAI211xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B(n_971), .C(n_972), .Y(n_967) );
INVx5_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_978), .A2(n_1253), .B1(n_1254), .B2(n_1255), .Y(n_1252) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_985), .A2(n_1307), .B1(n_1308), .B2(n_1312), .Y(n_1306) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_996), .B(n_1008), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_996), .B(n_1257), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_996), .B(n_1534), .Y(n_1566) );
INVx2_ASAP7_75t_L g1066 ( .A(n_997), .Y(n_1066) );
XOR2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1064), .Y(n_997) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_999), .B(n_1030), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1010), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1006), .Y(n_1002) );
NAND2xp5_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1009), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1171 ( .A(n_1009), .B(n_1172), .C(n_1174), .Y(n_1171) );
NAND4xp25_ASAP7_75t_L g1563 ( .A(n_1009), .B(n_1564), .C(n_1566), .D(n_1567), .Y(n_1563) );
AOI33xp33_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1012), .A3(n_1015), .B1(n_1018), .B2(n_1020), .B3(n_1021), .Y(n_1010) );
AOI33xp33_ASAP7_75t_L g1126 ( .A1(n_1011), .A2(n_1083), .A3(n_1127), .B1(n_1128), .B2(n_1131), .B3(n_1134), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1011), .B(n_1166), .Y(n_1165) );
AOI33xp33_ASAP7_75t_L g1209 ( .A1(n_1011), .A2(n_1210), .A3(n_1211), .B1(n_1212), .B2(n_1214), .B3(n_1215), .Y(n_1209) );
AOI33xp33_ASAP7_75t_L g1258 ( .A1(n_1011), .A2(n_1083), .A3(n_1259), .B1(n_1260), .B2(n_1262), .B3(n_1263), .Y(n_1258) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1020), .Y(n_1845) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1048), .B(n_1062), .Y(n_1030) );
NAND3xp33_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1035), .C(n_1047), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_1033), .A2(n_1234), .B1(n_1235), .B2(n_1236), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_1033), .A2(n_1275), .B1(n_1276), .B2(n_1277), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1929 ( .A1(n_1033), .A2(n_1276), .B1(n_1930), .B2(n_1931), .Y(n_1929) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1038), .Y(n_1184) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1038), .Y(n_1353) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1039), .Y(n_1109) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_SL g1045 ( .A(n_1046), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_1046), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_1051), .A2(n_1280), .B1(n_1281), .B2(n_1282), .C(n_1283), .Y(n_1279) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx4_ASAP7_75t_L g1856 ( .A(n_1052), .Y(n_1856) );
INVx4_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1057), .B1(n_1059), .B2(n_1060), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_1057), .A2(n_1060), .B1(n_1095), .B2(n_1096), .C(n_1097), .Y(n_1094) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1862 ( .A(n_1058), .Y(n_1862) );
OAI22xp33_ASAP7_75t_L g1853 ( .A1(n_1060), .A2(n_1828), .B1(n_1847), .B2(n_1854), .Y(n_1853) );
OAI22xp5_ASAP7_75t_L g1861 ( .A1(n_1060), .A2(n_1836), .B1(n_1844), .B2(n_1862), .Y(n_1861) );
INVx5_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
OAI21xp5_ASAP7_75t_SL g1384 ( .A1(n_1062), .A2(n_1385), .B(n_1392), .Y(n_1384) );
OAI21xp5_ASAP7_75t_L g1520 ( .A1(n_1062), .A2(n_1521), .B(n_1525), .Y(n_1520) );
OAI21xp5_ASAP7_75t_SL g1571 ( .A1(n_1062), .A2(n_1572), .B(n_1580), .Y(n_1571) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1063), .Y(n_1337) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1067), .Y(n_1151) );
XNOR2x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1114), .Y(n_1067) );
NAND3xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1088), .C(n_1091), .Y(n_1069) );
NOR3xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1085), .C(n_1087), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1075), .Y(n_1071) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1083), .Y(n_1435) );
NOR4xp25_ASAP7_75t_L g1900 ( .A(n_1087), .B(n_1901), .C(n_1903), .D(n_1904), .Y(n_1900) );
OAI21xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1101), .B(n_1113), .Y(n_1091) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1100), .Y(n_1229) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
AOI21xp5_ASAP7_75t_SL g1177 ( .A1(n_1113), .A2(n_1178), .B(n_1198), .Y(n_1177) );
O2A1O1Ixp5_ASAP7_75t_L g1265 ( .A1(n_1113), .A2(n_1266), .B(n_1278), .C(n_1287), .Y(n_1265) );
AND3x1_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1123), .C(n_1126), .Y(n_1119) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
OAI21xp5_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1144), .B(n_1150), .Y(n_1136) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g1607 ( .A(n_1153), .Y(n_1607) );
AOI22xp5_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1155), .B1(n_1293), .B2(n_1606), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
XNOR2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1249), .Y(n_1156) );
OAI22x1_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B1(n_1202), .B2(n_1248), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
XNOR2x1_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
AND3x2_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1177), .C(n_1200), .Y(n_1161) );
NOR2xp33_ASAP7_75t_SL g1162 ( .A(n_1163), .B(n_1171), .Y(n_1162) );
OAI21xp5_ASAP7_75t_SL g1163 ( .A1(n_1164), .A2(n_1165), .B(n_1168), .Y(n_1163) );
NAND3xp33_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1182), .C(n_1188), .Y(n_1178) );
AOI31xp33_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1190), .A3(n_1193), .B(n_1194), .Y(n_1188) );
INVx2_ASAP7_75t_SL g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1192), .Y(n_1325) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1192), .Y(n_1398) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1197), .B(n_1387), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_1197), .A2(n_1527), .B1(n_1528), .B2(n_1531), .Y(n_1526) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1197), .B(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1202), .Y(n_1248) );
NAND3xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1218), .C(n_1221), .Y(n_1203) );
NOR3xp33_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1216), .C(n_1217), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1209), .Y(n_1205) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1213), .Y(n_1430) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1213), .Y(n_1841) );
NOR3xp33_ASAP7_75t_L g1405 ( .A(n_1217), .B(n_1406), .C(n_1414), .Y(n_1405) );
OAI21xp5_ASAP7_75t_L g1221 ( .A1(n_1222), .A2(n_1238), .B(n_1246), .Y(n_1221) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1243), .Y(n_1239) );
OAI21xp5_ASAP7_75t_L g1920 ( .A1(n_1246), .A2(n_1921), .B(n_1924), .Y(n_1920) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
XOR2x2_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1292), .Y(n_1249) );
NAND3x1_ASAP7_75t_SL g1250 ( .A(n_1251), .B(n_1265), .C(n_1290), .Y(n_1250) );
INVx1_ASAP7_75t_L g1902 ( .A(n_1255), .Y(n_1902) );
HB1xp67_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1293), .Y(n_1606) );
AOI22xp5_ASAP7_75t_L g1293 ( .A1(n_1294), .A2(n_1295), .B1(n_1378), .B2(n_1379), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1340), .B1(n_1376), .B2(n_1377), .Y(n_1295) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1296), .Y(n_1376) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
NAND4xp75_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1305), .C(n_1320), .D(n_1338), .Y(n_1298) );
INVx1_ASAP7_75t_SL g1302 ( .A(n_1303), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g1826 ( .A1(n_1307), .A2(n_1827), .A3(n_1834), .B1(n_1840), .B2(n_1845), .B3(n_1846), .Y(n_1826) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1329), .B(n_1337), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1326), .Y(n_1321) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1332), .B1(n_1333), .B2(n_1335), .C(n_1336), .Y(n_1330) );
BUFx3_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AOI21xp5_ASAP7_75t_L g1347 ( .A1(n_1337), .A2(n_1348), .B(n_1362), .Y(n_1347) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1340), .Y(n_1377) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
NAND3xp33_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1347), .C(n_1364), .Y(n_1344) );
NAND3xp33_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1355), .C(n_1359), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1367), .Y(n_1365) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
AO22x2_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1515), .B1(n_1604), .B2(n_1605), .Y(n_1379) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1380), .Y(n_1604) );
XNOR2xp5_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1415), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
NAND3xp33_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1402), .C(n_1405), .Y(n_1383) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1409), .Y(n_1406) );
NAND3xp33_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1452), .C(n_1482), .Y(n_1416) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1439), .Y(n_1417) );
OAI33xp33_ASAP7_75t_L g1418 ( .A1(n_1419), .A2(n_1421), .A3(n_1426), .B1(n_1429), .B2(n_1435), .B3(n_1436), .Y(n_1418) );
BUFx3_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1421 ( .A1(n_1422), .A2(n_1423), .B1(n_1424), .B2(n_1425), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_1422), .A2(n_1437), .B1(n_1442), .B2(n_1444), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1431), .B1(n_1432), .B2(n_1434), .Y(n_1429) );
BUFx6f_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx2_ASAP7_75t_L g1492 ( .A(n_1433), .Y(n_1492) );
OAI33xp33_ASAP7_75t_L g1439 ( .A1(n_1440), .A2(n_1441), .A3(n_1446), .B1(n_1447), .B2(n_1448), .B3(n_1449), .Y(n_1439) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx2_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVx2_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
OAI31xp33_ASAP7_75t_SL g1452 ( .A1(n_1453), .A2(n_1465), .A3(n_1475), .B(n_1479), .Y(n_1452) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1455), .Y(n_1866) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1461), .B1(n_1462), .B2(n_1463), .Y(n_1457) );
BUFx3_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1867 ( .A1(n_1459), .A2(n_1868), .B1(n_1869), .B2(n_1870), .Y(n_1867) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_1461), .A2(n_1496), .B1(n_1500), .B2(n_1503), .Y(n_1495) );
BUFx3_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1871 ( .A(n_1464), .Y(n_1871) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
BUFx2_ASAP7_75t_L g1873 ( .A(n_1468), .Y(n_1873) );
INVx2_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx2_ASAP7_75t_L g1875 ( .A(n_1474), .Y(n_1875) );
INVx3_ASAP7_75t_SL g1477 ( .A(n_1478), .Y(n_1477) );
CKINVDCx16_ASAP7_75t_R g1877 ( .A(n_1478), .Y(n_1877) );
OAI31xp33_ASAP7_75t_SL g1863 ( .A1(n_1479), .A2(n_1864), .A3(n_1872), .B(n_1876), .Y(n_1863) );
BUFx3_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
OAI31xp33_ASAP7_75t_SL g1482 ( .A1(n_1483), .A2(n_1490), .A3(n_1504), .B(n_1510), .Y(n_1482) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx2_ASAP7_75t_L g1880 ( .A(n_1488), .Y(n_1880) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
CKINVDCx8_ASAP7_75t_R g1493 ( .A(n_1494), .Y(n_1493) );
CKINVDCx8_ASAP7_75t_R g1882 ( .A(n_1494), .Y(n_1882) );
BUFx3_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
AND2x4_ASAP7_75t_L g1501 ( .A(n_1498), .B(n_1502), .Y(n_1501) );
AND2x4_ASAP7_75t_L g1884 ( .A(n_1498), .B(n_1499), .Y(n_1884) );
BUFx6f_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
AOI22xp33_ASAP7_75t_SL g1883 ( .A1(n_1501), .A2(n_1868), .B1(n_1884), .B2(n_1885), .Y(n_1883) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVx2_ASAP7_75t_SL g1506 ( .A(n_1507), .Y(n_1506) );
BUFx3_ASAP7_75t_L g1887 ( .A(n_1507), .Y(n_1887) );
BUFx3_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1889 ( .A(n_1509), .Y(n_1889) );
OAI31xp33_ASAP7_75t_L g1878 ( .A1(n_1510), .A2(n_1879), .A3(n_1881), .B(n_1886), .Y(n_1878) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1513), .Y(n_1510) );
INVx1_ASAP7_75t_SL g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1515), .Y(n_1605) );
AOI22xp5_ASAP7_75t_L g1515 ( .A1(n_1516), .A2(n_1517), .B1(n_1569), .B2(n_1603), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NOR3xp33_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1563), .C(n_1568), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1537), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1524), .Y(n_1522) );
NAND3xp33_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1532), .C(n_1535), .Y(n_1525) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_1530), .Y(n_1529) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_1541), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1540) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OAI22xp33_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1549), .B1(n_1550), .B2(n_1551), .Y(n_1547) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx2_ASAP7_75t_L g1848 ( .A(n_1552), .Y(n_1848) );
OAI22xp5_ASAP7_75t_L g1557 ( .A1(n_1558), .A2(n_1559), .B1(n_1560), .B2(n_1562), .Y(n_1557) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1569), .Y(n_1603) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1570), .Y(n_1602) );
NAND3xp33_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1588), .C(n_1591), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1595), .Y(n_1592) );
OAI22xp5_ASAP7_75t_SL g1704 ( .A1(n_1601), .A2(n_1705), .B1(n_1706), .B2(n_1707), .Y(n_1704) );
OAI221xp5_ASAP7_75t_L g1608 ( .A1(n_1609), .A2(n_1818), .B1(n_1821), .B2(n_1890), .C(n_1893), .Y(n_1608) );
NOR3xp33_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1780), .C(n_1793), .Y(n_1609) );
NAND4xp25_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1708), .C(n_1730), .D(n_1763), .Y(n_1610) );
OAI31xp33_ASAP7_75t_L g1611 ( .A1(n_1612), .A2(n_1663), .A3(n_1693), .B(n_1702), .Y(n_1611) );
OAI21xp33_ASAP7_75t_L g1612 ( .A1(n_1613), .A2(n_1634), .B(n_1652), .Y(n_1612) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1614), .B(n_1728), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1614), .B(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1630), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1615), .B(n_1676), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1615), .B(n_1658), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1615), .B(n_1700), .Y(n_1699) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1615), .B(n_1630), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1615), .B(n_1702), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1615), .B(n_1667), .Y(n_1745) );
NAND3xp33_ASAP7_75t_L g1775 ( .A(n_1615), .B(n_1671), .C(n_1776), .Y(n_1775) );
CKINVDCx6p67_ASAP7_75t_R g1615 ( .A(n_1616), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1664 ( .A(n_1616), .B(n_1665), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1616), .B(n_1630), .Y(n_1715) );
OR2x2_ASAP7_75t_L g1724 ( .A(n_1616), .B(n_1630), .Y(n_1724) );
CKINVDCx5p33_ASAP7_75t_R g1749 ( .A(n_1616), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1616), .B(n_1703), .Y(n_1761) );
OR2x6_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1624), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1742 ( .A(n_1617), .B(n_1624), .Y(n_1742) );
INVx2_ASAP7_75t_L g1705 ( .A(n_1618), .Y(n_1705) );
AND2x6_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1620), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1619), .B(n_1623), .Y(n_1622) );
AND2x4_ASAP7_75t_L g1625 ( .A(n_1619), .B(n_1626), .Y(n_1625) );
AND2x6_ASAP7_75t_L g1628 ( .A(n_1619), .B(n_1629), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1619), .B(n_1623), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1619), .B(n_1623), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1820 ( .A(n_1619), .B(n_1626), .Y(n_1820) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1621), .B(n_1627), .Y(n_1626) );
HB1xp67_ASAP7_75t_L g1939 ( .A(n_1626), .Y(n_1939) );
OR2x2_ASAP7_75t_L g1659 ( .A(n_1630), .B(n_1660), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1630), .B(n_1667), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1630), .B(n_1660), .Y(n_1692) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1630), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1630), .B(n_1771), .Y(n_1770) );
INVx3_ASAP7_75t_L g1786 ( .A(n_1630), .Y(n_1786) );
OAI21xp5_ASAP7_75t_L g1796 ( .A1(n_1630), .A2(n_1711), .B(n_1797), .Y(n_1796) );
AND2x4_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1633), .Y(n_1630) );
INVxp67_ASAP7_75t_L g1707 ( .A(n_1632), .Y(n_1707) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1634), .Y(n_1791) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1640), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1635), .B(n_1641), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1635), .B(n_1690), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1635), .B(n_1653), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1635), .B(n_1654), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1635), .B(n_1766), .Y(n_1765) );
AND3x1_ASAP7_75t_L g1801 ( .A(n_1635), .B(n_1649), .C(n_1654), .Y(n_1801) );
INVx2_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
BUFx2_ASAP7_75t_L g1674 ( .A(n_1636), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1636), .B(n_1690), .Y(n_1697) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1636), .B(n_1755), .Y(n_1754) );
OR2x2_ASAP7_75t_L g1798 ( .A(n_1636), .B(n_1679), .Y(n_1798) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1636), .B(n_1645), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1640), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1645), .Y(n_1640) );
NOR2xp33_ASAP7_75t_L g1669 ( .A(n_1641), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1641), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1641), .B(n_1676), .Y(n_1685) );
NOR2xp33_ASAP7_75t_L g1752 ( .A(n_1641), .B(n_1753), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1641), .B(n_1684), .Y(n_1774) );
INVx2_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1642), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1642), .B(n_1645), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1642), .B(n_1674), .Y(n_1691) );
NOR2xp33_ASAP7_75t_L g1737 ( .A(n_1642), .B(n_1738), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1762 ( .A(n_1642), .B(n_1667), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1642), .B(n_1660), .Y(n_1771) );
OR2x2_ASAP7_75t_L g1777 ( .A(n_1642), .B(n_1660), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .Y(n_1642) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1645), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1649), .Y(n_1645) );
INVx2_ASAP7_75t_L g1654 ( .A(n_1646), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1646), .B(n_1655), .Y(n_1690) );
OR2x2_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1648), .Y(n_1646) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1649), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1649), .B(n_1654), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1649), .B(n_1674), .Y(n_1684) );
OR2x2_ASAP7_75t_L g1753 ( .A(n_1649), .B(n_1674), .Y(n_1753) );
AOI32xp33_ASAP7_75t_L g1769 ( .A1(n_1649), .A2(n_1749), .A3(n_1770), .B1(n_1772), .B2(n_1773), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1651), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1656), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1653), .B(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1653), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1653), .B(n_1657), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1655), .Y(n_1653) );
OR2x2_ASAP7_75t_L g1738 ( .A(n_1654), .B(n_1674), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1654), .B(n_1674), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1655), .B(n_1674), .Y(n_1673) );
OAI211xp5_ASAP7_75t_L g1739 ( .A1(n_1656), .A2(n_1740), .B(n_1741), .C(n_1742), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1658), .Y(n_1656) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1657), .Y(n_1696) );
INVx2_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
AOI211xp5_ASAP7_75t_L g1757 ( .A1(n_1659), .A2(n_1696), .B(n_1749), .C(n_1758), .Y(n_1757) );
OAI22xp5_ASAP7_75t_L g1781 ( .A1(n_1659), .A2(n_1782), .B1(n_1786), .B2(n_1787), .Y(n_1781) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1660), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1660), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1662), .Y(n_1660) );
OAI211xp5_ASAP7_75t_SL g1663 ( .A1(n_1664), .A2(n_1668), .B(n_1672), .C(n_1686), .Y(n_1663) );
OAI21xp5_ASAP7_75t_L g1693 ( .A1(n_1665), .A2(n_1694), .B(n_1698), .Y(n_1693) );
A2O1A1Ixp33_ASAP7_75t_L g1802 ( .A1(n_1665), .A2(n_1778), .B(n_1803), .C(n_1804), .Y(n_1802) );
CKINVDCx6p67_ASAP7_75t_R g1665 ( .A(n_1666), .Y(n_1665) );
AOI31xp33_ASAP7_75t_L g1746 ( .A1(n_1666), .A2(n_1691), .A3(n_1747), .B(n_1749), .Y(n_1746) );
INVx2_ASAP7_75t_L g1676 ( .A(n_1667), .Y(n_1676) );
OAI211xp5_ASAP7_75t_SL g1768 ( .A1(n_1668), .A2(n_1723), .B(n_1769), .C(n_1775), .Y(n_1768) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
AOI211xp5_ASAP7_75t_L g1759 ( .A1(n_1670), .A2(n_1760), .B(n_1761), .C(n_1762), .Y(n_1759) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1726 ( .A(n_1671), .B(n_1688), .Y(n_1726) );
OR2x2_ASAP7_75t_L g1748 ( .A(n_1671), .B(n_1690), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1812 ( .A(n_1671), .B(n_1674), .Y(n_1812) );
AOI321xp33_ASAP7_75t_L g1672 ( .A1(n_1673), .A2(n_1675), .A3(n_1677), .B1(n_1678), .B2(n_1680), .C(n_1682), .Y(n_1672) );
AOI221xp5_ASAP7_75t_L g1743 ( .A1(n_1675), .A2(n_1725), .B1(n_1744), .B2(n_1745), .C(n_1746), .Y(n_1743) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1675), .Y(n_1767) );
INVx2_ASAP7_75t_L g1712 ( .A(n_1676), .Y(n_1712) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AOI21xp33_ASAP7_75t_SL g1764 ( .A1(n_1679), .A2(n_1765), .B(n_1767), .Y(n_1764) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
NOR2xp33_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1685), .Y(n_1682) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
OAI21xp33_ASAP7_75t_L g1686 ( .A1(n_1687), .A2(n_1689), .B(n_1692), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1687), .B(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1687), .Y(n_1744) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1689), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1691), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1690), .B(n_1699), .Y(n_1698) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1691), .Y(n_1721) );
INVx2_ASAP7_75t_L g1792 ( .A(n_1692), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1697), .Y(n_1694) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1696), .B(n_1714), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1696), .B(n_1733), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1696), .B(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1697), .Y(n_1758) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1699), .Y(n_1756) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1700), .Y(n_1790) );
AOI211xp5_ASAP7_75t_L g1806 ( .A1(n_1700), .A2(n_1709), .B(n_1807), .C(n_1808), .Y(n_1806) );
OAI32xp33_ASAP7_75t_L g1813 ( .A1(n_1701), .A2(n_1778), .A3(n_1814), .B1(n_1815), .B2(n_1816), .Y(n_1813) );
OAI321xp33_ASAP7_75t_L g1731 ( .A1(n_1702), .A2(n_1711), .A3(n_1732), .B1(n_1734), .B2(n_1735), .C(n_1739), .Y(n_1731) );
INVx2_ASAP7_75t_SL g1702 ( .A(n_1703), .Y(n_1702) );
INVx2_ASAP7_75t_SL g1779 ( .A(n_1703), .Y(n_1779) );
O2A1O1Ixp33_ASAP7_75t_L g1708 ( .A1(n_1709), .A2(n_1713), .B(n_1715), .C(n_1716), .Y(n_1708) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1711), .B(n_1719), .Y(n_1718) );
A2O1A1Ixp33_ASAP7_75t_L g1794 ( .A1(n_1711), .A2(n_1737), .B(n_1786), .C(n_1795), .Y(n_1794) );
INVx2_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1712), .B(n_1729), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1783 ( .A(n_1712), .B(n_1784), .Y(n_1783) );
NAND2xp5_ASAP7_75t_L g1788 ( .A(n_1712), .B(n_1713), .Y(n_1788) );
AOI21xp33_ASAP7_75t_SL g1799 ( .A1(n_1712), .A2(n_1800), .B(n_1802), .Y(n_1799) );
OAI221xp5_ASAP7_75t_L g1716 ( .A1(n_1717), .A2(n_1723), .B1(n_1724), .B2(n_1725), .C(n_1727), .Y(n_1716) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
OR2x2_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1722), .Y(n_1720) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1724), .Y(n_1772) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
NOR5xp2_ASAP7_75t_SL g1730 ( .A(n_1731), .B(n_1743), .C(n_1750), .D(n_1757), .E(n_1759), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1732), .B(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1734), .Y(n_1817) );
INVxp67_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1738), .Y(n_1741) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
AOI21xp33_ASAP7_75t_SL g1750 ( .A1(n_1751), .A2(n_1754), .B(n_1756), .Y(n_1750) );
INVxp33_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1754), .Y(n_1814) );
O2A1O1Ixp33_ASAP7_75t_L g1780 ( .A1(n_1758), .A2(n_1761), .B(n_1781), .C(n_1789), .Y(n_1780) );
OAI211xp5_ASAP7_75t_L g1795 ( .A1(n_1758), .A2(n_1777), .B(n_1785), .C(n_1796), .Y(n_1795) );
OAI21xp5_ASAP7_75t_L g1763 ( .A1(n_1764), .A2(n_1768), .B(n_1778), .Y(n_1763) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1766), .Y(n_1805) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx3_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NAND2xp5_ASAP7_75t_L g1816 ( .A(n_1779), .B(n_1786), .Y(n_1816) );
INVxp67_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
AOI221xp5_ASAP7_75t_L g1793 ( .A1(n_1788), .A2(n_1794), .B1(n_1799), .B2(n_1806), .C(n_1817), .Y(n_1793) );
OAI21xp5_ASAP7_75t_SL g1789 ( .A1(n_1790), .A2(n_1791), .B(n_1792), .Y(n_1789) );
OAI21xp5_ASAP7_75t_SL g1808 ( .A1(n_1792), .A2(n_1809), .B(n_1813), .Y(n_1808) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVx2_ASAP7_75t_L g1803 ( .A(n_1801), .Y(n_1803) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
CKINVDCx20_ASAP7_75t_R g1818 ( .A(n_1819), .Y(n_1818) );
CKINVDCx5p33_ASAP7_75t_R g1819 ( .A(n_1820), .Y(n_1819) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
NAND3xp33_ASAP7_75t_L g1824 ( .A(n_1825), .B(n_1863), .C(n_1878), .Y(n_1824) );
NOR2xp33_ASAP7_75t_L g1825 ( .A(n_1826), .B(n_1850), .Y(n_1825) );
OAI22xp33_ASAP7_75t_L g1827 ( .A1(n_1828), .A2(n_1829), .B1(n_1831), .B2(n_1832), .Y(n_1827) );
OAI22xp33_ASAP7_75t_L g1846 ( .A1(n_1829), .A2(n_1847), .B1(n_1848), .B2(n_1849), .Y(n_1846) );
BUFx4f_ASAP7_75t_SL g1829 ( .A(n_1830), .Y(n_1829) );
OAI22xp5_ASAP7_75t_L g1858 ( .A1(n_1831), .A2(n_1849), .B1(n_1856), .B2(n_1859), .Y(n_1858) );
INVxp67_ASAP7_75t_SL g1832 ( .A(n_1833), .Y(n_1832) );
OAI22xp33_ASAP7_75t_L g1855 ( .A1(n_1835), .A2(n_1842), .B1(n_1856), .B2(n_1857), .Y(n_1855) );
INVx3_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
BUFx2_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
OAI22xp5_ASAP7_75t_L g1840 ( .A1(n_1841), .A2(n_1842), .B1(n_1843), .B2(n_1844), .Y(n_1840) );
OAI33xp33_ASAP7_75t_L g1850 ( .A1(n_1851), .A2(n_1853), .A3(n_1855), .B1(n_1858), .B2(n_1860), .B3(n_1861), .Y(n_1850) );
BUFx6f_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx2_ASAP7_75t_L g1870 ( .A(n_1871), .Y(n_1870) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1875), .Y(n_1874) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
INVx3_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
HB1xp67_ASAP7_75t_L g1894 ( .A(n_1895), .Y(n_1894) );
BUFx3_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
INVxp33_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
AND3x2_ASAP7_75t_L g1899 ( .A(n_1900), .B(n_1920), .C(n_1932), .Y(n_1899) );
INVx1_ASAP7_75t_L g1909 ( .A(n_1910), .Y(n_1909) );
HB1xp67_ASAP7_75t_L g1935 ( .A(n_1936), .Y(n_1935) );
HB1xp67_ASAP7_75t_L g1936 ( .A(n_1937), .Y(n_1936) );
OAI21xp5_ASAP7_75t_L g1937 ( .A1(n_1938), .A2(n_1939), .B(n_1940), .Y(n_1937) );
INVx1_ASAP7_75t_L g1940 ( .A(n_1941), .Y(n_1940) );
endmodule