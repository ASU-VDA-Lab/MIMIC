module real_jpeg_23621_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_292;
wire n_288;
wire n_221;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_216;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_295;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_47),
.B1(n_72),
.B2(n_73),
.Y(n_125)
);

INVx8_ASAP7_75t_SL g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_88),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_162),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_26),
.B(n_42),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_119),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_23),
.B1(n_241),
.B2(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_72),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_77),
.B1(n_80),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_6),
.A2(n_72),
.B1(n_73),
.B2(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_170),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_170),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_51),
.B1(n_72),
.B2(n_73),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_51),
.B1(n_77),
.B2(n_113),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_72),
.B1(n_73),
.B2(n_83),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_83),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_83),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_11),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_72),
.B1(n_73),
.B2(n_114),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_114),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_114),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_64),
.B1(n_72),
.B2(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_33),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_33),
.B1(n_72),
.B2(n_73),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_128)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_20),
.B(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_20),
.B(n_148),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_53),
.CI(n_99),
.CON(n_20),
.SN(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_22),
.B(n_35),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_22),
.A2(n_52),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_31),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_23),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_23),
.A2(n_59),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_23),
.A2(n_61),
.B1(n_233),
.B2(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_23),
.A2(n_31),
.B(n_105),
.Y(n_269)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_24),
.B(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_24),
.A2(n_60),
.B1(n_104),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_24),
.A2(n_106),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_25),
.B(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_29),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_29),
.A2(n_57),
.B(n_167),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_46),
.B(n_48),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_45),
.B1(n_46),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_36),
.A2(n_45),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_36),
.A2(n_127),
.B(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_37),
.A2(n_49),
.B(n_128),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_37),
.A2(n_129),
.B1(n_217),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_37),
.A2(n_129),
.B1(n_225),
.B2(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_45),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_40),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_39),
.B(n_92),
.Y(n_268)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_40),
.A2(n_44),
.B(n_162),
.C(n_219),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_40),
.A2(n_72),
.A3(n_91),
.B1(n_261),
.B2(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_45),
.A2(n_63),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_45),
.B(n_162),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_50),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_98),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_54),
.B(n_66),
.C(n_89),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_56),
.B(n_62),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_89),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_81),
.B(n_84),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_68),
.B1(n_81),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_76),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_70),
.B1(n_77),
.B2(n_80),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_69),
.A2(n_73),
.A3(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_159)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_70),
.B(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_73),
.B1(n_91),
.B2(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_73),
.B(n_162),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_80),
.A2(n_161),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_85),
.Y(n_137)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_88),
.B(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_88),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_88),
.A2(n_169),
.B1(n_171),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_117),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_90),
.A2(n_116),
.B1(n_201),
.B2(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_95),
.A2(n_119),
.B1(n_156),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_95),
.A2(n_119),
.B1(n_186),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.C(n_115),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_101),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_107),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_115),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_143),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_131),
.B1(n_141),
.B2(n_142),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B(n_130),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_140),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_173),
.B(n_296),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_149),
.B(n_177),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.CI(n_154),
.CON(n_149),
.SN(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_168),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_168),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_164),
.B1(n_165),
.B2(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_162),
.B(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_206),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_188),
.B(n_205),
.Y(n_175)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_187),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_179),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_187),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.C(n_185),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_185),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_189),
.B(n_192),
.Y(n_295)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_195),
.Y(n_292)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_199),
.B(n_278),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_202),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_294),
.C(n_295),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_288),
.B(n_293),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_273),
.B(n_287),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_254),
.B(n_272),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_229),
.B(n_253),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_226),
.C(n_227),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_237),
.B(n_252),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_235),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_251),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_265),
.C(n_270),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_283),
.C(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);


endmodule