module real_aes_7151_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_1), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_1), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_2), .A2(n_132), .B(n_137), .C(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_3), .A2(n_127), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_4), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g487 ( .A(n_5), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_6), .B(n_165), .Y(n_231) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_7), .A2(n_127), .B(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_L g132 ( .A(n_8), .B(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_9), .A2(n_262), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g144 ( .A(n_10), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_11), .B(n_43), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_12), .B(n_142), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_13), .B(n_189), .Y(n_466) );
INVx1_ASAP7_75t_L g500 ( .A(n_14), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_15), .A2(n_33), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_15), .Y(n_734) );
INVx1_ASAP7_75t_L g125 ( .A(n_16), .Y(n_125) );
INVx1_ASAP7_75t_L g478 ( .A(n_17), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_18), .A2(n_145), .B(n_159), .C(n_163), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_19), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_20), .B(n_457), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_21), .B(n_127), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_22), .B(n_271), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_23), .A2(n_189), .B(n_190), .C(n_192), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_24), .B(n_165), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_25), .B(n_142), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_26), .A2(n_161), .B(n_163), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_27), .B(n_142), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
INVx1_ASAP7_75t_L g201 ( .A(n_29), .Y(n_201) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_30), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_31), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_32), .B(n_142), .Y(n_488) );
INVx1_ASAP7_75t_L g733 ( .A(n_33), .Y(n_733) );
INVx1_ASAP7_75t_L g267 ( .A(n_34), .Y(n_267) );
INVx1_ASAP7_75t_L g508 ( .A(n_35), .Y(n_508) );
INVx2_ASAP7_75t_L g130 ( .A(n_36), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_37), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_38), .A2(n_189), .B(n_227), .C(n_229), .Y(n_226) );
INVxp67_ASAP7_75t_L g268 ( .A(n_39), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_40), .A2(n_137), .B(n_200), .C(n_206), .Y(n_199) );
CKINVDCx14_ASAP7_75t_R g225 ( .A(n_41), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_42), .A2(n_132), .B(n_137), .C(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g507 ( .A(n_44), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_45), .A2(n_141), .B(n_143), .C(n_146), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_46), .B(n_142), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_47), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_48), .Y(n_264) );
INVx1_ASAP7_75t_L g187 ( .A(n_49), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_50), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_51), .B(n_127), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_52), .A2(n_137), .B1(n_192), .B2(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_53), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_54), .Y(n_484) );
CKINVDCx14_ASAP7_75t_R g135 ( .A(n_55), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_56), .A2(n_141), .B(n_229), .C(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_57), .Y(n_545) );
INVx1_ASAP7_75t_L g497 ( .A(n_58), .Y(n_497) );
INVx1_ASAP7_75t_L g133 ( .A(n_59), .Y(n_133) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
INVx1_ASAP7_75t_SL g228 ( .A(n_61), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_62), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_63), .B(n_165), .Y(n_194) );
INVx1_ASAP7_75t_L g216 ( .A(n_64), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_SL g516 ( .A1(n_65), .A2(n_229), .B(n_457), .C(n_517), .Y(n_516) );
INVxp67_ASAP7_75t_L g518 ( .A(n_66), .Y(n_518) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_67), .A2(n_444), .B1(n_729), .B2(n_735), .C1(n_736), .C2(n_740), .Y(n_443) );
INVx1_ASAP7_75t_L g441 ( .A(n_68), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_69), .A2(n_127), .B(n_134), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_70), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_71), .A2(n_127), .B(n_156), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_72), .Y(n_511) );
INVx1_ASAP7_75t_L g539 ( .A(n_73), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_74), .A2(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g157 ( .A(n_75), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_76), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g427 ( .A1(n_77), .A2(n_78), .B1(n_428), .B2(n_429), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_77), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_78), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_79), .A2(n_132), .B(n_137), .C(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_80), .A2(n_127), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g160 ( .A(n_81), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_82), .B(n_202), .Y(n_455) );
INVx2_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
INVx1_ASAP7_75t_L g176 ( .A(n_84), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_85), .B(n_457), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_86), .A2(n_132), .B(n_137), .C(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g726 ( .A(n_87), .Y(n_726) );
OR2x2_ASAP7_75t_L g728 ( .A(n_87), .B(n_109), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_88), .A2(n_137), .B(n_215), .C(n_218), .Y(n_214) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_89), .A2(n_103), .B1(n_433), .B2(n_442), .C1(n_741), .C2(n_745), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_89), .A2(n_113), .B1(n_114), .B2(n_430), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_89), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_90), .B(n_121), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_91), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_92), .A2(n_132), .B(n_137), .C(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_93), .Y(n_470) );
INVx1_ASAP7_75t_L g515 ( .A(n_94), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_95), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_96), .B(n_202), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_97), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_98), .B(n_150), .Y(n_479) );
INVx2_ASAP7_75t_L g191 ( .A(n_99), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_100), .B(n_441), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_101), .A2(n_127), .B(n_514), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_112), .B(n_431), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g432 ( .A(n_107), .Y(n_432) );
BUFx2_ASAP7_75t_L g747 ( .A(n_107), .Y(n_747) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_108), .B(n_726), .Y(n_735) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g725 ( .A(n_109), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
XOR2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_427), .Y(n_114) );
INVx2_ASAP7_75t_L g727 ( .A(n_115), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_115), .A2(n_728), .B1(n_737), .B2(n_738), .Y(n_736) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_357), .Y(n_115) );
NAND5xp2_ASAP7_75t_L g116 ( .A(n_117), .B(n_272), .C(n_304), .D(n_321), .E(n_344), .Y(n_116) );
AOI221xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_195), .B1(n_232), .B2(n_236), .C(n_240), .Y(n_117) );
INVx1_ASAP7_75t_L g384 ( .A(n_118), .Y(n_384) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_167), .Y(n_118) );
AND3x2_ASAP7_75t_L g359 ( .A(n_119), .B(n_169), .C(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_152), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_120), .B(n_238), .Y(n_237) );
BUFx3_ASAP7_75t_L g247 ( .A(n_120), .Y(n_247) );
AND2x2_ASAP7_75t_L g251 ( .A(n_120), .B(n_183), .Y(n_251) );
INVx2_ASAP7_75t_L g281 ( .A(n_120), .Y(n_281) );
OR2x2_ASAP7_75t_L g292 ( .A(n_120), .B(n_184), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_120), .B(n_168), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_120), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g371 ( .A(n_120), .B(n_184), .Y(n_371) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_126), .B(n_149), .Y(n_120) );
INVx1_ASAP7_75t_L g170 ( .A(n_121), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_121), .A2(n_173), .B(n_198), .C(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g221 ( .A(n_121), .Y(n_221) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_121), .A2(n_473), .B(n_479), .Y(n_472) );
AND2x2_ASAP7_75t_SL g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_L g151 ( .A(n_122), .B(n_123), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
BUFx2_ASAP7_75t_L g262 ( .A(n_127), .Y(n_262) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_128), .B(n_132), .Y(n_173) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g205 ( .A(n_129), .Y(n_205) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
INVx1_ASAP7_75t_L g193 ( .A(n_130), .Y(n_193) );
INVx1_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
INVx3_ASAP7_75t_L g145 ( .A(n_131), .Y(n_145) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
INVx1_ASAP7_75t_L g457 ( .A(n_131), .Y(n_457) );
INVx4_ASAP7_75t_SL g148 ( .A(n_132), .Y(n_148) );
BUFx3_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_136), .B(n_140), .C(n_148), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_136), .A2(n_148), .B(n_157), .C(n_158), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g186 ( .A1(n_136), .A2(n_148), .B(n_187), .C(n_188), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_136), .A2(n_148), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_136), .A2(n_148), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_136), .A2(n_148), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_136), .A2(n_148), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_136), .A2(n_148), .B(n_515), .C(n_516), .Y(n_514) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx3_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_138), .Y(n_230) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx5_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_145), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_145), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_148), .A2(n_173), .B1(n_505), .B2(n_509), .Y(n_504) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_150), .Y(n_154) );
INVx4_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_150), .A2(n_513), .B(n_519), .Y(n_512) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g259 ( .A(n_151), .Y(n_259) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_152), .Y(n_250) );
AND2x2_ASAP7_75t_L g312 ( .A(n_152), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_152), .B(n_168), .Y(n_331) );
INVx1_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g239 ( .A(n_153), .B(n_168), .Y(n_239) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_153), .Y(n_246) );
AND2x2_ASAP7_75t_L g298 ( .A(n_153), .B(n_184), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_153), .B(n_167), .C(n_281), .Y(n_323) );
AND2x2_ASAP7_75t_L g388 ( .A(n_153), .B(n_169), .Y(n_388) );
AND2x2_ASAP7_75t_L g422 ( .A(n_153), .B(n_168), .Y(n_422) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_164), .Y(n_153) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_154), .A2(n_185), .B(n_194), .Y(n_184) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_154), .A2(n_223), .B(n_231), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_161), .B(n_191), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_161), .A2(n_202), .B1(n_267), .B2(n_268), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_161), .B(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g178 ( .A(n_162), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g506 ( .A1(n_162), .A2(n_178), .B1(n_507), .B2(n_508), .Y(n_506) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_165), .A2(n_495), .B(n_501), .Y(n_494) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_166), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_166), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_212), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_166), .B(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_L g248 ( .A(n_167), .Y(n_248) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_168), .B(n_281), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_168), .B(n_312), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_168), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g398 ( .A(n_168), .Y(n_398) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g305 ( .A(n_169), .B(n_298), .Y(n_305) );
BUFx3_ASAP7_75t_L g337 ( .A(n_169), .Y(n_337) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_181), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_170), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_170), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_170), .B(n_545), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_173), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_173), .A2(n_484), .B(n_485), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_173), .A2(n_539), .B(n_540), .Y(n_538) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .C(n_180), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_177), .A2(n_180), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_180), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_180), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g313 ( .A(n_183), .Y(n_313) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_189), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g489 ( .A(n_192), .Y(n_489) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_195), .A2(n_373), .B1(n_375), .B2(n_376), .Y(n_372) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_209), .Y(n_195) );
AND2x2_ASAP7_75t_L g232 ( .A(n_196), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_SL g243 ( .A(n_196), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_196), .B(n_276), .Y(n_308) );
OR2x2_ASAP7_75t_L g327 ( .A(n_196), .B(n_210), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_196), .B(n_284), .Y(n_332) );
AND2x2_ASAP7_75t_L g335 ( .A(n_196), .B(n_277), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_196), .B(n_222), .Y(n_347) );
AND2x2_ASAP7_75t_L g363 ( .A(n_196), .B(n_211), .Y(n_363) );
AND2x4_ASAP7_75t_L g366 ( .A(n_196), .B(n_234), .Y(n_366) );
OR2x2_ASAP7_75t_L g383 ( .A(n_196), .B(n_319), .Y(n_383) );
OR2x2_ASAP7_75t_L g414 ( .A(n_196), .B(n_256), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_196), .B(n_342), .Y(n_416) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_204), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_202), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_205), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g290 ( .A(n_209), .B(n_254), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_209), .B(n_277), .Y(n_409) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_222), .Y(n_209) );
AND2x2_ASAP7_75t_L g242 ( .A(n_210), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g276 ( .A(n_210), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g284 ( .A(n_210), .B(n_256), .Y(n_284) );
AND2x2_ASAP7_75t_L g302 ( .A(n_210), .B(n_234), .Y(n_302) );
OR2x2_ASAP7_75t_L g319 ( .A(n_210), .B(n_277), .Y(n_319) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
AND2x2_ASAP7_75t_L g342 ( .A(n_211), .B(n_222), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_221), .A2(n_462), .B(n_469), .Y(n_461) );
INVx2_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
INVx1_ASAP7_75t_L g354 ( .A(n_222), .Y(n_354) );
AND2x2_ASAP7_75t_L g404 ( .A(n_222), .B(n_243), .Y(n_404) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_230), .Y(n_467) );
AND2x2_ASAP7_75t_L g253 ( .A(n_233), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g288 ( .A(n_233), .B(n_243), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_233), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x2_ASAP7_75t_L g275 ( .A(n_234), .B(n_243), .Y(n_275) );
OR2x2_ASAP7_75t_L g391 ( .A(n_235), .B(n_365), .Y(n_391) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_238), .B(n_371), .Y(n_377) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OAI32xp33_ASAP7_75t_L g333 ( .A1(n_239), .A2(n_334), .A3(n_336), .B1(n_338), .B2(n_339), .Y(n_333) );
OR2x2_ASAP7_75t_L g350 ( .A(n_239), .B(n_292), .Y(n_350) );
OAI21xp33_ASAP7_75t_SL g375 ( .A1(n_239), .A2(n_249), .B(n_280), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B1(n_249), .B2(n_252), .Y(n_240) );
INVxp33_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_242), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_243), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g301 ( .A(n_243), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g401 ( .A(n_243), .B(n_342), .Y(n_401) );
OR2x2_ASAP7_75t_L g425 ( .A(n_243), .B(n_319), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_244), .A2(n_307), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g285 ( .A(n_246), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_246), .B(n_251), .Y(n_303) );
AND2x2_ASAP7_75t_L g325 ( .A(n_247), .B(n_298), .Y(n_325) );
INVx1_ASAP7_75t_L g338 ( .A(n_247), .Y(n_338) );
OR2x2_ASAP7_75t_L g343 ( .A(n_247), .B(n_277), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_250), .B(n_292), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_274), .B1(n_279), .B2(n_283), .Y(n_273) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_254), .A2(n_316), .B1(n_323), .B2(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g400 ( .A(n_254), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_256), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g419 ( .A(n_256), .B(n_302), .Y(n_419) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B(n_269), .Y(n_256) );
INVx1_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_257), .A2(n_538), .B(n_544), .Y(n_537) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AOI21xp5_ASAP7_75t_SL g451 ( .A1(n_258), .A2(n_452), .B(n_453), .Y(n_451) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_259), .A2(n_483), .B(n_490), .Y(n_482) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_259), .A2(n_504), .B(n_510), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_259), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_261), .A2(n_270), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_285), .B1(n_286), .B2(n_291), .C(n_293), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_275), .B(n_277), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_275), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_276), .A2(n_382), .B(n_383), .C(n_384), .Y(n_381) );
AND2x2_ASAP7_75t_L g386 ( .A(n_276), .B(n_366), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_SL g424 ( .A1(n_276), .A2(n_365), .B(n_425), .C(n_426), .Y(n_424) );
BUFx3_ASAP7_75t_L g316 ( .A(n_277), .Y(n_316) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_280), .B(n_337), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_280), .A2(n_400), .B(n_402), .C(n_408), .Y(n_399) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVxp67_ASAP7_75t_L g360 ( .A(n_282), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_284), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AOI211xp5_ASAP7_75t_L g304 ( .A1(n_288), .A2(n_305), .B(n_306), .C(n_314), .Y(n_304) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g389 ( .A(n_292), .Y(n_389) );
OR2x2_ASAP7_75t_L g406 ( .A(n_292), .B(n_336), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B1(n_300), .B2(n_303), .Y(n_293) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_295), .A2(n_307), .B1(n_308), .B2(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OR2x2_ASAP7_75t_L g393 ( .A(n_297), .B(n_337), .Y(n_393) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g348 ( .A(n_298), .B(n_338), .Y(n_348) );
INVx1_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_302), .B(n_316), .Y(n_364) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_312), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g421 ( .A(n_313), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_320), .Y(n_314) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_316), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_316), .B(n_347), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_316), .B(n_342), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_316), .B(n_363), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_316), .A2(n_326), .B(n_366), .C(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_326), .B1(n_328), .B2(n_332), .C(n_333), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_330), .B(n_338), .Y(n_412) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g423 ( .A1(n_332), .A2(n_347), .B(n_349), .C(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_335), .B(n_342), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_336), .B(n_389), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g336 ( .A(n_337), .Y(n_336) );
INVxp33_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AOI21xp33_ASAP7_75t_SL g352 ( .A1(n_341), .A2(n_353), .B(n_355), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_341), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_342), .B(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B1(n_349), .B2(n_351), .C(n_352), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_348), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
NAND5xp2_ASAP7_75t_L g357 ( .A(n_358), .B(n_385), .C(n_399), .D(n_410), .E(n_423), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_368), .C(n_381), .Y(n_358) );
INVx2_ASAP7_75t_SL g405 ( .A(n_359), .Y(n_405) );
NAND4xp25_ASAP7_75t_SL g361 ( .A(n_362), .B(n_364), .C(n_365), .D(n_367), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_367), .A2(n_369), .B(n_372), .C(n_378), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_411), .B1(n_413), .B2(n_415), .C(n_417), .Y(n_410) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .B1(n_390), .B2(n_392), .C(n_394), .Y(n_385) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_406), .B2(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_SL g744 ( .A(n_432), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
CKINVDCx6p67_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_SL g743 ( .A(n_438), .B(n_440), .Y(n_743) );
OA21x2_ASAP7_75t_L g746 ( .A1(n_438), .A2(n_439), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_444) );
INVx2_ASAP7_75t_L g737 ( .A(n_445), .Y(n_737) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_694), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_587), .C(n_660), .Y(n_446) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_480), .B(n_520), .C(n_571), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_460), .Y(n_449) );
AND2x2_ASAP7_75t_L g536 ( .A(n_450), .B(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g554 ( .A(n_450), .Y(n_554) );
INVx2_ASAP7_75t_L g569 ( .A(n_450), .Y(n_569) );
INVx1_ASAP7_75t_L g599 ( .A(n_450), .Y(n_599) );
AND2x2_ASAP7_75t_L g649 ( .A(n_450), .B(n_570), .Y(n_649) );
AOI32xp33_ASAP7_75t_L g676 ( .A1(n_450), .A2(n_604), .A3(n_677), .B1(n_679), .B2(n_680), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_450), .B(n_526), .Y(n_682) );
AND2x2_ASAP7_75t_L g709 ( .A(n_450), .B(n_552), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_450), .B(n_718), .Y(n_717) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .Y(n_450) );
AND2x2_ASAP7_75t_L g598 ( .A(n_460), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g620 ( .A(n_460), .Y(n_620) );
AND2x2_ASAP7_75t_L g705 ( .A(n_460), .B(n_536), .Y(n_705) );
AND2x2_ASAP7_75t_L g708 ( .A(n_460), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_471), .Y(n_460) );
INVx2_ASAP7_75t_L g528 ( .A(n_461), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_461), .B(n_552), .Y(n_558) );
AND2x2_ASAP7_75t_L g568 ( .A(n_461), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g604 ( .A(n_461), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_468), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_467), .Y(n_464) );
AND2x2_ASAP7_75t_L g546 ( .A(n_471), .B(n_528), .Y(n_546) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g529 ( .A(n_472), .Y(n_529) );
AND2x2_ASAP7_75t_L g570 ( .A(n_472), .B(n_552), .Y(n_570) );
AND2x2_ASAP7_75t_L g639 ( .A(n_472), .B(n_537), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
OR2x2_ASAP7_75t_L g534 ( .A(n_481), .B(n_503), .Y(n_534) );
INVx1_ASAP7_75t_L g612 ( .A(n_481), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_481), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_481), .B(n_502), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_481), .B(n_624), .Y(n_678) );
AND2x2_ASAP7_75t_L g686 ( .A(n_481), .B(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g524 ( .A(n_482), .Y(n_524) );
AND2x2_ASAP7_75t_L g593 ( .A(n_482), .B(n_503), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_492), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g720 ( .A(n_492), .Y(n_720) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_493), .B(n_564), .Y(n_586) );
OR2x2_ASAP7_75t_L g615 ( .A(n_493), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g647 ( .A(n_493), .B(n_627), .Y(n_647) );
INVx1_ASAP7_75t_SL g667 ( .A(n_493), .Y(n_667) );
AND2x2_ASAP7_75t_L g671 ( .A(n_493), .B(n_533), .Y(n_671) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_SL g525 ( .A(n_494), .B(n_502), .Y(n_525) );
AND2x2_ASAP7_75t_L g532 ( .A(n_494), .B(n_512), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_494), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_556), .Y(n_574) );
INVx1_ASAP7_75t_SL g581 ( .A(n_494), .Y(n_581) );
BUFx2_ASAP7_75t_L g592 ( .A(n_494), .Y(n_592) );
AND2x2_ASAP7_75t_L g608 ( .A(n_494), .B(n_524), .Y(n_608) );
AND2x2_ASAP7_75t_L g623 ( .A(n_494), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g687 ( .A(n_494), .B(n_503), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_502), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g611 ( .A(n_502), .B(n_612), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_502), .A2(n_629), .B1(n_632), .B2(n_635), .C(n_640), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_502), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx3_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
BUFx2_ASAP7_75t_L g566 ( .A(n_512), .Y(n_566) );
AND2x2_ASAP7_75t_L g580 ( .A(n_512), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g597 ( .A(n_512), .Y(n_597) );
OR2x2_ASAP7_75t_L g616 ( .A(n_512), .B(n_556), .Y(n_616) );
INVx3_ASAP7_75t_L g624 ( .A(n_512), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_512), .B(n_556), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_526), .B1(n_530), .B2(n_535), .C(n_547), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_523), .B(n_596), .Y(n_721) );
OR2x2_ASAP7_75t_L g724 ( .A(n_523), .B(n_555), .Y(n_724) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
OAI221xp5_ASAP7_75t_SL g547 ( .A1(n_524), .A2(n_548), .B1(n_555), .B2(n_557), .C(n_560), .Y(n_547) );
AND2x2_ASAP7_75t_L g564 ( .A(n_524), .B(n_556), .Y(n_564) );
AND2x2_ASAP7_75t_L g572 ( .A(n_524), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_524), .B(n_580), .Y(n_579) );
NAND2x1_ASAP7_75t_L g622 ( .A(n_524), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g674 ( .A(n_524), .B(n_616), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_526), .A2(n_634), .B1(n_663), .B2(n_665), .Y(n_662) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI322xp5_ASAP7_75t_L g571 ( .A1(n_527), .A2(n_536), .A3(n_572), .B1(n_575), .B2(n_578), .C1(n_582), .C2(n_585), .Y(n_571) );
OR2x2_ASAP7_75t_L g583 ( .A(n_527), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_528), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g562 ( .A(n_528), .B(n_537), .Y(n_562) );
INVx1_ASAP7_75t_L g577 ( .A(n_528), .Y(n_577) );
AND2x2_ASAP7_75t_L g643 ( .A(n_528), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g553 ( .A(n_529), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_529), .B(n_552), .Y(n_718) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_533), .B(n_667), .Y(n_666) );
INVx3_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g618 ( .A(n_534), .B(n_565), .Y(n_618) );
OR2x2_ASAP7_75t_L g715 ( .A(n_534), .B(n_566), .Y(n_715) );
INVx1_ASAP7_75t_L g696 ( .A(n_535), .Y(n_696) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_546), .Y(n_535) );
INVx4_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_536), .B(n_603), .Y(n_609) );
INVx2_ASAP7_75t_L g552 ( .A(n_537), .Y(n_552) );
INVx1_ASAP7_75t_L g634 ( .A(n_546), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_546), .B(n_606), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_548), .A2(n_622), .B(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g606 ( .A(n_552), .Y(n_606) );
INVx1_ASAP7_75t_L g633 ( .A(n_552), .Y(n_633) );
INVx1_ASAP7_75t_L g559 ( .A(n_553), .Y(n_559) );
AND2x2_ASAP7_75t_L g561 ( .A(n_553), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g657 ( .A(n_554), .B(n_643), .Y(n_657) );
AND2x2_ASAP7_75t_L g679 ( .A(n_554), .B(n_639), .Y(n_679) );
BUFx2_ASAP7_75t_L g631 ( .A(n_556), .Y(n_631) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AOI32xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .A3(n_564), .B1(n_565), .B2(n_567), .Y(n_560) );
INVx1_ASAP7_75t_L g641 ( .A(n_561), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_561), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_564), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_564), .B(n_623), .Y(n_664) );
AND2x2_ASAP7_75t_L g711 ( .A(n_564), .B(n_596), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_565), .B(n_612), .Y(n_659) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g712 ( .A(n_567), .Y(n_712) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_570), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g684 ( .A(n_570), .B(n_604), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_570), .B(n_599), .Y(n_691) );
INVx1_ASAP7_75t_SL g673 ( .A(n_572), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_573), .B(n_624), .Y(n_651) );
NOR4xp25_ASAP7_75t_L g697 ( .A(n_573), .B(n_596), .C(n_698), .D(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_574), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVxp67_ASAP7_75t_L g654 ( .A(n_577), .Y(n_654) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_580), .A2(n_671), .B(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g596 ( .A(n_581), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g645 ( .A(n_584), .Y(n_645) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND4xp25_ASAP7_75t_SL g587 ( .A(n_588), .B(n_613), .C(n_628), .D(n_648), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_594), .B(n_598), .C(n_600), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g680 ( .A(n_593), .B(n_623), .Y(n_680) );
AND2x2_ASAP7_75t_L g689 ( .A(n_593), .B(n_667), .Y(n_689) );
INVx3_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_596), .B(n_631), .Y(n_693) );
AND2x2_ASAP7_75t_L g605 ( .A(n_599), .B(n_606), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_607), .B1(n_609), .B2(n_610), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
AND2x2_ASAP7_75t_L g703 ( .A(n_603), .B(n_649), .Y(n_703) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_605), .B(n_654), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_606), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B(n_619), .C(n_621), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_614), .A2(n_649), .B1(n_650), .B2(n_652), .C(n_655), .Y(n_648) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_622), .A2(n_707), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_623), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_631), .B(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_636), .A2(n_656), .B1(n_658), .B2(n_659), .Y(n_655) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_645), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_656), .A2(n_682), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g701 ( .A(n_658), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_668), .C(n_688), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_681), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_675), .C(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g700 ( .A(n_678), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g722 ( .A1(n_679), .A2(n_705), .B(n_723), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_691), .A2(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .C(n_719), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_702), .C(n_704), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
CKINVDCx14_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g739 ( .A(n_725), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_729), .Y(n_740) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule