module fake_ibex_1619_n_1820 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1820);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1820;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_981;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_864;
wire n_608;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_1179;
wire n_907;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_1491;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_341),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_76),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_328),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_8),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_23),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_258),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_78),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_10),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_160),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_59),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_133),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_249),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_270),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_171),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_82),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_245),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_234),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_339),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_321),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_247),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_122),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_59),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_36),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_261),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_169),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_292),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_223),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_271),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_127),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_364),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_297),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_126),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_82),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_31),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_340),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_20),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_298),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_202),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_268),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_301),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_372),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_324),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_121),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_124),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_116),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_138),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_181),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_205),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_149),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_199),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_52),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_16),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_212),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_166),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_344),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_79),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_107),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_120),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_143),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_327),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_38),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_154),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_330),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_375),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_182),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_317),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_110),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_291),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_307),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_123),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_305),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_282),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_136),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_45),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_132),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_44),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_27),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_108),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_294),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_352),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_21),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_16),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_356),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_224),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_44),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_204),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_37),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_345),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_9),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_218),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_10),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_129),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_306),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_242),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_368),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_315),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_359),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_34),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_144),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_48),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_248),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_313),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_179),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_58),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_320),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_265),
.Y(n_488)
);

BUFx5_ASAP7_75t_L g489 ( 
.A(n_188),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_173),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_333),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_323),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_334),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_194),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_288),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_262),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_94),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_272),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_280),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_342),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_326),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_347),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_263),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_111),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_308),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_252),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_196),
.Y(n_507)
);

BUFx2_ASAP7_75t_SL g508 ( 
.A(n_183),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_158),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_164),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_31),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_43),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_81),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_348),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_134),
.Y(n_515)
);

BUFx8_ASAP7_75t_SL g516 ( 
.A(n_189),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_331),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_186),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_29),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_279),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_64),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_237),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_311),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_336),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_350),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_351),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_363),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_25),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_353),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_21),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_230),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_142),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_260),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_277),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_29),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_314),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_289),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_346),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_64),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_309),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_190),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_150),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_243),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_155),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_176),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_22),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_303),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_235),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_355),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_365),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_361),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_13),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_228),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_293),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_170),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_366),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_318),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_34),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_172),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_117),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_358),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_259),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_231),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_57),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_72),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_69),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_203),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_125),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_290),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_319),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_76),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_325),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_72),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_267),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_275),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_360),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_81),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_338),
.Y(n_578)
);

BUFx5_ASAP7_75t_L g579 ( 
.A(n_238),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_362),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_349),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_286),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_257),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_103),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_201),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_198),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_148),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_70),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_310),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_107),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_370),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_80),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_46),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_329),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_17),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_141),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_278),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_151),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_264),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_12),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_121),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_332),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_89),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_266),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_87),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_281),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_213),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_316),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_337),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_369),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_161),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_115),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_71),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_232),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_343),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_269),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_357),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_88),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_191),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_221),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_283),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_285),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_335),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_276),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_25),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_226),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_284),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_214),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_63),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_97),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_6),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_322),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_516),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_440),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_538),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_516),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_382),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_385),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_620),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_436),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_406),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_463),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_425),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_458),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_463),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_471),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_459),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_471),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_590),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_457),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_379),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_592),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_592),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_401),
.B(n_0),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_456),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_403),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_434),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_468),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_483),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_595),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_460),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_480),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_497),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_488),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_498),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_423),
.B(n_381),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_511),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_512),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_544),
.Y(n_673)
);

CKINVDCx16_ASAP7_75t_R g674 ( 
.A(n_520),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_535),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_564),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_534),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_585),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_565),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_573),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_577),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_534),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_591),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_612),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_613),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_630),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_393),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_393),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_466),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_466),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_388),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_392),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_551),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_395),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_551),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_397),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_383),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_489),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_415),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_419),
.B(n_421),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_387),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_402),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_426),
.B(n_0),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_389),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_430),
.Y(n_708)
);

INVxp33_ASAP7_75t_SL g709 ( 
.A(n_394),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_413),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_431),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_402),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_386),
.B(n_414),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_417),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_482),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_427),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_648),
.B(n_482),
.Y(n_717)
);

BUFx8_ASAP7_75t_L g718 ( 
.A(n_716),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_659),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_678),
.A2(n_438),
.B1(n_439),
.B2(n_433),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_701),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_701),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_660),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_699),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_699),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_645),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_643),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_646),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_694),
.B(n_462),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_647),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_656),
.B(n_443),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_667),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_649),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_712),
.B(n_508),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_713),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_635),
.B(n_519),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_675),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_638),
.B(n_519),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_676),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_690),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_677),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_680),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_681),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_657),
.A2(n_518),
.B(n_462),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_682),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_709),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_687),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_650),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_689),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_654),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_655),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_695),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_697),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_698),
.B(n_489),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_702),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_672),
.B(n_449),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_691),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_672),
.B(n_464),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_711),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_670),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_703),
.A2(n_531),
.B(n_518),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_706),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_700),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_664),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_641),
.B(n_467),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_692),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_685),
.B(n_531),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_686),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_693),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_639),
.A2(n_473),
.B1(n_504),
.B2(n_469),
.Y(n_776)
);

CKINVDCx6p67_ASAP7_75t_R g777 ( 
.A(n_674),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_640),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_707),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_696),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_710),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_714),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_633),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_715),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_715),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_636),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_705),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_705),
.B(n_532),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_637),
.B(n_513),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_642),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_644),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_652),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_661),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_662),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_668),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_669),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_673),
.Y(n_799)
);

OA21x2_ASAP7_75t_L g800 ( 
.A1(n_679),
.A2(n_550),
.B(n_532),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_634),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_678),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_683),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_684),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_684),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_688),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_653),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_688),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_663),
.Y(n_810)
);

NOR2x1_ASAP7_75t_L g811 ( 
.A(n_653),
.B(n_435),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_658),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_658),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_663),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_659),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_659),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_633),
.Y(n_817)
);

CKINVDCx8_ASAP7_75t_R g818 ( 
.A(n_641),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_701),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_635),
.B(n_519),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_659),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_699),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_699),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_701),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_701),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_716),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_659),
.Y(n_828)
);

OA21x2_ASAP7_75t_L g829 ( 
.A1(n_701),
.A2(n_594),
.B(n_550),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_635),
.B(n_519),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_699),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_694),
.B(n_594),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_659),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_638),
.B(n_404),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_635),
.B(n_397),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_699),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_659),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_701),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_699),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_701),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_699),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_701),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_699),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_699),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_701),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_648),
.B(n_521),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_659),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_599),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_659),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_648),
.B(n_528),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_701),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_701),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_659),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_701),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_699),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_699),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_698),
.B(n_489),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_701),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_659),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_648),
.B(n_530),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_701),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_738),
.A2(n_726),
.B1(n_774),
.B2(n_778),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_725),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_766),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_759),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_759),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_726),
.B(n_539),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_769),
.B(n_378),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_759),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_829),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_737),
.B(n_475),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_718),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_829),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_728),
.Y(n_879)
);

BUFx10_ASAP7_75t_L g880 ( 
.A(n_784),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_728),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_725),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_725),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_738),
.B(n_546),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_760),
.B(n_763),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_728),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_804),
.A2(n_424),
.B1(n_384),
.B2(n_441),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_725),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_739),
.Y(n_889)
);

AND3x4_ASAP7_75t_L g890 ( 
.A(n_814),
.B(n_576),
.C(n_541),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_739),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_820),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_728),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_765),
.A2(n_448),
.B1(n_452),
.B2(n_442),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_756),
.B(n_380),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_827),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_775),
.A2(n_566),
.B1(n_571),
.B2(n_552),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_749),
.A2(n_588),
.B1(n_593),
.B2(n_584),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_767),
.B(n_489),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_761),
.B(n_428),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_L g901 ( 
.A(n_767),
.B(n_489),
.Y(n_901)
);

BUFx4f_ASAP7_75t_L g902 ( 
.A(n_777),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_733),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_718),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_757),
.B(n_762),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_848),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_735),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_831),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_735),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_781),
.B(n_782),
.Y(n_910)
);

XNOR2xp5_ASAP7_75t_L g911 ( 
.A(n_720),
.B(n_600),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_749),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_779),
.B(n_541),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_761),
.B(n_390),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_820),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_768),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_773),
.A2(n_603),
.B1(n_605),
.B2(n_601),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_830),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_735),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_771),
.B(n_767),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_818),
.A2(n_625),
.B1(n_631),
.B2(n_618),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_800),
.A2(n_767),
.B1(n_719),
.B2(n_730),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_824),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_852),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_762),
.B(n_391),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_764),
.B(n_396),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_864),
.B(n_576),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_735),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_755),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_830),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_771),
.B(n_398),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_743),
.B(n_836),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_831),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_764),
.B(n_399),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_R g935 ( 
.A(n_817),
.B(n_799),
.Y(n_935)
);

NOR2x1p5_ASAP7_75t_L g936 ( 
.A(n_817),
.B(n_400),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_741),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_723),
.B(n_405),
.Y(n_938)
);

INVx6_ASAP7_75t_L g939 ( 
.A(n_784),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_755),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_755),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_407),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_734),
.B(n_408),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_736),
.B(n_409),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_740),
.B(n_410),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_845),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_737),
.B(n_580),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_755),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_742),
.B(n_411),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_790),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_824),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_744),
.B(n_412),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_732),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_814),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_808),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_745),
.B(n_416),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_845),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_858),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_743),
.B(n_418),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_722),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_732),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_721),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_721),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_741),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_836),
.B(n_422),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_859),
.B(n_746),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_754),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_791),
.Y(n_968)
);

BUFx10_ASAP7_75t_L g969 ( 
.A(n_784),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_808),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_791),
.B(n_429),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_780),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_858),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_727),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_751),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_859),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_748),
.B(n_437),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_750),
.B(n_446),
.Y(n_978)
);

AND2x6_ASAP7_75t_L g979 ( 
.A(n_784),
.B(n_580),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_SL g980 ( 
.A(n_789),
.B(n_451),
.C(n_450),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_717),
.B(n_432),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_770),
.B(n_444),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_860),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_752),
.B(n_454),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_753),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_860),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_722),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_772),
.B(n_776),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_724),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_855),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_815),
.B(n_465),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_835),
.B(n_445),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_822),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_800),
.A2(n_461),
.B1(n_476),
.B2(n_453),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_787),
.B(n_485),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_816),
.B(n_470),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_855),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_798),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_772),
.B(n_447),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_837),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_841),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_780),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_786),
.B(n_1),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_474),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_823),
.B(n_472),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_843),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_SL g1007 ( 
.A1(n_729),
.A2(n_509),
.B(n_496),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_846),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_828),
.B(n_477),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_722),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_788),
.B(n_1),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_833),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_834),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_787),
.B(n_515),
.Y(n_1014)
);

BUFx8_ASAP7_75t_SL g1015 ( 
.A(n_812),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_787),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_737),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_722),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_819),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_838),
.B(n_478),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_839),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_849),
.A2(n_522),
.B1(n_524),
.B2(n_517),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_851),
.B(n_479),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_797),
.B(n_2),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_856),
.B(n_863),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_835),
.B(n_481),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_747),
.A2(n_529),
.B1(n_543),
.B2(n_527),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_729),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_832),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_787),
.B(n_484),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_819),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_832),
.B(n_850),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_850),
.B(n_847),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_847),
.B(n_487),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_819),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_819),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_792),
.B(n_501),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_825),
.Y(n_1039)
);

AO21x2_ASAP7_75t_L g1040 ( 
.A1(n_857),
.A2(n_553),
.B(n_549),
.Y(n_1040)
);

NOR2x1p5_ASAP7_75t_L g1041 ( 
.A(n_799),
.B(n_490),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_747),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_825),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_825),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_825),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_826),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_789),
.A2(n_570),
.B1(n_572),
.B2(n_555),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_857),
.B(n_492),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_793),
.B(n_578),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_847),
.B(n_493),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_826),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_865),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_826),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_826),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_840),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_840),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_840),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_794),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_840),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_798),
.B(n_582),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_842),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_842),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_847),
.B(n_795),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_796),
.B(n_583),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_794),
.B(n_587),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_758),
.B(n_494),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_842),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_842),
.B(n_495),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_844),
.Y(n_1070)
);

NOR2x1p5_ASAP7_75t_L g1071 ( 
.A(n_812),
.B(n_785),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_783),
.B(n_628),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_844),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_844),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_797),
.B(n_2),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_758),
.A2(n_604),
.B1(n_606),
.B2(n_598),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_844),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_794),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_794),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_811),
.B(n_499),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_853),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_810),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_801),
.B(n_632),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_861),
.B(n_500),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_861),
.B(n_502),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_853),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_853),
.B(n_503),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_853),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_862),
.Y(n_1089)
);

INVx11_ASAP7_75t_L g1090 ( 
.A(n_810),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_862),
.A2(n_608),
.B1(n_609),
.B2(n_607),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_862),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_802),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_962),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_1017),
.B(n_505),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_912),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_962),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_988),
.A2(n_885),
.B1(n_1030),
.B2(n_1029),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_871),
.B(n_802),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_866),
.B(n_805),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1033),
.B(n_862),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_905),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1012),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_903),
.B(n_807),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_896),
.A2(n_803),
.B1(n_802),
.B2(n_806),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1013),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_968),
.B(n_802),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_906),
.B(n_809),
.Y(n_1108)
);

OAI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_924),
.A2(n_813),
.B1(n_803),
.B2(n_806),
.C(n_610),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_999),
.B(n_506),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1082),
.A2(n_803),
.B1(n_806),
.B2(n_615),
.C(n_507),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_890),
.A2(n_803),
.B1(n_806),
.B2(n_602),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1017),
.B(n_510),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1021),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_916),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_L g1116 ( 
.A(n_910),
.B(n_489),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1024),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_971),
.B(n_627),
.Y(n_1118)
);

OAI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_972),
.A2(n_525),
.B1(n_526),
.B2(n_514),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1026),
.A2(n_602),
.B1(n_599),
.B2(n_455),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_889),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_891),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_892),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_SL g1124 ( 
.A(n_998),
.B(n_533),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_915),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_918),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_SL g1127 ( 
.A(n_980),
.B(n_536),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_930),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_884),
.B(n_537),
.Y(n_1129)
);

INVx8_ASAP7_75t_L g1130 ( 
.A(n_1078),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1005),
.B(n_540),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_950),
.B(n_542),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_963),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_963),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_982),
.A2(n_548),
.B1(n_554),
.B2(n_545),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_932),
.B(n_556),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_917),
.B(n_557),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1078),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1002),
.B(n_3),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_L g1140 ( 
.A(n_921),
.B(n_561),
.C(n_559),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_937),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_898),
.B(n_624),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_562),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_927),
.B(n_563),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_876),
.B(n_567),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1047),
.B(n_569),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_947),
.B(n_900),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_876),
.B(n_574),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_923),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_990),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_981),
.A2(n_581),
.B1(n_586),
.B2(n_575),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1090),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1061),
.B(n_3),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1049),
.B(n_589),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_947),
.B(n_596),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1049),
.B(n_597),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_L g1157 ( 
.A(n_970),
.B(n_616),
.C(n_611),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_990),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_877),
.B(n_4),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1071),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1061),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_994),
.B(n_617),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1041),
.B(n_4),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_922),
.A2(n_455),
.B1(n_523),
.B2(n_420),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1007),
.B(n_619),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_904),
.B(n_5),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1049),
.B(n_621),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1049),
.B(n_622),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_895),
.B(n_623),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1065),
.B(n_579),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_938),
.B(n_579),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1065),
.B(n_579),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_964),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1065),
.B(n_579),
.Y(n_1174)
);

OAI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_894),
.A2(n_523),
.B1(n_547),
.B2(n_455),
.C(n_420),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_965),
.B(n_1083),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1065),
.A2(n_579),
.B1(n_455),
.B2(n_523),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1080),
.B(n_5),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_942),
.B(n_579),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1072),
.B(n_6),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_953),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_997),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_974),
.B(n_7),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_880),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_997),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_875),
.B(n_420),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_975),
.B(n_7),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_887),
.A2(n_547),
.B1(n_568),
.B2(n_523),
.C(n_420),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_992),
.A2(n_568),
.B1(n_547),
.B2(n_614),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_887),
.B(n_8),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_985),
.B(n_897),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_953),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_902),
.A2(n_568),
.B1(n_614),
.B2(n_547),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_911),
.B(n_9),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_943),
.B(n_11),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_944),
.B(n_11),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_945),
.B(n_949),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_SL g1198 ( 
.A(n_935),
.B(n_614),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1027),
.B(n_12),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_961),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_952),
.B(n_13),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_961),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_902),
.B(n_14),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_956),
.B(n_568),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_977),
.B(n_614),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_978),
.B(n_14),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_SL g1207 ( 
.A(n_1015),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1025),
.A2(n_18),
.B(n_15),
.C(n_17),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1038),
.B(n_15),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_984),
.B(n_18),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1075),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_868),
.A2(n_130),
.B(n_128),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_989),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_996),
.B(n_1004),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1003),
.B(n_19),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_993),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1009),
.B(n_19),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_880),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1023),
.B(n_20),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_873),
.B(n_22),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1000),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1011),
.A2(n_26),
.B(n_23),
.C(n_24),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_936),
.B(n_24),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1053),
.B(n_26),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1022),
.B(n_27),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1028),
.B(n_28),
.C(n_30),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1076),
.B(n_28),
.Y(n_1227)
);

NOR3xp33_ASAP7_75t_L g1228 ( 
.A(n_914),
.B(n_30),
.C(n_32),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_920),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_910),
.B(n_32),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_908),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_910),
.B(n_33),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_910),
.B(n_131),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1052),
.B(n_925),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_991),
.B(n_33),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_926),
.B(n_35),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_955),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_934),
.B(n_35),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_868),
.A2(n_137),
.B(n_135),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_954),
.B(n_36),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_983),
.B(n_37),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1020),
.B(n_38),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_951),
.B(n_39),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1093),
.B(n_39),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_888),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_976),
.B(n_40),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_933),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_983),
.B(n_40),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1042),
.B(n_41),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_875),
.B(n_41),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_946),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_957),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_931),
.B(n_42),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_969),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_878),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_L g1256 ( 
.A(n_878),
.B(n_139),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1064),
.B(n_959),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1040),
.B(n_46),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_986),
.B(n_47),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1001),
.Y(n_1260)
);

INVx8_ASAP7_75t_L g1261 ( 
.A(n_1066),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1006),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_958),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1059),
.B(n_47),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_L g1265 ( 
.A(n_979),
.B(n_140),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1079),
.B(n_48),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1008),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1066),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1067),
.B(n_49),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_969),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_986),
.B(n_49),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1016),
.B(n_50),
.Y(n_1272)
);

BUFx5_ASAP7_75t_L g1273 ( 
.A(n_1054),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1040),
.B(n_50),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_L g1275 ( 
.A(n_979),
.B(n_145),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_973),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_879),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1085),
.B(n_51),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1084),
.B(n_51),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_913),
.B(n_52),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_939),
.B(n_53),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1034),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1098),
.B(n_1102),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1096),
.B(n_1153),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1161),
.B(n_939),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1103),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1239),
.A2(n_901),
.B(n_899),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1130),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1106),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1186),
.A2(n_1048),
.B(n_966),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1114),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1211),
.B(n_913),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1117),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1095),
.B(n_919),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1208),
.A2(n_1069),
.B(n_1050),
.C(n_1035),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1115),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1095),
.B(n_919),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1186),
.A2(n_1063),
.B(n_1054),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1207),
.B(n_979),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1222),
.A2(n_1091),
.B(n_1087),
.C(n_886),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1130),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1100),
.B(n_1191),
.Y(n_1302)
);

INVxp67_ASAP7_75t_SL g1303 ( 
.A(n_1101),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1197),
.A2(n_1073),
.B(n_1063),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1094),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1214),
.A2(n_1088),
.B(n_1073),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1101),
.A2(n_1092),
.B(n_1088),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1234),
.A2(n_1092),
.B(n_870),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1097),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1209),
.A2(n_886),
.B(n_928),
.C(n_879),
.Y(n_1310)
);

AOI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1132),
.A2(n_929),
.B(n_928),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1099),
.B(n_913),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1178),
.B(n_913),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1133),
.A2(n_919),
.B1(n_987),
.B2(n_960),
.Y(n_1314)
);

AO21x1_ASAP7_75t_L g1315 ( 
.A1(n_1239),
.A2(n_870),
.B(n_869),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1256),
.A2(n_872),
.B(n_869),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1171),
.A2(n_874),
.B(n_872),
.Y(n_1317)
);

CKINVDCx10_ASAP7_75t_R g1318 ( 
.A(n_1237),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1147),
.B(n_1031),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1104),
.A2(n_1066),
.B1(n_995),
.B2(n_1014),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1179),
.A2(n_874),
.B(n_1055),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1181),
.A2(n_1057),
.B(n_1018),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1109),
.A2(n_1279),
.B(n_1225),
.C(n_1105),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1192),
.A2(n_1202),
.B(n_1200),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1162),
.A2(n_1019),
.B(n_1010),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1124),
.B(n_960),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1164),
.A2(n_882),
.B(n_867),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1119),
.B(n_960),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_1258),
.B(n_1274),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1270),
.B(n_987),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_L g1331 ( 
.A(n_1270),
.B(n_987),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1143),
.A2(n_1036),
.B(n_1032),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1134),
.A2(n_1158),
.B(n_1150),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1182),
.A2(n_1044),
.B(n_1037),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1176),
.B(n_1066),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1217),
.A2(n_1269),
.B(n_1278),
.C(n_1227),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1185),
.A2(n_1074),
.B1(n_1046),
.B2(n_893),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1121),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1180),
.A2(n_948),
.B(n_929),
.C(n_893),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1107),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1152),
.B(n_881),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1130),
.B(n_1138),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1138),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1160),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1122),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1184),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1245),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1277),
.A2(n_1051),
.B(n_1045),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1108),
.A2(n_1014),
.B1(n_995),
.B2(n_979),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1218),
.B(n_1046),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1116),
.A2(n_1110),
.B(n_1224),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1129),
.B(n_881),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1195),
.A2(n_1060),
.B(n_1056),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1250),
.A2(n_948),
.B(n_1062),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1250),
.A2(n_1081),
.B(n_1068),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1240),
.B(n_1190),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1236),
.A2(n_1089),
.B(n_1086),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1238),
.A2(n_1201),
.B(n_1196),
.Y(n_1358)
);

OAI21xp33_ASAP7_75t_L g1359 ( 
.A1(n_1131),
.A2(n_1144),
.B(n_1112),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1254),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1123),
.B(n_995),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1149),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1206),
.A2(n_883),
.B(n_1043),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1149),
.B(n_1268),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1163),
.B(n_1046),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1125),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1245),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1163),
.B(n_888),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1210),
.A2(n_1070),
.B(n_1043),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1261),
.B(n_888),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1219),
.A2(n_1077),
.B(n_1070),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1155),
.B(n_907),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1126),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1165),
.A2(n_1120),
.B(n_1246),
.C(n_1243),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1128),
.B(n_1074),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1169),
.A2(n_1077),
.B(n_909),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1220),
.A2(n_909),
.B(n_940),
.C(n_907),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1136),
.A2(n_941),
.B(n_940),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1141),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1173),
.B(n_995),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_941),
.B(n_1074),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_L g1383 ( 
.A1(n_1198),
.A2(n_1014),
.B(n_1058),
.C(n_1039),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1229),
.A2(n_1039),
.B(n_1058),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1120),
.A2(n_1014),
.B(n_56),
.C(n_54),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1213),
.A2(n_1039),
.B(n_1058),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1215),
.B(n_55),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1261),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1216),
.A2(n_147),
.B(n_146),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1221),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1203),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1245),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1151),
.B(n_56),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1199),
.B(n_57),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1260),
.A2(n_153),
.B(n_152),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1183),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1187),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1111),
.A2(n_61),
.B1(n_58),
.B2(n_60),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1249),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1135),
.B(n_62),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1262),
.A2(n_157),
.B(n_156),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1157),
.B(n_63),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1267),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1166),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1223),
.B(n_65),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1233),
.A2(n_162),
.B(n_159),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1231),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1139),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1247),
.A2(n_165),
.B(n_163),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1235),
.B(n_65),
.Y(n_1410)
);

NOR3xp33_ASAP7_75t_L g1411 ( 
.A(n_1194),
.B(n_66),
.C(n_67),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1204),
.A2(n_168),
.B(n_167),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1251),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1255),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1252),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1255),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1263),
.A2(n_175),
.B(n_174),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1242),
.B(n_66),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1205),
.A2(n_178),
.B(n_177),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1188),
.A2(n_1228),
.B1(n_1226),
.B2(n_1253),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1140),
.B(n_67),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1282),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1276),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1154),
.B(n_68),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1145),
.B(n_71),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1258),
.A2(n_73),
.B(n_74),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1148),
.B(n_73),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1404),
.B(n_1137),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1301),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1414),
.A2(n_1127),
.B1(n_1142),
.B2(n_1226),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1286),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1316),
.A2(n_1212),
.B(n_1172),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1301),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1288),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1289),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1351),
.A2(n_1174),
.B(n_1170),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1344),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1298),
.A2(n_1248),
.B(n_1241),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1358),
.A2(n_1271),
.B(n_1259),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_SL g1440 ( 
.A(n_1411),
.B(n_1113),
.C(n_1189),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1318),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1290),
.A2(n_1275),
.B(n_1265),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1336),
.A2(n_1264),
.B(n_1257),
.C(n_1230),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1305),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1315),
.A2(n_1384),
.B(n_1386),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1343),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1302),
.B(n_1146),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1353),
.A2(n_1266),
.B(n_1232),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1332),
.A2(n_1175),
.B(n_1167),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1347),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1355),
.A2(n_1168),
.B(n_1156),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1420),
.A2(n_1323),
.B(n_1300),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1375),
.A2(n_1159),
.B(n_1280),
.C(n_1177),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1365),
.B(n_1272),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1391),
.B(n_1281),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1347),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1283),
.B(n_1244),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1318),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1294),
.A2(n_1118),
.B(n_1193),
.C(n_1273),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1347),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1296),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1329),
.A2(n_1273),
.B(n_273),
.C(n_274),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1291),
.B(n_1273),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1343),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1293),
.B(n_1273),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1340),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1342),
.B(n_74),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1356),
.B(n_1273),
.Y(n_1469)
);

AND2x6_ASAP7_75t_L g1470 ( 
.A(n_1416),
.B(n_75),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1284),
.B(n_75),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1304),
.A2(n_184),
.B(n_180),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1306),
.A2(n_187),
.B(n_185),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1393),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1359),
.A2(n_1422),
.B(n_1420),
.C(n_1397),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1346),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1338),
.B(n_1374),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1408),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1345),
.B(n_77),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1360),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1402),
.A2(n_80),
.B(n_83),
.C(n_84),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1363),
.A2(n_193),
.B(n_192),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1376),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1376),
.B(n_83),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1396),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_1485)
);

OAI21xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1303),
.A2(n_1417),
.B(n_1409),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1366),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1310),
.A2(n_197),
.B(n_195),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1385),
.A2(n_85),
.B(n_86),
.C(n_87),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1320),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1297),
.A2(n_287),
.B(n_377),
.C(n_376),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1380),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1308),
.A2(n_206),
.B(n_200),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1339),
.A2(n_208),
.B(n_207),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1423),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1369),
.A2(n_210),
.B(n_209),
.Y(n_1496)
);

AOI22x1_ASAP7_75t_L g1497 ( 
.A1(n_1406),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1371),
.A2(n_215),
.B(n_211),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1373),
.B(n_91),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1367),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1287),
.A2(n_217),
.B(n_216),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1421),
.A2(n_92),
.B(n_93),
.C(n_94),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1407),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1307),
.A2(n_222),
.B(n_219),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1354),
.A2(n_1357),
.B(n_1334),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_SL g1506 ( 
.A1(n_1378),
.A2(n_296),
.B(n_374),
.C(n_373),
.Y(n_1506)
);

BUFx5_ASAP7_75t_L g1507 ( 
.A(n_1362),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1295),
.A2(n_93),
.B(n_95),
.C(n_96),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1367),
.Y(n_1509)
);

OAI321xp33_ASAP7_75t_L g1510 ( 
.A1(n_1426),
.A2(n_95),
.A3(n_96),
.B1(n_97),
.B2(n_98),
.C(n_99),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1427),
.B(n_98),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1352),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1349),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1373),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1299),
.B(n_102),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1348),
.A2(n_302),
.B(n_371),
.Y(n_1516)
);

AO31x2_ASAP7_75t_L g1517 ( 
.A1(n_1445),
.A2(n_1387),
.A3(n_1399),
.B(n_1389),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1453),
.A2(n_1327),
.B(n_1382),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1505),
.A2(n_1401),
.A3(n_1395),
.B(n_1324),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1486),
.A2(n_1333),
.B(n_1367),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1442),
.A2(n_1313),
.B(n_1383),
.Y(n_1521)
);

INVx4_ASAP7_75t_SL g1522 ( 
.A(n_1429),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1456),
.B(n_1425),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1511),
.A2(n_1455),
.B1(n_1474),
.B2(n_1458),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1468),
.B(n_1368),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_1467),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1481),
.A2(n_1398),
.B(n_1319),
.C(n_1394),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1462),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1413),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1475),
.A2(n_1418),
.B(n_1410),
.C(n_1405),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1439),
.A2(n_1325),
.B(n_1322),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1431),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1447),
.B(n_1400),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1438),
.A2(n_1292),
.B(n_1392),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1435),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1455),
.A2(n_1335),
.B1(n_1415),
.B2(n_1312),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1433),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1463),
.A2(n_1392),
.B(n_1321),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1432),
.A2(n_1317),
.B(n_1379),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1436),
.A2(n_1419),
.B(n_1412),
.Y(n_1541)
);

AO32x2_ASAP7_75t_L g1542 ( 
.A1(n_1490),
.A2(n_1314),
.A3(n_1337),
.B1(n_1424),
.B2(n_1311),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1441),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_SL g1544 ( 
.A(n_1437),
.B(n_1388),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1448),
.A2(n_1377),
.B(n_1415),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1471),
.A2(n_1285),
.B1(n_1372),
.B2(n_1361),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_L g1547 ( 
.A(n_1429),
.B(n_1507),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1477),
.Y(n_1548)
);

AO22x2_ASAP7_75t_L g1549 ( 
.A1(n_1484),
.A2(n_1326),
.B1(n_1350),
.B2(n_1328),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1449),
.A2(n_1381),
.B(n_1370),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1454),
.A2(n_1370),
.B(n_1390),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1487),
.Y(n_1552)
);

AOI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1430),
.A2(n_1370),
.B(n_1341),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1428),
.A2(n_1331),
.B1(n_1330),
.B2(n_1388),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1489),
.A2(n_1403),
.B(n_1364),
.C(n_1331),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1503),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1480),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1451),
.A2(n_1330),
.B(n_304),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1499),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1478),
.B(n_103),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1444),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1443),
.A2(n_300),
.B(n_367),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1524),
.A2(n_1512),
.B1(n_1469),
.B2(n_1485),
.Y(n_1563)
);

INVx6_ASAP7_75t_L g1564 ( 
.A(n_1522),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1523),
.A2(n_1470),
.B1(n_1440),
.B2(n_1513),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1537),
.A2(n_1508),
.B1(n_1483),
.B2(n_1497),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1532),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1535),
.B(n_1452),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1518),
.Y(n_1569)
);

INVx6_ASAP7_75t_L g1570 ( 
.A(n_1522),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1518),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1561),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1556),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1533),
.A2(n_1470),
.B1(n_1525),
.B2(n_1553),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1543),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

BUFx12f_ASAP7_75t_L g1577 ( 
.A(n_1529),
.Y(n_1577)
);

BUFx2_ASAP7_75t_SL g1578 ( 
.A(n_1554),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1559),
.A2(n_1464),
.B1(n_1466),
.B2(n_1479),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1528),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1546),
.A2(n_1515),
.B1(n_1465),
.B2(n_1502),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1549),
.A2(n_1470),
.B1(n_1459),
.B2(n_1437),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.Y(n_1583)
);

INVx6_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1548),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1545),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1536),
.A2(n_1507),
.B1(n_1446),
.B2(n_1514),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1526),
.Y(n_1589)
);

CKINVDCx11_ASAP7_75t_R g1590 ( 
.A(n_1547),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1540),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1560),
.A2(n_1510),
.B1(n_1476),
.B2(n_1434),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1567),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1583),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1588),
.Y(n_1597)
);

INVx4_ASAP7_75t_L g1598 ( 
.A(n_1590),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1585),
.B(n_1530),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1567),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1583),
.B(n_1517),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1517),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1577),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1589),
.B(n_1551),
.Y(n_1605)
);

AO21x2_ASAP7_75t_L g1606 ( 
.A1(n_1591),
.A2(n_1520),
.B(n_1521),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

AO21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1587),
.A2(n_1542),
.B(n_1507),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1584),
.A2(n_1562),
.B1(n_1558),
.B2(n_1501),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1576),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1588),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1594),
.B(n_1542),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1569),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1571),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.Y(n_1619)
);

BUFx5_ASAP7_75t_L g1620 ( 
.A(n_1592),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1568),
.B(n_1542),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1621),
.B(n_1571),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1604),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1604),
.B(n_1575),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1601),
.B(n_1603),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1621),
.B(n_1591),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1578),
.Y(n_1629)
);

CKINVDCx16_ASAP7_75t_R g1630 ( 
.A(n_1598),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1613),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1618),
.A2(n_1531),
.B(n_1534),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_SL g1633 ( 
.A1(n_1597),
.A2(n_1565),
.B(n_1574),
.C(n_1581),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1601),
.Y(n_1634)
);

AND2x4_ASAP7_75t_SL g1635 ( 
.A(n_1598),
.B(n_1592),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1618),
.A2(n_1550),
.B(n_1538),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1595),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1598),
.A2(n_1582),
.B1(n_1584),
.B2(n_1579),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1578),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1619),
.B(n_1586),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1615),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1634),
.B(n_1605),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1623),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1630),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1637),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1631),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1640),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1627),
.B(n_1616),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1635),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1634),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1629),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1615),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1627),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1640),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1644),
.B(n_1622),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1646),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1650),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1658),
.B(n_1622),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1646),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1647),
.A2(n_1638),
.B(n_1625),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1647),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1648),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1658),
.B(n_1639),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1652),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1649),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1655),
.B(n_1639),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1644),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1628),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1652),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

AOI33xp33_ASAP7_75t_L g1675 ( 
.A1(n_1645),
.A2(n_1635),
.A3(n_1631),
.B1(n_1612),
.B2(n_1593),
.B3(n_1628),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1651),
.B(n_1635),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1650),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1671),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1673),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1675),
.B(n_1654),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1666),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1665),
.B(n_1656),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1666),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1679),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1679),
.A2(n_1664),
.B(n_1638),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1678),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1681),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1683),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1684),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1685),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1685),
.B(n_1680),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1689),
.Y(n_1692)
);

AOI222xp33_ASAP7_75t_L g1693 ( 
.A1(n_1690),
.A2(n_1686),
.B1(n_1669),
.B2(n_1687),
.C1(n_1688),
.C2(n_1674),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1691),
.B(n_1673),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1690),
.A2(n_1630),
.B1(n_1674),
.B2(n_1668),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1689),
.B(n_1659),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_SL g1697 ( 
.A(n_1692),
.B(n_1564),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1696),
.B(n_1659),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1694),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1695),
.A2(n_1626),
.B1(n_1633),
.B2(n_1668),
.C(n_1607),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1693),
.Y(n_1701)
);

AOI222xp33_ASAP7_75t_L g1702 ( 
.A1(n_1692),
.A2(n_1682),
.B1(n_1668),
.B2(n_1676),
.C1(n_1663),
.C2(n_1660),
.Y(n_1702)
);

NAND4xp25_ASAP7_75t_L g1703 ( 
.A(n_1692),
.B(n_1676),
.C(n_1563),
.D(n_1599),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1698),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1701),
.A2(n_1575),
.B(n_1676),
.C(n_1682),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1699),
.A2(n_1670),
.B1(n_1651),
.B2(n_1620),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1703),
.Y(n_1707)
);

OAI22x1_ASAP7_75t_L g1708 ( 
.A1(n_1700),
.A2(n_1616),
.B1(n_1670),
.B2(n_1651),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1702),
.B(n_1660),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1697),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1701),
.B(n_1663),
.Y(n_1711)
);

OAI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1701),
.A2(n_1584),
.B1(n_1570),
.B2(n_1564),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1701),
.B(n_1661),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1701),
.B(n_1620),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1699),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1704),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1707),
.B(n_1564),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1710),
.B(n_1677),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1713),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1715),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1705),
.A2(n_1570),
.B1(n_1564),
.B2(n_1620),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1711),
.A2(n_1570),
.B1(n_1677),
.B2(n_1661),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1712),
.B(n_1620),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_SL g1724 ( 
.A(n_1709),
.B(n_1706),
.C(n_1708),
.D(n_1714),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_L g1725 ( 
.A(n_1707),
.B(n_1491),
.C(n_1527),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1704),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1704),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1704),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1704),
.B(n_1667),
.Y(n_1729)
);

NAND4xp25_ASAP7_75t_L g1730 ( 
.A(n_1705),
.B(n_1566),
.C(n_1667),
.D(n_1570),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1712),
.A2(n_1611),
.B(n_1655),
.C(n_1460),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1704),
.B(n_1662),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1726),
.B(n_1662),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1716),
.A2(n_1620),
.B1(n_1657),
.B2(n_1609),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1727),
.B(n_1620),
.Y(n_1735)
);

AOI211x1_ASAP7_75t_L g1736 ( 
.A1(n_1728),
.A2(n_1719),
.B(n_1724),
.C(n_1720),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1717),
.A2(n_1672),
.B1(n_1662),
.B2(n_1605),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1662),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1729),
.A2(n_1506),
.B(n_1488),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1723),
.A2(n_1725),
.B(n_1721),
.C(n_1722),
.Y(n_1740)
);

O2A1O1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1730),
.A2(n_1718),
.B(n_1722),
.C(n_1731),
.Y(n_1741)
);

OAI21xp33_ASAP7_75t_L g1742 ( 
.A1(n_1717),
.A2(n_1657),
.B(n_1600),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1717),
.A2(n_1595),
.B(n_1600),
.C(n_1494),
.Y(n_1743)
);

NOR4xp25_ASAP7_75t_L g1744 ( 
.A(n_1716),
.B(n_104),
.C(n_105),
.D(n_106),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1716),
.A2(n_1642),
.B1(n_1504),
.B2(n_1496),
.C(n_1498),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1726),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1716),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1716),
.A2(n_108),
.B(n_109),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1716),
.A2(n_1642),
.B1(n_1493),
.B2(n_1472),
.C(n_1473),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1746),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1736),
.A2(n_1516),
.B1(n_1482),
.B2(n_1642),
.C(n_1619),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1733),
.B(n_109),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1744),
.A2(n_1741),
.B1(n_1748),
.B2(n_1740),
.C(n_1747),
.Y(n_1753)
);

OAI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1735),
.A2(n_1642),
.B(n_1641),
.Y(n_1754)
);

OAI31xp33_ASAP7_75t_L g1755 ( 
.A1(n_1743),
.A2(n_1590),
.A3(n_111),
.B(n_112),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1738),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1742),
.A2(n_1608),
.B1(n_1610),
.B2(n_1617),
.Y(n_1757)
);

AOI211xp5_ASAP7_75t_L g1758 ( 
.A1(n_1737),
.A2(n_110),
.B(n_112),
.C(n_113),
.Y(n_1758)
);

OAI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1734),
.A2(n_1749),
.B(n_1739),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1745),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1746),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1746),
.A2(n_1620),
.B1(n_1507),
.B2(n_1592),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1746),
.A2(n_1620),
.B1(n_1641),
.B2(n_1632),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1746),
.A2(n_1632),
.B1(n_1606),
.B2(n_1608),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1746),
.A2(n_113),
.B(n_114),
.C(n_115),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1746),
.B(n_114),
.Y(n_1766)
);

NAND2xp33_ASAP7_75t_R g1767 ( 
.A(n_1746),
.B(n_116),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1746),
.A2(n_1632),
.B1(n_1606),
.B2(n_1586),
.Y(n_1768)
);

NAND4xp75_ASAP7_75t_L g1769 ( 
.A(n_1753),
.B(n_117),
.C(n_118),
.D(n_119),
.Y(n_1769)
);

BUFx12f_ASAP7_75t_L g1770 ( 
.A(n_1761),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1750),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1752),
.Y(n_1772)
);

NAND2x1p5_ASAP7_75t_L g1773 ( 
.A(n_1766),
.B(n_1450),
.Y(n_1773)
);

XOR2x2_ASAP7_75t_L g1774 ( 
.A(n_1758),
.B(n_118),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1762),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1760),
.B(n_1609),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1768),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1765),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1763),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_L g1780 ( 
.A(n_1759),
.B(n_119),
.Y(n_1780)
);

AOI22x1_ASAP7_75t_L g1781 ( 
.A1(n_1770),
.A2(n_1778),
.B1(n_1771),
.B2(n_1772),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1769),
.Y(n_1782)
);

NAND4xp75_ASAP7_75t_L g1783 ( 
.A(n_1780),
.B(n_1755),
.C(n_1751),
.D(n_1767),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1774),
.Y(n_1784)
);

AND3x4_ASAP7_75t_L g1785 ( 
.A(n_1779),
.B(n_1754),
.C(n_1764),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1778),
.B(n_1757),
.C(n_120),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1769),
.B(n_1775),
.C(n_1777),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1776),
.A2(n_1450),
.B1(n_1500),
.B2(n_1457),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1773),
.B(n_1457),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1770),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1771),
.B(n_1610),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1771),
.B(n_1632),
.Y(n_1792)
);

INVxp33_ASAP7_75t_SL g1793 ( 
.A(n_1790),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1781),
.A2(n_1787),
.B(n_1782),
.C(n_1786),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1791),
.B(n_225),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1792),
.B(n_1606),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1785),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1784),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1789),
.A2(n_1509),
.B(n_1500),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1783),
.B(n_227),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1788),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1798),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1797),
.B(n_1636),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1793),
.A2(n_1509),
.B1(n_1461),
.B2(n_1586),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1794),
.A2(n_1461),
.B1(n_1636),
.B2(n_1541),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1802),
.B(n_1800),
.Y(n_1806)
);

AOI22x1_ASAP7_75t_L g1807 ( 
.A1(n_1803),
.A2(n_1801),
.B1(n_1796),
.B2(n_1795),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1805),
.Y(n_1808)
);

AOI22x1_ASAP7_75t_SL g1809 ( 
.A1(n_1808),
.A2(n_1804),
.B1(n_1799),
.B2(n_236),
.Y(n_1809)
);

XNOR2xp5_ASAP7_75t_L g1810 ( 
.A(n_1806),
.B(n_229),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1807),
.B(n_1617),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1809),
.A2(n_1636),
.B1(n_239),
.B2(n_240),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1810),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1811),
.B(n_233),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1812),
.A2(n_1636),
.B1(n_1519),
.B2(n_246),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1813),
.B(n_241),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1814),
.A2(n_244),
.B(n_250),
.Y(n_1817)
);

BUFx4_ASAP7_75t_R g1818 ( 
.A(n_1817),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_R g1819 ( 
.A1(n_1818),
.A2(n_1815),
.B1(n_1816),
.B2(n_254),
.C(n_255),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_251),
.B(n_253),
.C(n_256),
.Y(n_1820)
);


endmodule