module fake_jpeg_1884_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_27),
.Y(n_28)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_26),
.B1(n_13),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_16),
.B1(n_13),
.B2(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_21),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_45),
.B1(n_31),
.B2(n_35),
.Y(n_50)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_35),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_42),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_38),
.B1(n_41),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_46),
.B1(n_45),
.B2(n_14),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_46),
.B1(n_15),
.B2(n_11),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_30),
.B(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.C(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_15),
.C(n_18),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_18),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_55),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_59),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_7),
.Y(n_64)
);


endmodule