module real_aes_16640_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_869;
wire n_613;
wire n_642;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g523 ( .A(n_0), .B(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_1), .A2(n_34), .B1(n_130), .B2(n_142), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_2), .A2(n_10), .B1(n_549), .B2(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g524 ( .A(n_3), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_4), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_11), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_6), .A2(n_859), .B1(n_865), .B2(n_866), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_6), .Y(n_865) );
OR2x2_ASAP7_75t_L g508 ( .A(n_7), .B(n_30), .Y(n_508) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_8), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_9), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_12), .B(n_181), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_13), .A2(n_100), .B1(n_178), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_14), .A2(n_31), .B1(n_572), .B2(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_15), .B(n_181), .Y(n_613) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_16), .A2(n_45), .B(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_17), .B(n_270), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_18), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_19), .A2(n_93), .B1(n_863), .B2(n_864), .Y(n_862) );
INVx1_ASAP7_75t_L g864 ( .A(n_19), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_20), .A2(n_38), .B1(n_168), .B2(n_186), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_21), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_22), .A2(n_43), .B1(n_168), .B2(n_549), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_23), .A2(n_81), .B1(n_497), .B2(n_498), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_23), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_24), .B(n_572), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_25), .B(n_133), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_26), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_27), .B(n_191), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_28), .Y(n_177) );
AOI22x1_ASAP7_75t_L g494 ( .A1(n_29), .A2(n_495), .B1(n_496), .B2(n_499), .Y(n_494) );
INVx1_ASAP7_75t_L g499 ( .A(n_29), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_32), .A2(n_84), .B1(n_130), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_33), .A2(n_37), .B1(n_130), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_35), .A2(n_48), .B1(n_549), .B2(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_36), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_39), .B(n_181), .Y(n_231) );
INVx2_ASAP7_75t_L g520 ( .A(n_40), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_41), .B(n_182), .Y(n_265) );
INVx1_ASAP7_75t_L g506 ( .A(n_42), .Y(n_506) );
BUFx3_ASAP7_75t_L g534 ( .A(n_42), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_44), .B(n_150), .Y(n_272) );
AND2x2_ASAP7_75t_L g170 ( .A(n_46), .B(n_150), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_47), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_49), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_50), .B(n_186), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_51), .A2(n_77), .B1(n_110), .B2(n_111), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_51), .Y(n_110) );
XNOR2x1_ASAP7_75t_L g535 ( .A(n_51), .B(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_52), .A2(n_69), .B1(n_186), .B2(n_551), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_53), .A2(n_72), .B1(n_130), .B2(n_562), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_54), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_55), .A2(n_135), .B(n_160), .C(n_161), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_56), .A2(n_97), .B1(n_549), .B2(n_560), .Y(n_622) );
INVx1_ASAP7_75t_L g126 ( .A(n_57), .Y(n_126) );
AND2x4_ASAP7_75t_L g147 ( .A(n_58), .B(n_148), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_59), .A2(n_60), .B1(n_168), .B2(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_61), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_62), .B(n_150), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_63), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_64), .B(n_168), .Y(n_234) );
INVx1_ASAP7_75t_L g148 ( .A(n_65), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_66), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_67), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_68), .B(n_191), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_70), .B(n_130), .Y(n_129) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_71), .B(n_142), .C(n_182), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_73), .B(n_130), .Y(n_212) );
INVx2_ASAP7_75t_L g137 ( .A(n_74), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_75), .B(n_181), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_76), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_78), .B(n_188), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_79), .A2(n_96), .B1(n_160), .B2(n_168), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_80), .Y(n_588) );
INVx1_ASAP7_75t_L g498 ( .A(n_81), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_82), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_82), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_83), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_85), .A2(n_90), .B1(n_133), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_86), .B(n_181), .Y(n_180) );
NAND2xp33_ASAP7_75t_SL g204 ( .A(n_87), .B(n_187), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_88), .B(n_179), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_89), .B(n_191), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_91), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_92), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g515 ( .A(n_92), .Y(n_515) );
INVx1_ASAP7_75t_L g863 ( .A(n_93), .Y(n_863) );
NAND2xp33_ASAP7_75t_L g616 ( .A(n_94), .B(n_181), .Y(n_616) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_95), .B(n_187), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_98), .B(n_150), .Y(n_149) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_99), .B(n_187), .C(n_199), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_101), .B(n_130), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_102), .B(n_133), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_103), .Y(n_516) );
AOI211xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_517), .B(n_525), .C(n_880), .Y(n_104) );
OAI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_501), .B(n_509), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_493), .B1(n_494), .B2(n_500), .Y(n_107) );
XNOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
XOR2x2_ASAP7_75t_L g500 ( .A(n_109), .B(n_112), .Y(n_500) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g536 ( .A(n_113), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g113 ( .A(n_114), .B(n_388), .Y(n_113) );
NOR2x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_323), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_246), .C(n_296), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_171), .B(n_206), .C(n_223), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g462 ( .A(n_118), .B(n_381), .Y(n_462) );
OR2x2_ASAP7_75t_L g473 ( .A(n_118), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_119), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g364 ( .A(n_119), .B(n_253), .Y(n_364) );
AND2x2_ASAP7_75t_L g485 ( .A(n_119), .B(n_295), .Y(n_485) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_151), .Y(n_119) );
INVx2_ASAP7_75t_L g315 ( .A(n_120), .Y(n_315) );
AND2x2_ASAP7_75t_L g330 ( .A(n_120), .B(n_282), .Y(n_330) );
AND2x2_ASAP7_75t_L g339 ( .A(n_120), .B(n_208), .Y(n_339) );
AND2x2_ASAP7_75t_L g408 ( .A(n_120), .B(n_294), .Y(n_408) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g221 ( .A(n_121), .Y(n_221) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_149), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_122), .A2(n_175), .B(n_190), .Y(n_174) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_122), .A2(n_175), .B(n_190), .Y(n_289) );
OAI21xp33_ASAP7_75t_SL g380 ( .A1(n_122), .A2(n_127), .B(n_149), .Y(n_380) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_123), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_123), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
INVx2_ASAP7_75t_L g245 ( .A(n_124), .Y(n_245) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_125), .Y(n_192) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_138), .B(n_146), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_135), .Y(n_128) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_130), .A2(n_167), .B1(n_168), .B2(n_169), .Y(n_166) );
INVx1_ASAP7_75t_L g551 ( .A(n_130), .Y(n_551) );
INVx1_ASAP7_75t_L g560 ( .A(n_130), .Y(n_560) );
INVx4_ASAP7_75t_L g562 ( .A(n_130), .Y(n_562) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g203 ( .A(n_131), .Y(n_203) );
INVx1_ASAP7_75t_L g242 ( .A(n_131), .Y(n_242) );
INVx1_ASAP7_75t_L g559 ( .A(n_133), .Y(n_559) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_135), .A2(n_202), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_135), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_135), .A2(n_230), .B(n_231), .Y(n_229) );
BUFx4f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx8_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
INVx1_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_143), .Y(n_138) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_176), .B(n_183), .Y(n_175) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_146), .A2(n_197), .B(n_201), .Y(n_196) );
AND2x4_ASAP7_75t_SL g218 ( .A(n_146), .B(n_192), .Y(n_218) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_146), .A2(n_229), .B(n_232), .Y(n_228) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_146), .A2(n_264), .B(n_267), .Y(n_263) );
BUFx10_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx10_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
INVx1_ASAP7_75t_L g586 ( .A(n_147), .Y(n_586) );
AND2x2_ASAP7_75t_L g379 ( .A(n_151), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g222 ( .A(n_152), .B(n_194), .Y(n_222) );
INVx2_ASAP7_75t_L g251 ( .A(n_152), .Y(n_251) );
AOI21x1_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_158), .B(n_170), .Y(n_152) );
NOR2xp67_ASAP7_75t_SL g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx2_ASAP7_75t_L g552 ( .A(n_154), .Y(n_552) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_155), .A2(n_157), .A3(n_237), .B(n_243), .Y(n_236) );
NOR2xp33_ASAP7_75t_SL g565 ( .A(n_155), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_155), .B(n_497), .Y(n_605) );
INVx1_ASAP7_75t_L g546 ( .A(n_156), .Y(n_546) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AO31x2_ASAP7_75t_L g556 ( .A1(n_157), .A2(n_557), .A3(n_564), .B(n_565), .Y(n_556) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_157), .A2(n_570), .A3(n_576), .B(n_577), .Y(n_569) );
AO31x2_ASAP7_75t_L g631 ( .A1(n_157), .A2(n_632), .A3(n_635), .B(n_636), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_164), .Y(n_158) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx2_ASAP7_75t_SL g602 ( .A(n_163), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_165), .A2(n_238), .B1(n_240), .B2(n_241), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_165), .A2(n_240), .B1(n_548), .B2(n_550), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_165), .A2(n_240), .B1(n_571), .B2(n_574), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_165), .A2(n_240), .B1(n_583), .B2(n_584), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_165), .A2(n_240), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx2_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_168), .A2(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g416 ( .A(n_171), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_193), .Y(n_172) );
INVx1_ASAP7_75t_L g436 ( .A(n_173), .Y(n_436) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g274 ( .A(n_174), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g357 ( .A(n_174), .B(n_262), .Y(n_357) );
O2A1O1Ixp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_180), .C(n_182), .Y(n_176) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_198), .B(n_200), .Y(n_197) );
INVx1_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
INVx3_ASAP7_75t_L g549 ( .A(n_181), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_233), .B(n_234), .Y(n_232) );
INVx6_ASAP7_75t_L g240 ( .A(n_182), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g611 ( .A1(n_182), .A2(n_562), .B(n_612), .C(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_188), .Y(n_183) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g572 ( .A(n_187), .Y(n_572) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_189), .A2(n_215), .B1(n_216), .B2(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g635 ( .A(n_191), .Y(n_635) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_SL g195 ( .A(n_192), .Y(n_195) );
INVx2_ASAP7_75t_L g227 ( .A(n_192), .Y(n_227) );
BUFx3_ASAP7_75t_L g576 ( .A(n_192), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_192), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g609 ( .A(n_192), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_192), .B(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_192), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g283 ( .A(n_193), .B(n_221), .Y(n_283) );
INVxp67_ASAP7_75t_L g432 ( .A(n_193), .Y(n_432) );
OR2x2_ASAP7_75t_L g474 ( .A(n_193), .B(n_208), .Y(n_474) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_205), .Y(n_194) );
INVx1_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
INVx1_ASAP7_75t_SL g563 ( .A(n_199), .Y(n_563) );
INVx1_ASAP7_75t_L g604 ( .A(n_199), .Y(n_604) );
INVx1_ASAP7_75t_L g573 ( .A(n_203), .Y(n_573) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
INVx1_ASAP7_75t_L g329 ( .A(n_207), .Y(n_329) );
AND2x2_ASAP7_75t_L g483 ( .A(n_207), .B(n_379), .Y(n_483) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g254 ( .A(n_208), .Y(n_254) );
INVx4_ASAP7_75t_L g294 ( .A(n_208), .Y(n_294) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_218), .Y(n_210) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
AND2x2_ASAP7_75t_L g310 ( .A(n_220), .B(n_293), .Y(n_310) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g347 ( .A(n_221), .B(n_295), .Y(n_347) );
INVx2_ASAP7_75t_L g313 ( .A(n_222), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_222), .B(n_318), .Y(n_481) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_225), .B(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g466 ( .A(n_225), .Y(n_466) );
AND2x2_ASAP7_75t_L g480 ( .A(n_225), .B(n_302), .Y(n_480) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_236), .Y(n_225) );
INVx1_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
AND2x2_ASAP7_75t_L g415 ( .A(n_226), .B(n_322), .Y(n_415) );
OR2x2_ASAP7_75t_L g452 ( .A(n_226), .B(n_236), .Y(n_452) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_235), .Y(n_226) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_227), .A2(n_263), .B(n_272), .Y(n_262) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_227), .A2(n_263), .B(n_272), .Y(n_275) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_227), .A2(n_228), .B(n_235), .Y(n_278) );
AND2x2_ASAP7_75t_L g261 ( .A(n_236), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g276 ( .A(n_236), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
OR2x2_ASAP7_75t_L g335 ( .A(n_236), .B(n_275), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_236), .B(n_275), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_240), .A2(n_558), .B1(n_561), .B2(n_563), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_240), .A2(n_601), .B1(n_603), .B2(n_604), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_240), .A2(n_615), .B(n_616), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_240), .A2(n_563), .B1(n_622), .B2(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g575 ( .A(n_242), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
BUFx2_ASAP7_75t_L g564 ( .A(n_245), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_256), .B(n_279), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI31xp33_ASAP7_75t_L g325 ( .A1(n_248), .A2(n_326), .A3(n_328), .B(n_331), .Y(n_325) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
AND2x2_ASAP7_75t_L g338 ( .A(n_249), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g348 ( .A(n_250), .Y(n_348) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_250), .Y(n_354) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
AND2x2_ASAP7_75t_L g311 ( .A(n_251), .B(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g361 ( .A(n_251), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_252), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g386 ( .A(n_253), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g435 ( .A(n_253), .B(n_436), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g490 ( .A1(n_253), .A2(n_320), .A3(n_330), .B1(n_357), .B2(n_466), .B3(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
INVx1_ASAP7_75t_L g382 ( .A(n_255), .Y(n_382) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_273), .Y(n_257) );
INVx2_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
AND2x2_ASAP7_75t_L g371 ( .A(n_258), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx1_ASAP7_75t_L g333 ( .A(n_259), .Y(n_333) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g401 ( .A(n_260), .B(n_288), .Y(n_401) );
AND2x2_ASAP7_75t_L g351 ( .A(n_261), .B(n_345), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_261), .B(n_369), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_261), .B(n_401), .Y(n_450) );
AND2x2_ASAP7_75t_L g287 ( .A(n_262), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_301), .Y(n_306) );
INVx1_ASAP7_75t_L g321 ( .A(n_262), .Y(n_321) );
AOI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_271), .Y(n_267) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g376 ( .A(n_274), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_274), .B(n_469), .Y(n_471) );
AND2x2_ASAP7_75t_L g484 ( .A(n_274), .B(n_300), .Y(n_484) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_288), .Y(n_302) );
INVx2_ASAP7_75t_L g284 ( .A(n_276), .Y(n_284) );
AND2x2_ASAP7_75t_L g398 ( .A(n_276), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g457 ( .A(n_276), .B(n_369), .Y(n_457) );
BUFx2_ASAP7_75t_L g439 ( .A(n_277), .Y(n_439) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx3_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
OAI32xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .A3(n_285), .B1(n_290), .B2(n_291), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g387 ( .A(n_282), .Y(n_387) );
AND2x2_ASAP7_75t_L g417 ( .A(n_282), .B(n_339), .Y(n_417) );
AND2x2_ASAP7_75t_L g359 ( .A(n_283), .B(n_360), .Y(n_359) );
AND3x2_ASAP7_75t_L g366 ( .A(n_283), .B(n_293), .C(n_361), .Y(n_366) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_286), .A2(n_308), .B1(n_317), .B2(n_319), .Y(n_316) );
OAI322xp33_ASAP7_75t_L g464 ( .A1(n_286), .A2(n_385), .A3(n_465), .B1(n_466), .B2(n_467), .C1(n_468), .C2(n_471), .Y(n_464) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g486 ( .A(n_287), .B(n_469), .Y(n_486) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_288), .Y(n_305) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_288), .Y(n_345) );
BUFx3_ASAP7_75t_L g369 ( .A(n_288), .Y(n_369) );
INVx1_ASAP7_75t_L g395 ( .A(n_288), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_288), .Y(n_399) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g353 ( .A(n_292), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g404 ( .A(n_293), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_293), .B(n_361), .Y(n_455) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_294), .B(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
AND2x2_ASAP7_75t_L g360 ( .A(n_294), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g381 ( .A(n_294), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_295), .B(n_408), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_303), .B(n_307), .C(n_316), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI31xp33_ASAP7_75t_L g458 ( .A1(n_298), .A2(n_459), .A3(n_461), .B(n_462), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
AND2x4_ASAP7_75t_L g411 ( .A(n_299), .B(n_320), .Y(n_411) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_301), .B(n_321), .Y(n_427) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g467 ( .A(n_310), .Y(n_467) );
AND2x2_ASAP7_75t_L g327 ( .A(n_311), .B(n_318), .Y(n_327) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_312), .A2(n_397), .B1(n_400), .B2(n_402), .Y(n_396) );
OR2x6_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g454 ( .A(n_315), .Y(n_454) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g424 ( .A(n_320), .B(n_369), .Y(n_424) );
INVx2_ASAP7_75t_L g470 ( .A(n_320), .Y(n_470) );
AND2x4_ASAP7_75t_L g478 ( .A(n_320), .B(n_399), .Y(n_478) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_340), .C(n_370), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_336), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_327), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g391 ( .A(n_329), .B(n_346), .Y(n_391) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_332), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g422 ( .A(n_334), .B(n_401), .Y(n_422) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_335), .Y(n_342) );
INVx1_ASAP7_75t_L g460 ( .A(n_335), .Y(n_460) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g489 ( .A(n_338), .Y(n_489) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_346), .B(n_349), .C(n_362), .Y(n_340) );
NOR3x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .C(n_344), .Y(n_341) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_344), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2x1p5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B1(n_355), .B2(n_358), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g443 ( .A(n_354), .Y(n_443) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g438 ( .A(n_357), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g492 ( .A(n_360), .Y(n_492) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_367), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g373 ( .A(n_369), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_427), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B(n_375), .Y(n_370) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_373), .B(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_383), .B2(n_385), .Y(n_375) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g403 ( .A(n_379), .B(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
INVx1_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_444), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_390), .B(n_405), .C(n_418), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g451 ( .A(n_394), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_403), .B(n_431), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_412), .B2(n_416), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_413), .A2(n_434), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_429), .B1(n_433), .B2(n_441), .Y(n_418) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_423), .Y(n_419) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g469 ( .A(n_439), .Y(n_469) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_463), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .C(n_458), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_453), .C(n_456), .Y(n_449) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_472), .C(n_487), .Y(n_463) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .B1(n_479), .B2(n_481), .C(n_482), .Y(n_472) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_482) );
OAI21xp33_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_497), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
CKINVDCx8_ASAP7_75t_R g877 ( .A(n_503), .Y(n_877) );
INVx3_ASAP7_75t_L g885 ( .A(n_503), .Y(n_885) );
AND2x6_ASAP7_75t_SL g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_506), .Y(n_513) );
AND3x2_ASAP7_75t_L g512 ( .A(n_507), .B(n_513), .C(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_508), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_511), .B(n_516), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g531 ( .A(n_515), .Y(n_531) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
BUFx2_ASAP7_75t_L g879 ( .A(n_519), .Y(n_879) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_520), .B(n_885), .Y(n_884) );
OR2x4_ASAP7_75t_L g883 ( .A(n_521), .B(n_884), .Y(n_883) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g878 ( .A(n_523), .B(n_879), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_867), .B(n_874), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_857), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_535), .B1(n_537), .B2(n_854), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g868 ( .A(n_529), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NOR2x1_ASAP7_75t_R g855 ( .A(n_530), .B(n_856), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g873 ( .A(n_531), .B(n_533), .Y(n_873) );
INVxp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g856 ( .A(n_533), .Y(n_856) );
A2O1A1O1Ixp25_ASAP7_75t_SL g867 ( .A1(n_535), .A2(n_858), .B(n_868), .C(n_869), .D(n_870), .Y(n_867) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_538), .B(n_854), .Y(n_869) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_763), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_702), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_653), .C(n_672), .D(n_683), .Y(n_540) );
O2A1O1Ixp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_589), .B(n_596), .C(n_626), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_567), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_543), .B(n_718), .C(n_719), .Y(n_717) );
AND2x2_ASAP7_75t_L g799 ( .A(n_543), .B(n_681), .Y(n_799) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x2_ASAP7_75t_L g643 ( .A(n_544), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g661 ( .A(n_544), .B(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g678 ( .A(n_544), .Y(n_678) );
AND2x2_ASAP7_75t_L g723 ( .A(n_544), .B(n_569), .Y(n_723) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
AND2x4_ASAP7_75t_L g671 ( .A(n_545), .B(n_662), .Y(n_671) );
AO31x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .A3(n_552), .B(n_553), .Y(n_545) );
AO31x2_ASAP7_75t_L g620 ( .A1(n_546), .A2(n_564), .A3(n_621), .B(n_624), .Y(n_620) );
AO31x2_ASAP7_75t_L g581 ( .A1(n_552), .A2(n_582), .A3(n_585), .B(n_587), .Y(n_581) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g646 ( .A(n_555), .B(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_555), .Y(n_669) );
INVx1_ASAP7_75t_L g680 ( .A(n_555), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_555), .B(n_579), .Y(n_689) );
INVx2_ASAP7_75t_L g696 ( .A(n_555), .Y(n_696) );
INVx4_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g641 ( .A(n_556), .B(n_569), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_556), .B(n_648), .Y(n_714) );
AND2x2_ASAP7_75t_L g722 ( .A(n_556), .B(n_581), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_556), .B(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g775 ( .A(n_556), .Y(n_775) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g791 ( .A(n_568), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_579), .Y(n_568) );
INVx1_ASAP7_75t_L g595 ( .A(n_569), .Y(n_595) );
INVx1_ASAP7_75t_L g648 ( .A(n_569), .Y(n_648) );
INVx2_ASAP7_75t_L g682 ( .A(n_569), .Y(n_682) );
OR2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_581), .Y(n_686) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_569), .Y(n_735) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_576), .A2(n_585), .A3(n_600), .B(n_605), .Y(n_599) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g708 ( .A(n_580), .B(n_593), .Y(n_708) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_581), .Y(n_644) );
INVx2_ASAP7_75t_L g662 ( .A(n_581), .Y(n_662) );
AND2x4_ASAP7_75t_L g681 ( .A(n_581), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g769 ( .A(n_581), .Y(n_769) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g617 ( .A(n_586), .Y(n_617) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g687 ( .A(n_592), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_592), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g750 ( .A(n_593), .Y(n_750) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_606), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_598), .B(n_607), .Y(n_700) );
INVx1_ASAP7_75t_L g798 ( .A(n_598), .Y(n_798) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g638 ( .A(n_599), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g652 ( .A(n_599), .B(n_631), .Y(n_652) );
AND2x4_ASAP7_75t_L g675 ( .A(n_599), .B(n_619), .Y(n_675) );
INVx2_ASAP7_75t_L g692 ( .A(n_599), .Y(n_692) );
AND2x2_ASAP7_75t_L g718 ( .A(n_599), .B(n_620), .Y(n_718) );
INVx1_ASAP7_75t_L g783 ( .A(n_599), .Y(n_783) );
AND2x2_ASAP7_75t_L g743 ( .A(n_606), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_619), .Y(n_606) );
AND2x2_ASAP7_75t_L g709 ( .A(n_607), .B(n_666), .Y(n_709) );
AND2x4_ASAP7_75t_L g725 ( .A(n_607), .B(n_692), .Y(n_725) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g719 ( .A(n_608), .Y(n_719) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_618), .Y(n_608) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_609), .A2(n_610), .B(n_618), .Y(n_640) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_614), .B(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g651 ( .A(n_619), .Y(n_651) );
INVx3_ASAP7_75t_L g657 ( .A(n_619), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_619), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_619), .B(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g691 ( .A(n_620), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g815 ( .A(n_620), .Y(n_815) );
OAI33xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_641), .A3(n_642), .B1(n_643), .B2(n_645), .B3(n_649), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_638), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g749 ( .A(n_630), .B(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g658 ( .A(n_631), .B(n_640), .Y(n_658) );
INVx2_ASAP7_75t_L g666 ( .A(n_631), .Y(n_666) );
INVx1_ASAP7_75t_L g674 ( .A(n_631), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_638), .A2(n_694), .B1(n_697), .B2(n_701), .Y(n_693) );
OR2x2_ASAP7_75t_L g833 ( .A(n_638), .B(n_651), .Y(n_833) );
AND2x4_ASAP7_75t_L g737 ( .A(n_639), .B(n_699), .Y(n_737) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_640), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_641), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g701 ( .A(n_641), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_641), .B(n_677), .Y(n_779) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g752 ( .A(n_643), .Y(n_752) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g810 ( .A(n_646), .B(n_678), .Y(n_810) );
NAND2x1_ASAP7_75t_L g828 ( .A(n_646), .B(n_677), .Y(n_828) );
AND2x2_ASAP7_75t_L g852 ( .A(n_646), .B(n_671), .Y(n_852) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g842 ( .A(n_650), .B(n_719), .Y(n_842) );
NOR2x1p5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g776 ( .A(n_651), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g744 ( .A(n_652), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_659), .B1(n_663), .B2(n_667), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
AND2x2_ASAP7_75t_L g751 ( .A(n_656), .B(n_719), .Y(n_751) );
AND2x2_ASAP7_75t_L g788 ( .A(n_656), .B(n_737), .Y(n_788) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g663 ( .A(n_657), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_657), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g829 ( .A(n_657), .B(n_658), .Y(n_829) );
AND2x2_ASAP7_75t_L g690 ( .A(n_658), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g809 ( .A(n_658), .B(n_675), .Y(n_809) );
AND2x2_ASAP7_75t_L g853 ( .A(n_658), .B(n_718), .Y(n_853) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_663), .A2(n_788), .B1(n_789), .B2(n_792), .C1(n_794), .C2(n_795), .Y(n_787) );
AND2x2_ASAP7_75t_L g710 ( .A(n_664), .B(n_678), .Y(n_710) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g741 ( .A(n_665), .Y(n_741) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_665), .Y(n_786) );
INVx2_ASAP7_75t_L g699 ( .A(n_666), .Y(n_699) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g756 ( .A(n_669), .Y(n_756) );
INVx2_ASAP7_75t_L g762 ( .A(n_670), .Y(n_762) );
INVx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g746 ( .A(n_671), .B(n_735), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x4_ASAP7_75t_L g777 ( .A(n_674), .B(n_725), .Y(n_777) );
INVx2_ASAP7_75t_L g824 ( .A(n_674), .Y(n_824) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx4_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g767 ( .A(n_678), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g801 ( .A(n_678), .B(n_686), .Y(n_801) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g706 ( .A(n_680), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_681), .B(n_771), .Y(n_770) );
AND2x4_ASAP7_75t_L g813 ( .A(n_681), .B(n_729), .Y(n_813) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_688), .B(n_690), .C(n_693), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OR2x2_ASAP7_75t_L g694 ( .A(n_686), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g730 ( .A(n_686), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_687), .B(n_722), .Y(n_826) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g802 ( .A(n_689), .B(n_771), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_691), .B(n_741), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_691), .A2(n_707), .B1(n_749), .B2(n_751), .Y(n_748) );
AND2x2_ASAP7_75t_L g754 ( .A(n_691), .B(n_719), .Y(n_754) );
AND2x2_ASAP7_75t_L g823 ( .A(n_691), .B(n_824), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_L g816 ( .A1(n_694), .A2(n_796), .B(n_817), .C(n_820), .Y(n_816) );
INVx2_ASAP7_75t_L g729 ( .A(n_696), .Y(n_729) );
OR2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g807 ( .A(n_699), .Y(n_807) );
INVx1_ASAP7_75t_L g732 ( .A(n_700), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_701), .A2(n_748), .B1(n_752), .B2(n_753), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_715), .C(n_738), .Y(n_702) );
AO22x1_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_708), .Y(n_841) );
OR2x2_ASAP7_75t_L g848 ( .A(n_708), .B(n_729), .Y(n_848) );
AND2x2_ASAP7_75t_L g760 ( .A(n_709), .B(n_718), .Y(n_760) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g836 ( .A(n_714), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .C(n_726), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g758 ( .A(n_718), .Y(n_758) );
AND2x4_ASAP7_75t_SL g794 ( .A(n_718), .B(n_737), .Y(n_794) );
INVx1_ASAP7_75t_SL g805 ( .A(n_718), .Y(n_805) );
OR2x2_ASAP7_75t_L g757 ( .A(n_719), .B(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AND2x4_ASAP7_75t_L g734 ( .A(n_722), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g792 ( .A(n_723), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g814 ( .A(n_725), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g839 ( .A(n_725), .B(n_819), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .B1(n_733), .B2(n_736), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x4_ASAP7_75t_L g774 ( .A(n_730), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g796 ( .A(n_730), .Y(n_796) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g851 ( .A(n_734), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_747), .C(n_755), .Y(n_738) );
AOI21xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .B(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g820 ( .A(n_741), .Y(n_820) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI222xp33_ASAP7_75t_L g843 ( .A1(n_746), .A2(n_844), .B1(n_847), .B2(n_849), .C1(n_851), .C2(n_853), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_749), .B(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g772 ( .A(n_750), .Y(n_772) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_759), .C(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_821), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_765), .B(n_787), .C(n_797), .D(n_808), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_776), .B1(n_778), .B2(n_780), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .C(n_773), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_767), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g793 ( .A(n_769), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_771), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g818 ( .A(n_783), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g832 ( .A(n_784), .Y(n_832) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_785), .Y(n_850) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g845 ( .A(n_794), .Y(n_845) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_800), .C(n_806), .Y(n_797) );
AOI21xp33_ASAP7_75t_SL g800 ( .A1(n_801), .A2(n_802), .B(n_803), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_801), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_811), .B2(n_814), .C(n_816), .Y(n_808) );
INVx1_ASAP7_75t_L g846 ( .A(n_809), .Y(n_846) );
AOI31xp33_ASAP7_75t_L g830 ( .A1(n_812), .A2(n_831), .A3(n_832), .B(n_833), .Y(n_830) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g819 ( .A(n_815), .Y(n_819) );
INVxp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_834), .C(n_843), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_825), .B1(n_827), .B2(n_829), .C(n_830), .Y(n_822) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_SL g831 ( .A(n_829), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_837), .B1(n_840), .B2(n_842), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g866 ( .A(n_859), .Y(n_866) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx6_ASAP7_75t_SL g881 ( .A(n_882), .Y(n_881) );
BUFx10_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
endmodule