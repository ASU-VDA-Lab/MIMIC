module fake_netlist_6_1727_n_1307 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1307);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1307;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1287;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_934;
wire n_482;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_216),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_42),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_19),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_24),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_192),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_181),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_139),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_111),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_21),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_209),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_24),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_175),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_120),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_86),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_141),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_171),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_164),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_107),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_122),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_189),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_128),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_146),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_94),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_153),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_261),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_109),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_132),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_200),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_170),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_129),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_117),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_279),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_65),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_215),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

BUFx8_ASAP7_75t_SL g341 ( 
.A(n_235),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_93),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_5),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_248),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_218),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_151),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_143),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_96),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_71),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_160),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_110),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_223),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_179),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_145),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_89),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_245),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_242),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_174),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_9),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_56),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_8),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_246),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_152),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_183),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_203),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_264),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_221),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_59),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_255),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_55),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_105),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_95),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_60),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_155),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_172),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_101),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_259),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_256),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_51),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_21),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_44),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_113),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_60),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_65),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_249),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_44),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_29),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_234),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_186),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_48),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_284),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_138),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_76),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_72),
.Y(n_399)
);

INVxp33_ASAP7_75t_R g400 ( 
.A(n_82),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_281),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_104),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_159),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_212),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_29),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_220),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_4),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_123),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_150),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_79),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_22),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_52),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_278),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_133),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_147),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_12),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_106),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_47),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_90),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_225),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_140),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_54),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_136),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_274),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_197),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_14),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_195),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_37),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_57),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_165),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_124),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_262),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_6),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_4),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_30),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_73),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_214),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_230),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_280),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_10),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_239),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_82),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_208),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_213),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_266),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_134),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_62),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_38),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_228),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_268),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_282),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_229),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_227),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_196),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_92),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_112),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_288),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_258),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_137),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_3),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_126),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_31),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_75),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_265),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_257),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_292),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_201),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_285),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_118),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_202),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_217),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_286),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_63),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_190),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_219),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_39),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_297),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_247),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_226),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_222),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_254),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_127),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_161),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_116),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_27),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_193),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_303),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_429),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_401),
.B(n_0),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_303),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_422),
.B(n_0),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_378),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_303),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_366),
.B(n_1),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_303),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_339),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_378),
.B(n_2),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_366),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_422),
.B(n_2),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_339),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_345),
.B(n_3),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_339),
.B(n_85),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_339),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_349),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_378),
.B(n_5),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_349),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_349),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_429),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_419),
.B(n_6),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_378),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_378),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_298),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_7),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_458),
.B(n_7),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_328),
.B(n_10),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_458),
.B(n_11),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_345),
.B(n_11),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_350),
.B(n_12),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_350),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_306),
.B(n_13),
.Y(n_526)
);

INVx6_ASAP7_75t_L g527 ( 
.A(n_344),
.Y(n_527)
);

BUFx8_ASAP7_75t_SL g528 ( 
.A(n_341),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_382),
.B(n_13),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_406),
.B(n_14),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_382),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_424),
.B(n_15),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_409),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_463),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_384),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_424),
.B(n_15),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_430),
.B(n_16),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_431),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_481),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_438),
.B(n_17),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_438),
.B(n_17),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_455),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_445),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_307),
.Y(n_549)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_464),
.B(n_18),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_19),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_343),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_299),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_300),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_392),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_308),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_317),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_321),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_323),
.B(n_20),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_392),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_309),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_325),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_368),
.B(n_22),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_369),
.B(n_23),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_362),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_334),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_375),
.B(n_23),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_335),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_338),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_363),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_372),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_340),
.B(n_25),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_312),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_347),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_352),
.B(n_25),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_354),
.Y(n_576)
);

BUFx12f_ASAP7_75t_L g577 ( 
.A(n_337),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_364),
.B(n_26),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_367),
.B(n_27),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_407),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_381),
.B(n_28),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_411),
.B(n_435),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_374),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_411),
.B(n_28),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_390),
.B(n_30),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_473),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_351),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_377),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_414),
.B(n_415),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_365),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_302),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_304),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_373),
.B(n_32),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_420),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_385),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_386),
.B(n_33),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_432),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_400),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_443),
.B(n_444),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_449),
.B(n_33),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_450),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_391),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_398),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_305),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_388),
.Y(n_608)
);

BUFx8_ASAP7_75t_SL g609 ( 
.A(n_389),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_457),
.B(n_459),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_461),
.B(n_34),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_466),
.B(n_35),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_395),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_467),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_490),
.A2(n_389),
.B1(n_399),
.B2(n_301),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_567),
.A2(n_412),
.B1(n_416),
.B2(n_410),
.Y(n_616)
);

AO22x2_ASAP7_75t_L g617 ( 
.A1(n_495),
.A2(n_405),
.B1(n_447),
.B2(n_418),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_503),
.B(n_469),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_523),
.A2(n_371),
.B1(n_376),
.B2(n_360),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_527),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_495),
.A2(n_483),
.B1(n_477),
.B2(n_453),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_556),
.B(n_441),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_527),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_311),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_525),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_551),
.A2(n_563),
.B1(n_564),
.B2(n_567),
.Y(n_629)
);

AO22x2_ASAP7_75t_L g630 ( 
.A1(n_512),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_489),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_556),
.B(n_313),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_492),
.A2(n_425),
.B1(n_360),
.B2(n_314),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_515),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_489),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_526),
.A2(n_425),
.B1(n_428),
.B2(n_426),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_510),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_510),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_549),
.B(n_592),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_487),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_545),
.A2(n_434),
.B1(n_436),
.B2(n_433),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_531),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_538),
.A2(n_442),
.B1(n_448),
.B2(n_440),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_491),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_577),
.B(n_460),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_491),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_315),
.Y(n_648)
);

AND2x2_ASAP7_75t_SL g649 ( 
.A(n_501),
.B(n_310),
.Y(n_649)
);

BUFx10_ASAP7_75t_L g650 ( 
.A(n_594),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_595),
.A2(n_333),
.B1(n_348),
.B2(n_320),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_491),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_573),
.B(n_316),
.Y(n_653)
);

OA22x2_ASAP7_75t_L g654 ( 
.A1(n_583),
.A2(n_476),
.B1(n_485),
.B2(n_462),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_588),
.A2(n_319),
.B1(n_322),
.B2(n_318),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_500),
.B(n_324),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_498),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_498),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_512),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_532),
.B(n_326),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_600),
.A2(n_329),
.B1(n_330),
.B2(n_327),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_498),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_546),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_532),
.B(n_331),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_505),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_528),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_505),
.Y(n_667)
);

AO22x2_ASAP7_75t_L g668 ( 
.A1(n_517),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_332),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_607),
.B(n_336),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_545),
.A2(n_346),
.B1(n_353),
.B2(n_342),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_519),
.A2(n_356),
.B1(n_357),
.B2(n_355),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_534),
.A2(n_359),
.B1(n_361),
.B2(n_358),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_504),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_505),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_506),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_530),
.A2(n_379),
.B1(n_380),
.B2(n_370),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_534),
.B(n_383),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_572),
.A2(n_393),
.B1(n_394),
.B2(n_387),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g681 ( 
.A(n_517),
.B(n_40),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_396),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_543),
.B(n_486),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_534),
.A2(n_403),
.B1(n_404),
.B2(n_397),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_506),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_539),
.B(n_408),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_518),
.B(n_413),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_506),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_539),
.B(n_540),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_518),
.B(n_417),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_540),
.B(n_421),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_520),
.A2(n_454),
.B1(n_482),
.B2(n_480),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_508),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_520),
.A2(n_484),
.B1(n_478),
.B2(n_475),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_544),
.A2(n_451),
.B1(n_472),
.B2(n_471),
.Y(n_695)
);

AO22x2_ASAP7_75t_L g696 ( 
.A1(n_524),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_508),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_600),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_SL g699 ( 
.A1(n_600),
.A2(n_474),
.B1(n_470),
.B2(n_465),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_598),
.B(n_584),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_SL g701 ( 
.A(n_524),
.B(n_423),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_508),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_673),
.B(n_535),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_657),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_700),
.B(n_513),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_677),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_677),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_642),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_649),
.B(n_529),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_685),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_685),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_693),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_634),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_693),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_639),
.B(n_541),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_700),
.A2(n_591),
.B(n_601),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_675),
.B(n_550),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_702),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_663),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_663),
.B(n_541),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_621),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_698),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_620),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_656),
.B(n_535),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_625),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_618),
.B(n_514),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_618),
.A2(n_701),
.B(n_643),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_640),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_695),
.B(n_542),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_652),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_658),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_665),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_675),
.B(n_550),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_667),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_651),
.B(n_542),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_676),
.Y(n_741)
);

INVxp33_ASAP7_75t_L g742 ( 
.A(n_615),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_687),
.B(n_601),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_688),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_648),
.B(n_542),
.Y(n_745)
);

XOR2xp5_ASAP7_75t_L g746 ( 
.A(n_633),
.B(n_427),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_689),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_697),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_619),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_529),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_629),
.B(n_552),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_642),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_642),
.Y(n_754)
);

XOR2xp5_ASAP7_75t_L g755 ( 
.A(n_655),
.B(n_437),
.Y(n_755)
);

BUFx5_ASAP7_75t_L g756 ( 
.A(n_637),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_645),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_653),
.B(n_552),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_645),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_645),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_690),
.B(n_493),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_623),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_631),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_635),
.Y(n_764)
);

INVxp33_ASAP7_75t_L g765 ( 
.A(n_636),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_626),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_638),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_617),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_660),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_617),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_681),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_671),
.B(n_552),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_690),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_627),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_632),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_664),
.B(n_497),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_669),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_679),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_686),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_650),
.B(n_605),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_624),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_624),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_641),
.B(n_497),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_682),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_661),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_704),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_767),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_756),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_768),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_720),
.Y(n_793)
);

AND2x2_ASAP7_75t_SL g794 ( 
.A(n_712),
.B(n_533),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_777),
.B(n_670),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_777),
.B(n_692),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_769),
.B(n_533),
.Y(n_797)
);

BUFx5_ASAP7_75t_L g798 ( 
.A(n_750),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_761),
.B(n_694),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_725),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_749),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_752),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_761),
.B(n_696),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_727),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_781),
.B(n_559),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_711),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_750),
.B(n_672),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_730),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_774),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_727),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_630),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_762),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_707),
.A2(n_680),
.B(n_507),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_707),
.B(n_659),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_773),
.B(n_537),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_720),
.B(n_678),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_738),
.B(n_616),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_756),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_763),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_750),
.B(n_683),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_659),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_764),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_751),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_711),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_756),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_776),
.B(n_668),
.Y(n_826)
);

AND2x2_ASAP7_75t_SL g827 ( 
.A(n_773),
.B(n_537),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_750),
.B(n_786),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_779),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_743),
.B(n_778),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_743),
.B(n_668),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_780),
.B(n_610),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_703),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_785),
.B(n_559),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_719),
.A2(n_499),
.B(n_602),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_766),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_719),
.A2(n_499),
.B(n_575),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_705),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_706),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_726),
.B(n_646),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_770),
.B(n_578),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_771),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_728),
.B(n_674),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_756),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_731),
.B(n_578),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_716),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_785),
.B(n_579),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_758),
.B(n_751),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_747),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_733),
.B(n_581),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_722),
.B(n_684),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_723),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_726),
.B(n_646),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_R g854 ( 
.A(n_784),
.B(n_605),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_740),
.B(n_644),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_754),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_772),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_783),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_708),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_782),
.B(n_610),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_745),
.B(n_586),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_732),
.B(n_611),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_709),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_759),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_711),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_710),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_753),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_713),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_714),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_715),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_757),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_717),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_724),
.B(n_691),
.Y(n_873)
);

INVxp33_ASAP7_75t_L g874 ( 
.A(n_746),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_760),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_721),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_734),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_801),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_829),
.Y(n_879)
);

INVx8_ASAP7_75t_L g880 ( 
.A(n_797),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_795),
.B(n_729),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_800),
.B(n_772),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_793),
.B(n_735),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_788),
.B(n_736),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_788),
.B(n_737),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_801),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_789),
.B(n_739),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_806),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_823),
.B(n_765),
.Y(n_889)
);

BUFx12f_ASAP7_75t_L g890 ( 
.A(n_846),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_789),
.B(n_741),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_857),
.B(n_742),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_831),
.B(n_666),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_808),
.B(n_744),
.Y(n_894)
);

BUFx8_ASAP7_75t_SL g895 ( 
.A(n_836),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_863),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_849),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_831),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_801),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_858),
.Y(n_900)
);

NAND2x1_ASAP7_75t_SL g901 ( 
.A(n_845),
.B(n_611),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_845),
.B(n_612),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_848),
.B(n_755),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_809),
.B(n_748),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_867),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_806),
.Y(n_906)
);

BUFx8_ASAP7_75t_SL g907 ( 
.A(n_849),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_SL g908 ( 
.A(n_794),
.B(n_793),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_806),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_802),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_867),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_806),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_810),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_830),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_804),
.B(n_699),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_809),
.B(n_787),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_830),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_804),
.B(n_598),
.Y(n_918)
);

BUFx12f_ASAP7_75t_L g919 ( 
.A(n_840),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_865),
.B(n_589),
.Y(n_920)
);

INVx6_ASAP7_75t_L g921 ( 
.A(n_853),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_865),
.B(n_589),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_790),
.B(n_553),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_SL g924 ( 
.A(n_794),
.B(n_609),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_852),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_863),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_866),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_792),
.B(n_554),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_821),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_824),
.B(n_597),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_866),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_842),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_814),
.B(n_584),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_868),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_834),
.B(n_531),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_869),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_805),
.B(n_561),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_805),
.B(n_871),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_832),
.B(n_605),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_832),
.B(n_606),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_565),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_847),
.B(n_547),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_796),
.B(n_582),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_841),
.B(n_582),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_871),
.B(n_570),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_878),
.Y(n_946)
);

INVx8_ASAP7_75t_L g947 ( 
.A(n_880),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_907),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_888),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_882),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_895),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_889),
.A2(n_850),
.B1(n_827),
.B2(n_815),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_892),
.B(n_803),
.Y(n_953)
);

CKINVDCx6p67_ASAP7_75t_R g954 ( 
.A(n_890),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_897),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_925),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_898),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_878),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_888),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_931),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_888),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_896),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_926),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_906),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_886),
.Y(n_965)
);

CKINVDCx6p67_ASAP7_75t_R g966 ( 
.A(n_893),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_893),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_921),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_906),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_919),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_938),
.B(n_812),
.Y(n_971)
);

BUFx2_ASAP7_75t_SL g972 ( 
.A(n_914),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_917),
.Y(n_973)
);

CKINVDCx6p67_ASAP7_75t_R g974 ( 
.A(n_915),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_927),
.Y(n_975)
);

INVx5_ASAP7_75t_SL g976 ( 
.A(n_933),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_943),
.B(n_799),
.Y(n_977)
);

INVx8_ASAP7_75t_L g978 ( 
.A(n_880),
.Y(n_978)
);

INVx6_ASAP7_75t_L g979 ( 
.A(n_929),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_886),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_900),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_881),
.B(n_815),
.Y(n_982)
);

INVx8_ASAP7_75t_L g983 ( 
.A(n_912),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_934),
.Y(n_984)
);

CKINVDCx6p67_ASAP7_75t_R g985 ( 
.A(n_915),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_938),
.B(n_819),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_912),
.Y(n_987)
);

BUFx2_ASAP7_75t_SL g988 ( 
.A(n_916),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_932),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_904),
.B(n_822),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_879),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_945),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_913),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_904),
.B(n_833),
.Y(n_994)
);

BUFx4_ASAP7_75t_SL g995 ( 
.A(n_933),
.Y(n_995)
);

BUFx2_ASAP7_75t_SL g996 ( 
.A(n_912),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_899),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_909),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_918),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_905),
.Y(n_1000)
);

BUFx2_ASAP7_75t_SL g1001 ( 
.A(n_909),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_905),
.B(n_802),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_920),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_922),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_918),
.Y(n_1005)
);

BUFx2_ASAP7_75t_SL g1006 ( 
.A(n_937),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_937),
.Y(n_1007)
);

BUFx4_ASAP7_75t_SL g1008 ( 
.A(n_944),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_970),
.Y(n_1009)
);

OAI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_952),
.A2(n_977),
.B1(n_982),
.B2(n_908),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_983),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_983),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_955),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_SL g1014 ( 
.A1(n_988),
.A2(n_924),
.B1(n_850),
.B2(n_903),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_946),
.Y(n_1015)
);

CKINVDCx6p67_ASAP7_75t_R g1016 ( 
.A(n_948),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_946),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_953),
.A2(n_843),
.B1(n_835),
.B2(n_837),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_958),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_960),
.A2(n_813),
.B1(n_855),
.B2(n_936),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_956),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_983),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_962),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_963),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_975),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_984),
.A2(n_855),
.B1(n_816),
.B2(n_817),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_958),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_974),
.A2(n_816),
.B1(n_817),
.B2(n_862),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_954),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_947),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_974),
.A2(n_862),
.B1(n_942),
.B2(n_935),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_950),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_968),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_947),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_965),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_968),
.Y(n_1036)
);

BUFx10_ASAP7_75t_L g1037 ( 
.A(n_979),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_965),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_993),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_985),
.A2(n_851),
.B1(n_894),
.B2(n_861),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_976),
.A2(n_876),
.B1(n_870),
.B2(n_923),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_976),
.A2(n_876),
.B1(n_870),
.B2(n_923),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_980),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_997),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_997),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_979),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_993),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_994),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_954),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_999),
.A2(n_928),
.B1(n_826),
.B2(n_839),
.Y(n_1050)
);

INVx6_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

CKINVDCx6p67_ASAP7_75t_R g1052 ( 
.A(n_948),
.Y(n_1052)
);

BUFx4_ASAP7_75t_R g1053 ( 
.A(n_951),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_989),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_990),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_957),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1005),
.A2(n_859),
.B1(n_872),
.B2(n_838),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1000),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_981),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1007),
.B(n_884),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_978),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_SL g1062 ( 
.A(n_1046),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1021),
.B(n_874),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1023),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1024),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1025),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1010),
.A2(n_986),
.B1(n_971),
.B2(n_941),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_1040),
.A2(n_940),
.B(n_939),
.Y(n_1068)
);

OAI222xp33_ASAP7_75t_L g1069 ( 
.A1(n_1018),
.A2(n_883),
.B1(n_899),
.B2(n_910),
.C1(n_807),
.C2(n_991),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1014),
.A2(n_986),
.B1(n_873),
.B2(n_885),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1040),
.A2(n_973),
.B1(n_972),
.B2(n_957),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_1028),
.B(n_860),
.C(n_877),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1027),
.Y(n_1073)
);

BUFx8_ASAP7_75t_SL g1074 ( 
.A(n_1049),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1031),
.A2(n_885),
.B1(n_887),
.B2(n_884),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1015),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1015),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1031),
.A2(n_891),
.B1(n_887),
.B2(n_967),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1035),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1032),
.A2(n_967),
.B1(n_811),
.B2(n_1008),
.Y(n_1080)
);

BUFx8_ASAP7_75t_L g1081 ( 
.A(n_1009),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1028),
.A2(n_1004),
.B1(n_1003),
.B2(n_1006),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1048),
.A2(n_966),
.B1(n_1007),
.B2(n_992),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_1022),
.Y(n_1084)
);

OAI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1055),
.A2(n_828),
.B1(n_910),
.B2(n_951),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1018),
.A2(n_860),
.B(n_820),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1041),
.A2(n_987),
.B1(n_969),
.B2(n_1001),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1019),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_1022),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1051),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_SL g1091 ( 
.A1(n_1053),
.A2(n_797),
.B1(n_902),
.B2(n_995),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1038),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1042),
.A2(n_969),
.B1(n_987),
.B2(n_1002),
.Y(n_1093)
);

OAI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1013),
.A2(n_1056),
.B1(n_1047),
.B2(n_1039),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1026),
.A2(n_902),
.B1(n_797),
.B2(n_864),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1053),
.A2(n_797),
.B1(n_902),
.B2(n_978),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1056),
.A2(n_797),
.B1(n_978),
.B2(n_504),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1042),
.A2(n_1002),
.B1(n_930),
.B2(n_996),
.Y(n_1098)
);

OAI222xp33_ASAP7_75t_L g1099 ( 
.A1(n_1020),
.A2(n_597),
.B1(n_608),
.B2(n_613),
.C1(n_446),
.C2(n_452),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1045),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1039),
.A2(n_1047),
.B1(n_1054),
.B2(n_1037),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1045),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1017),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1043),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1050),
.B(n_1060),
.Y(n_1105)
);

BUFx12f_ASAP7_75t_L g1106 ( 
.A(n_1037),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1057),
.B(n_854),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1077),
.B(n_1088),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1068),
.A2(n_1057),
.B1(n_1016),
.B2(n_1052),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1072),
.A2(n_875),
.B1(n_571),
.B2(n_1058),
.Y(n_1110)
);

OAI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1070),
.A2(n_613),
.B1(n_608),
.B2(n_1059),
.C(n_901),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1078),
.A2(n_1044),
.B1(n_1033),
.B2(n_1036),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1105),
.A2(n_911),
.B1(n_856),
.B2(n_1030),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1077),
.B(n_1030),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1103),
.B(n_1034),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1067),
.A2(n_856),
.B1(n_1034),
.B2(n_798),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1086),
.A2(n_1029),
.B1(n_1022),
.B2(n_1061),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1080),
.A2(n_798),
.B1(n_1011),
.B2(n_1061),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_L g1119 ( 
.A(n_1099),
.B(n_1012),
.C(n_998),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1088),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1063),
.A2(n_1011),
.B1(n_1061),
.B2(n_1012),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1104),
.B(n_949),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1075),
.A2(n_798),
.B1(n_557),
.B2(n_562),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1091),
.A2(n_798),
.B1(n_557),
.B2(n_562),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1091),
.A2(n_1101),
.B1(n_1107),
.B2(n_1096),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1071),
.A2(n_557),
.B1(n_562),
.B2(n_558),
.Y(n_1126)
);

OAI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1096),
.A2(n_901),
.B1(n_585),
.B2(n_536),
.C(n_587),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1082),
.A2(n_558),
.B1(n_568),
.B2(n_566),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1085),
.A2(n_558),
.B1(n_568),
.B2(n_566),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1085),
.A2(n_568),
.B1(n_569),
.B2(n_566),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1073),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1083),
.A2(n_574),
.B1(n_576),
.B2(n_569),
.Y(n_1132)
);

OAI221xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1095),
.A2(n_560),
.B1(n_536),
.B2(n_585),
.C(n_587),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1094),
.A2(n_959),
.B1(n_961),
.B2(n_949),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1083),
.A2(n_569),
.B1(n_576),
.B2(n_574),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1064),
.B(n_949),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1094),
.A2(n_574),
.B1(n_590),
.B2(n_576),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_SL g1138 ( 
.A1(n_1098),
.A2(n_961),
.B1(n_964),
.B2(n_959),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1065),
.B(n_1066),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1062),
.A2(n_1087),
.B1(n_1081),
.B2(n_1093),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1079),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1092),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1106),
.A2(n_590),
.B1(n_599),
.B2(n_596),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1097),
.A2(n_596),
.B1(n_603),
.B2(n_599),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1076),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1097),
.A2(n_603),
.B1(n_614),
.B2(n_604),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1090),
.A2(n_964),
.B1(n_961),
.B2(n_791),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1069),
.A2(n_580),
.B(n_555),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1100),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1102),
.B(n_548),
.Y(n_1151)
);

OAI21xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1084),
.A2(n_825),
.B(n_844),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1108),
.B(n_1074),
.Y(n_1153)
);

OAI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1109),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1131),
.B(n_49),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1117),
.B(n_509),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1139),
.B(n_50),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_SL g1158 ( 
.A(n_1119),
.B(n_50),
.C(n_51),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1111),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1148),
.A2(n_1141),
.B(n_1131),
.Y(n_1160)
);

AND2x2_ASAP7_75t_SL g1161 ( 
.A(n_1129),
.B(n_509),
.Y(n_1161)
);

AOI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_1125),
.A2(n_509),
.B1(n_511),
.B2(n_516),
.C(n_521),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1114),
.B(n_58),
.Y(n_1163)
);

AND2x2_ASAP7_75t_SL g1164 ( 
.A(n_1130),
.B(n_511),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1114),
.B(n_58),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1140),
.A2(n_59),
.B(n_61),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1141),
.B(n_61),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1110),
.A2(n_818),
.B(n_496),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1112),
.B(n_521),
.C(n_516),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1143),
.B(n_522),
.C(n_496),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1118),
.A2(n_522),
.B1(n_502),
.B2(n_496),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1142),
.B(n_63),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1145),
.B(n_64),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1138),
.B(n_522),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1120),
.A2(n_66),
.B(n_67),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1150),
.B(n_68),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1120),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1123),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1124),
.A2(n_502),
.B1(n_494),
.B2(n_74),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1149),
.B(n_87),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1136),
.B(n_70),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1134),
.B(n_494),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1115),
.B(n_73),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1151),
.A2(n_75),
.B(n_77),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1113),
.B(n_494),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1122),
.B(n_77),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1121),
.B(n_78),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_1126),
.B(n_502),
.C(n_80),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1137),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1116),
.B(n_84),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1128),
.B(n_295),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1132),
.B(n_88),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1177),
.B(n_1149),
.Y(n_1193)
);

OAI211xp5_ASAP7_75t_L g1194 ( 
.A1(n_1166),
.A2(n_1135),
.B(n_1146),
.C(n_1144),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_SL g1195 ( 
.A(n_1158),
.B(n_1127),
.C(n_1133),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1175),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1175),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_L g1198 ( 
.A(n_1154),
.B(n_1152),
.C(n_1147),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1153),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1163),
.B(n_91),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1155),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1155),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1167),
.B(n_97),
.Y(n_1203)
);

NAND4xp75_ASAP7_75t_L g1204 ( 
.A(n_1156),
.B(n_98),
.C(n_99),
.D(n_100),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1159),
.B(n_102),
.C(n_103),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1180),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_1206)
);

XNOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1187),
.B(n_119),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1183),
.B(n_121),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1184),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1157),
.B(n_125),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1184),
.B(n_130),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_L g1212 ( 
.A(n_1188),
.B(n_131),
.C(n_135),
.Y(n_1212)
);

XNOR2x2_ASAP7_75t_L g1213 ( 
.A(n_1211),
.B(n_1174),
.Y(n_1213)
);

XNOR2xp5_ASAP7_75t_L g1214 ( 
.A(n_1207),
.B(n_1165),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1209),
.B(n_1160),
.Y(n_1215)
);

NOR3xp33_ASAP7_75t_L g1216 ( 
.A(n_1205),
.B(n_1190),
.C(n_1162),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1193),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1199),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1201),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1212),
.B(n_1181),
.C(n_1186),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1200),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1202),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1210),
.B(n_1173),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1196),
.B(n_1160),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1197),
.B(n_1172),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1203),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1198),
.B(n_1176),
.Y(n_1227)
);

NAND4xp75_ASAP7_75t_L g1228 ( 
.A(n_1195),
.B(n_1174),
.C(n_1182),
.D(n_1161),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1208),
.B(n_1182),
.Y(n_1229)
);

NOR3xp33_ASAP7_75t_L g1230 ( 
.A(n_1205),
.B(n_1169),
.C(n_1179),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1215),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1218),
.Y(n_1232)
);

XNOR2xp5_ASAP7_75t_L g1233 ( 
.A(n_1214),
.B(n_1206),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1222),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1225),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1227),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1227),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1224),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1221),
.Y(n_1239)
);

XOR2x2_ASAP7_75t_L g1240 ( 
.A(n_1223),
.B(n_1204),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1217),
.B(n_1185),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1219),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1236),
.Y(n_1243)
);

AOI22x1_ASAP7_75t_SL g1244 ( 
.A1(n_1236),
.A2(n_1226),
.B1(n_1213),
.B2(n_1228),
.Y(n_1244)
);

AO22x2_ASAP7_75t_L g1245 ( 
.A1(n_1239),
.A2(n_1220),
.B1(n_1216),
.B2(n_1229),
.Y(n_1245)
);

XNOR2x1_ASAP7_75t_L g1246 ( 
.A(n_1233),
.B(n_1192),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1237),
.A2(n_1221),
.B1(n_1230),
.B2(n_1170),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1240),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1232),
.A2(n_1178),
.B1(n_1189),
.B2(n_1194),
.Y(n_1249)
);

AOI22x1_ASAP7_75t_L g1250 ( 
.A1(n_1239),
.A2(n_1191),
.B1(n_1168),
.B2(n_1164),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1234),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1242),
.Y(n_1252)
);

OA22x2_ASAP7_75t_L g1253 ( 
.A1(n_1235),
.A2(n_1171),
.B1(n_1164),
.B2(n_1161),
.Y(n_1253)
);

XOR2xp5_ASAP7_75t_L g1254 ( 
.A(n_1241),
.B(n_142),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1251),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1243),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1252),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1245),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1247),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1245),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1244),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1248),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1255),
.Y(n_1263)
);

NAND2x1_ASAP7_75t_SL g1264 ( 
.A(n_1261),
.B(n_1238),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1256),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1258),
.A2(n_1253),
.B1(n_1249),
.B2(n_1246),
.Y(n_1266)
);

OAI322xp33_ASAP7_75t_L g1267 ( 
.A1(n_1260),
.A2(n_1231),
.A3(n_1254),
.B1(n_1250),
.B2(n_154),
.C1(n_156),
.C2(n_157),
.Y(n_1267)
);

OAI322xp33_ASAP7_75t_L g1268 ( 
.A1(n_1259),
.A2(n_144),
.A3(n_148),
.B1(n_149),
.B2(n_158),
.C1(n_162),
.C2(n_163),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1265),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1264),
.Y(n_1270)
);

O2A1O1Ixp5_ASAP7_75t_SL g1271 ( 
.A1(n_1263),
.A2(n_1257),
.B(n_1262),
.C(n_169),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1266),
.A2(n_166),
.B1(n_168),
.B2(n_173),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1267),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1268),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1269),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1270),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1272),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1273),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1274),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1271),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1275),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1276),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1281),
.B(n_1277),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1282),
.A2(n_1280),
.B1(n_1279),
.B2(n_1278),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1281),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1285),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_1283),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1284),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1285),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1287),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1287),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_1291)
);

AOI31xp33_ASAP7_75t_L g1292 ( 
.A1(n_1288),
.A2(n_240),
.A3(n_241),
.B(n_244),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1286),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1289),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1291),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1294),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1293),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1295),
.A2(n_1290),
.B1(n_1292),
.B2(n_252),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1297),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1298),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1299),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1300),
.A2(n_1296),
.B1(n_267),
.B2(n_272),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1301),
.A2(n_263),
.B1(n_273),
.B2(n_275),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1302),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1303),
.Y(n_1305)
);

AOI221xp5_ASAP7_75t_L g1306 ( 
.A1(n_1304),
.A2(n_1305),
.B1(n_287),
.B2(n_289),
.C(n_291),
.Y(n_1306)
);

AOI211xp5_ASAP7_75t_L g1307 ( 
.A1(n_1306),
.A2(n_283),
.B(n_293),
.C(n_294),
.Y(n_1307)
);


endmodule