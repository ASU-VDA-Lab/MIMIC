module real_aes_2046_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g571 ( .A(n_0), .B(n_226), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_1), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g149 ( .A(n_2), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_3), .B(n_508), .Y(n_507) );
NAND2xp33_ASAP7_75t_SL g563 ( .A(n_4), .B(n_166), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_5), .B(n_210), .Y(n_218) );
INVx1_ASAP7_75t_L g556 ( .A(n_6), .Y(n_556) );
INVx1_ASAP7_75t_L g157 ( .A(n_7), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
OAI22x1_ASAP7_75t_R g800 ( .A1(n_9), .A2(n_76), .B1(n_801), .B2(n_802), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_9), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_10), .Y(n_183) );
AND2x2_ASAP7_75t_L g505 ( .A(n_11), .B(n_198), .Y(n_505) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g227 ( .A(n_14), .Y(n_227) );
AOI221x1_ASAP7_75t_L g559 ( .A1(n_15), .A2(n_170), .B1(n_510), .B2(n_560), .C(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_16), .B(n_508), .Y(n_543) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g224 ( .A(n_18), .Y(n_224) );
INVx1_ASAP7_75t_SL g239 ( .A(n_19), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_20), .B(n_160), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_21), .A2(n_27), .B1(n_496), .B2(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_21), .Y(n_835) );
AOI33xp33_ASAP7_75t_L g264 ( .A1(n_22), .A2(n_51), .A3(n_144), .B1(n_152), .B2(n_265), .B3(n_266), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_23), .A2(n_510), .B(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_24), .B(n_226), .Y(n_512) );
AOI221xp5_ASAP7_75t_SL g535 ( .A1(n_25), .A2(n_41), .B1(n_508), .B2(n_510), .C(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g175 ( .A(n_26), .Y(n_175) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_27), .B(n_129), .C(n_320), .Y(n_128) );
INVx1_ASAP7_75t_SL g496 ( .A(n_27), .Y(n_496) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_28), .A2(n_89), .B(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g199 ( .A(n_28), .B(n_89), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_29), .B(n_229), .Y(n_547) );
INVxp67_ASAP7_75t_L g558 ( .A(n_30), .Y(n_558) );
AND2x2_ASAP7_75t_L g531 ( .A(n_31), .B(n_197), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_32), .B(n_150), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_33), .A2(n_510), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_34), .B(n_229), .Y(n_537) );
INVx1_ASAP7_75t_L g143 ( .A(n_35), .Y(n_143) );
AND2x2_ASAP7_75t_L g155 ( .A(n_35), .B(n_146), .Y(n_155) );
AND2x2_ASAP7_75t_L g166 ( .A(n_35), .B(n_149), .Y(n_166) );
OR2x6_ASAP7_75t_L g114 ( .A(n_36), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_37), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_38), .B(n_150), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_39), .A2(n_171), .B1(n_206), .B2(n_210), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_40), .B(n_215), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_42), .A2(n_80), .B1(n_141), .B2(n_510), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_43), .B(n_160), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_44), .B(n_226), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_45), .B(n_137), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_46), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_47), .Y(n_209) );
AND2x2_ASAP7_75t_L g574 ( .A(n_48), .B(n_197), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_49), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_50), .B(n_197), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_52), .B(n_160), .Y(n_195) );
INVx1_ASAP7_75t_L g148 ( .A(n_53), .Y(n_148) );
INVx1_ASAP7_75t_L g162 ( .A(n_53), .Y(n_162) );
AND2x2_ASAP7_75t_L g196 ( .A(n_54), .B(n_197), .Y(n_196) );
AOI221xp5_ASAP7_75t_L g140 ( .A1(n_55), .A2(n_72), .B1(n_141), .B2(n_150), .C(n_156), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_56), .B(n_150), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_57), .B(n_508), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_58), .B(n_171), .Y(n_185) );
AOI21xp5_ASAP7_75t_SL g248 ( .A1(n_59), .A2(n_141), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g522 ( .A(n_60), .B(n_197), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_61), .B(n_229), .Y(n_572) );
INVx1_ASAP7_75t_L g221 ( .A(n_62), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_63), .B(n_226), .Y(n_520) );
AND2x2_ASAP7_75t_SL g548 ( .A(n_64), .B(n_198), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_65), .A2(n_510), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g194 ( .A(n_66), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_67), .B(n_229), .Y(n_513) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_68), .B(n_137), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_69), .A2(n_141), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g146 ( .A(n_70), .Y(n_146) );
INVx1_ASAP7_75t_L g164 ( .A(n_70), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_71), .B(n_150), .Y(n_267) );
AND2x2_ASAP7_75t_L g241 ( .A(n_73), .B(n_170), .Y(n_241) );
INVx1_ASAP7_75t_L g222 ( .A(n_74), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_75), .A2(n_141), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_76), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_77), .A2(n_141), .B(n_212), .C(n_216), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_78), .B(n_508), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_79), .A2(n_83), .B1(n_150), .B2(n_508), .Y(n_584) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_82), .B(n_170), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_84), .A2(n_141), .B1(n_262), .B2(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_85), .B(n_226), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_86), .B(n_226), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_87), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_88), .A2(n_510), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g250 ( .A(n_90), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_91), .B(n_229), .Y(n_519) );
AND2x2_ASAP7_75t_L g268 ( .A(n_92), .B(n_170), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_93), .A2(n_173), .B(n_174), .C(n_177), .Y(n_172) );
INVxp67_ASAP7_75t_L g561 ( .A(n_94), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_95), .B(n_508), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_96), .B(n_229), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_97), .A2(n_510), .B(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_SL g108 ( .A(n_98), .Y(n_108) );
BUFx2_ASAP7_75t_L g819 ( .A(n_98), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_99), .B(n_160), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_100), .A2(n_102), .B1(n_120), .B2(n_813), .C(n_821), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g832 ( .A1(n_100), .A2(n_833), .B1(n_834), .B2(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_100), .Y(n_833) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B(n_118), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx8_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g820 ( .A(n_111), .Y(n_820) );
BUFx3_ASAP7_75t_L g826 ( .A(n_111), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_112), .B(n_114), .Y(n_126) );
OR2x6_ASAP7_75t_SL g798 ( .A(n_112), .B(n_113), .Y(n_798) );
OR2x2_ASAP7_75t_L g807 ( .A(n_112), .B(n_114), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx2_ASAP7_75t_L g818 ( .A(n_118), .Y(n_818) );
OR2x2_ASAP7_75t_SL g839 ( .A(n_118), .B(n_819), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_808), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_799), .B(n_803), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B1(n_498), .B2(n_796), .Y(n_122) );
CKINVDCx6p67_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
CKINVDCx11_ASAP7_75t_R g812 ( .A(n_124), .Y(n_812) );
INVx3_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
AOI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_391), .B(n_494), .C(n_497), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_128), .A2(n_391), .B(n_494), .Y(n_810) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_130), .A2(n_392), .B(n_496), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_130), .B(n_469), .Y(n_830) );
NOR2x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_298), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_281), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_200), .B1(n_242), .B2(n_256), .C(n_271), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_187), .Y(n_133) );
NAND2x1_ASAP7_75t_SL g307 ( .A(n_134), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g334 ( .A(n_134), .B(n_304), .Y(n_334) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_134), .Y(n_380) );
AND2x2_ASAP7_75t_L g388 ( .A(n_134), .B(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g492 ( .A(n_134), .Y(n_492) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_136), .Y(n_270) );
INVx1_ASAP7_75t_L g286 ( .A(n_136), .Y(n_286) );
AND2x4_ASAP7_75t_L g293 ( .A(n_136), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_136), .B(n_168), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_136), .B(n_289), .Y(n_330) );
INVx1_ASAP7_75t_L g341 ( .A(n_136), .Y(n_341) );
INVxp67_ASAP7_75t_L g375 ( .A(n_136), .Y(n_375) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B(n_167), .Y(n_136) );
INVx2_ASAP7_75t_SL g216 ( .A(n_137), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_137), .A2(n_543), .B(n_544), .Y(n_542) );
BUFx4f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_139), .B(n_199), .Y(n_198) );
AND2x4_ASAP7_75t_L g210 ( .A(n_139), .B(n_199), .Y(n_210) );
INVxp67_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_141), .A2(n_150), .B1(n_555), .B2(n_557), .Y(n_554) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
NOR2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g266 ( .A(n_144), .Y(n_266) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x6_ASAP7_75t_L g158 ( .A(n_145), .B(n_152), .Y(n_158) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g226 ( .A(n_146), .B(n_161), .Y(n_226) );
AND2x6_ASAP7_75t_L g510 ( .A(n_147), .B(n_155), .Y(n_510) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx2_ASAP7_75t_L g152 ( .A(n_148), .Y(n_152) );
AND2x4_ASAP7_75t_L g229 ( .A(n_148), .B(n_163), .Y(n_229) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_149), .Y(n_153) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
INVx1_ASAP7_75t_L g207 ( .A(n_151), .Y(n_207) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVxp33_ASAP7_75t_L g265 ( .A(n_152), .Y(n_265) );
INVx1_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_158), .B(n_159), .C(n_165), .Y(n_156) );
INVxp67_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_158), .A2(n_165), .B(n_194), .C(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_176), .B1(n_221), .B2(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_158), .A2(n_165), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_158), .A2(n_165), .B(n_250), .C(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
AND2x4_ASAP7_75t_L g508 ( .A(n_160), .B(n_166), .Y(n_508) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_165), .B(n_210), .Y(n_230) );
INVx1_ASAP7_75t_L g262 ( .A(n_165), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_165), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_165), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_165), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_165), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_165), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_165), .A2(n_571), .B(n_572), .Y(n_570) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_166), .Y(n_177) );
INVx2_ASAP7_75t_L g258 ( .A(n_168), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_168), .B(n_189), .Y(n_274) );
INVx1_ASAP7_75t_L g292 ( .A(n_168), .Y(n_292) );
INVx1_ASAP7_75t_L g339 ( .A(n_168), .Y(n_339) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_180), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B1(n_178), .B2(n_179), .Y(n_169) );
INVx3_ASAP7_75t_L g179 ( .A(n_170), .Y(n_179) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_171), .B(n_182), .Y(n_181) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_171), .A2(n_568), .B(n_574), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_176), .B(n_210), .C(n_563), .Y(n_562) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_196), .Y(n_189) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_179), .A2(n_190), .B(n_196), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_187), .B(n_311), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_187), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g347 ( .A(n_187), .B(n_293), .Y(n_347) );
INVx1_ASAP7_75t_L g356 ( .A(n_187), .Y(n_356) );
AND2x2_ASAP7_75t_L g404 ( .A(n_187), .B(n_303), .Y(n_404) );
OR2x2_ASAP7_75t_L g447 ( .A(n_187), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x4_ASAP7_75t_L g287 ( .A(n_188), .B(n_288), .Y(n_287) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_188), .B(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g269 ( .A(n_189), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_189), .B(n_289), .Y(n_367) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_189), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_197), .Y(n_234) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_197), .A2(n_535), .B(n_539), .Y(n_534) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_231), .Y(n_201) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_202), .B(n_326), .Y(n_371) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g333 ( .A(n_203), .B(n_324), .Y(n_333) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
INVx1_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
AND2x4_ASAP7_75t_L g279 ( .A(n_204), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g283 ( .A(n_204), .Y(n_283) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_204), .Y(n_319) );
AND2x2_ASAP7_75t_L g489 ( .A(n_204), .B(n_245), .Y(n_489) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_211), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .C(n_209), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_210), .A2(n_248), .B(n_252), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_210), .A2(n_507), .B(n_509), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_210), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_210), .B(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_210), .B(n_561), .Y(n_560) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_216), .A2(n_260), .B(n_268), .Y(n_259) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_216), .A2(n_260), .B(n_268), .Y(n_289) );
AOI21x1_ASAP7_75t_L g582 ( .A1(n_216), .A2(n_583), .B(n_586), .Y(n_582) );
INVx3_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
INVx2_ASAP7_75t_L g297 ( .A(n_217), .Y(n_297) );
NOR2x1_ASAP7_75t_SL g314 ( .A(n_217), .B(n_245), .Y(n_314) );
AND2x2_ASAP7_75t_L g352 ( .A(n_217), .B(n_233), .Y(n_352) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_223), .B(n_230), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B1(n_227), .B2(n_228), .Y(n_223) );
INVxp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g426 ( .A(n_231), .Y(n_426) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g255 ( .A(n_232), .Y(n_255) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
INVx1_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
INVx1_ASAP7_75t_L g384 ( .A(n_233), .Y(n_384) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_233), .Y(n_403) );
OR2x2_ASAP7_75t_L g409 ( .A(n_233), .B(n_245), .Y(n_409) );
AND2x2_ASAP7_75t_L g453 ( .A(n_233), .B(n_280), .Y(n_453) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_234), .A2(n_516), .B(n_522), .Y(n_515) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_234), .A2(n_525), .B(n_531), .Y(n_524) );
AO21x2_ASAP7_75t_L g663 ( .A1(n_234), .A2(n_525), .B(n_531), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_254), .Y(n_243) );
AND2x2_ASAP7_75t_L g295 ( .A(n_244), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g449 ( .A(n_244), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g454 ( .A(n_244), .Y(n_454) );
AND2x2_ASAP7_75t_L g466 ( .A(n_244), .B(n_352), .Y(n_466) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_253), .Y(n_244) );
INVx4_ASAP7_75t_L g277 ( .A(n_245), .Y(n_277) );
INVx2_ASAP7_75t_L g327 ( .A(n_245), .Y(n_327) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_245), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_245), .B(n_385), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_245), .B(n_255), .Y(n_458) );
AND2x2_ASAP7_75t_L g484 ( .A(n_245), .B(n_297), .Y(n_484) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x4_ASAP7_75t_L g386 ( .A(n_253), .B(n_277), .Y(n_386) );
AND2x2_ASAP7_75t_L g313 ( .A(n_254), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_254), .B(n_318), .Y(n_331) );
INVx1_ASAP7_75t_L g365 ( .A(n_254), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_254), .B(n_279), .Y(n_421) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_255), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_256), .A2(n_338), .B1(n_482), .B2(n_485), .Y(n_481) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_269), .Y(n_256) );
INVx1_ASAP7_75t_L g411 ( .A(n_257), .Y(n_411) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g285 ( .A(n_258), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g434 ( .A(n_258), .B(n_306), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_258), .B(n_306), .Y(n_443) );
INVx2_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
AND2x4_ASAP7_75t_L g304 ( .A(n_259), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_261), .B(n_267), .Y(n_260) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_270), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_273), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_273), .B(n_293), .Y(n_378) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g416 ( .A(n_274), .B(n_330), .Y(n_416) );
INVxp33_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_L g397 ( .A(n_276), .Y(n_397) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x4_ASAP7_75t_SL g318 ( .A(n_277), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_277), .Y(n_343) );
INVx2_ASAP7_75t_L g407 ( .A(n_278), .Y(n_407) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_278), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g348 ( .A(n_279), .B(n_327), .Y(n_348) );
AND2x2_ASAP7_75t_L g282 ( .A(n_280), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g385 ( .A(n_280), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B1(n_290), .B2(n_295), .Y(n_281) );
AND2x2_ASAP7_75t_L g310 ( .A(n_282), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g415 ( .A(n_282), .Y(n_415) );
INVx1_ASAP7_75t_L g364 ( .A(n_283), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g322 ( .A1(n_284), .A2(n_323), .B1(n_328), .B2(n_331), .Y(n_322) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_L g448 ( .A(n_285), .Y(n_448) );
BUFx3_ASAP7_75t_L g413 ( .A(n_286), .Y(n_413) );
INVx1_ASAP7_75t_L g436 ( .A(n_287), .Y(n_436) );
AND2x2_ASAP7_75t_L g374 ( .A(n_288), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g441 ( .A(n_288), .B(n_306), .Y(n_441) );
INVx1_ASAP7_75t_L g475 ( .A(n_288), .Y(n_475) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI21xp33_ASAP7_75t_L g312 ( .A1(n_290), .A2(n_313), .B(n_315), .Y(n_312) );
OA21x2_ASAP7_75t_L g346 ( .A1(n_290), .A2(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g423 ( .A(n_292), .Y(n_423) );
AND2x2_ASAP7_75t_L g440 ( .A(n_292), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g430 ( .A(n_293), .B(n_389), .Y(n_430) );
AND2x2_ASAP7_75t_L g433 ( .A(n_293), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g442 ( .A(n_293), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g387 ( .A(n_296), .B(n_386), .Y(n_387) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2x1_ASAP7_75t_L g325 ( .A(n_297), .B(n_326), .Y(n_325) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_297), .B(n_402), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_309), .B(n_312), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_307), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_302), .A2(n_318), .B1(n_343), .B2(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_306), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_308), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_308), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g450 ( .A(n_311), .Y(n_450) );
AND2x2_ASAP7_75t_L g437 ( .A(n_314), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_R g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_318), .B(n_401), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_320), .Y(n_495) );
OR3x2_ASAP7_75t_L g829 ( .A(n_320), .B(n_393), .C(n_830), .Y(n_829) );
NAND3x1_ASAP7_75t_SL g320 ( .A(n_321), .B(n_335), .C(n_349), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_332), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_323), .A2(n_433), .B1(n_435), .B2(n_437), .Y(n_432) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_324), .B(n_363), .Y(n_377) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_329), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g398 ( .A(n_329), .B(n_339), .Y(n_398) );
AND2x2_ASAP7_75t_L g422 ( .A(n_329), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_333), .A2(n_429), .B(n_430), .Y(n_428) );
AND2x2_ASAP7_75t_L g480 ( .A(n_333), .B(n_359), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_334), .A2(n_487), .B1(n_490), .B2(n_493), .Y(n_486) );
AOI21xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_342), .B(n_346), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
BUFx2_ASAP7_75t_L g456 ( .A(n_339), .Y(n_456) );
INVx1_ASAP7_75t_SL g463 ( .A(n_339), .Y(n_463) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_340), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_350), .B(n_369), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g358 ( .A(n_352), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_352), .B(n_363), .Y(n_444) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_360), .B(n_366), .Y(n_357) );
OR2x6_ASAP7_75t_L g414 ( .A(n_359), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g464 ( .A(n_367), .Y(n_464) );
OR2x2_ASAP7_75t_L g491 ( .A(n_367), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_368), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_379), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_376), .B2(n_378), .Y(n_370) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_373), .Y(n_471) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_387), .B2(n_388), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_467), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_417), .C(n_445), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_405), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_399), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp33_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_410), .B1(n_414), .B2(n_416), .Y(n_405) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_407), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_409), .B(n_415), .Y(n_485) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx3_ASAP7_75t_L g473 ( .A(n_413), .Y(n_473) );
INVx2_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_431), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_428), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B1(n_424), .B2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_427), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_432), .B(n_439), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_434), .B(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g459 ( .A(n_442), .Y(n_459) );
AOI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B(n_451), .C(n_460), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g478 ( .A1(n_448), .A2(n_479), .B(n_481), .C(n_486), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B1(n_457), .B2(n_459), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVxp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_SL g494 ( .A1(n_467), .A2(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_470), .B(n_478), .Y(n_469) );
AOI21xp33_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_472), .B(n_476), .Y(n_470) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp33_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_497), .B(n_812), .Y(n_811) );
AO22x2_ASAP7_75t_L g809 ( .A1(n_498), .A2(n_797), .B1(n_810), .B2(n_811), .Y(n_809) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_707), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_629), .C(n_679), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_596), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_532), .B1(n_549), .B2(n_579), .C(n_588), .Y(n_502) );
INVx1_ASAP7_75t_SL g678 ( .A(n_503), .Y(n_678) );
AND2x4_ASAP7_75t_SL g503 ( .A(n_504), .B(n_514), .Y(n_503) );
INVx2_ASAP7_75t_L g600 ( .A(n_504), .Y(n_600) );
OR2x2_ASAP7_75t_L g622 ( .A(n_504), .B(n_613), .Y(n_622) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_504), .Y(n_637) );
INVx5_ASAP7_75t_L g644 ( .A(n_504), .Y(n_644) );
AND2x4_ASAP7_75t_L g650 ( .A(n_504), .B(n_524), .Y(n_650) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_504), .B(n_581), .Y(n_653) );
OR2x2_ASAP7_75t_L g662 ( .A(n_504), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g669 ( .A(n_504), .B(n_515), .Y(n_669) );
AND2x2_ASAP7_75t_L g770 ( .A(n_504), .B(n_523), .Y(n_770) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx3_ASAP7_75t_SL g621 ( .A(n_514), .Y(n_621) );
AND2x2_ASAP7_75t_L g665 ( .A(n_514), .B(n_581), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_514), .A2(n_669), .B(n_670), .Y(n_668) );
AND2x2_ASAP7_75t_L g706 ( .A(n_514), .B(n_644), .Y(n_706) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_515), .B(n_524), .Y(n_587) );
OR2x2_ASAP7_75t_L g591 ( .A(n_515), .B(n_524), .Y(n_591) );
INVx1_ASAP7_75t_L g599 ( .A(n_515), .Y(n_599) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_515), .Y(n_611) );
INVx2_ASAP7_75t_L g619 ( .A(n_515), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_515), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g728 ( .A(n_515), .B(n_613), .Y(n_728) );
AND2x2_ASAP7_75t_L g743 ( .A(n_515), .B(n_581), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g612 ( .A(n_524), .B(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_524), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_532), .B(n_736), .Y(n_735) );
NOR2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_540), .Y(n_532) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g565 ( .A(n_534), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_534), .B(n_541), .Y(n_594) );
INVx1_ASAP7_75t_L g604 ( .A(n_534), .Y(n_604) );
INVx2_ASAP7_75t_L g627 ( .A(n_534), .Y(n_627) );
INVx2_ASAP7_75t_L g633 ( .A(n_534), .Y(n_633) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_534), .Y(n_703) );
OR2x2_ASAP7_75t_L g734 ( .A(n_534), .B(n_541), .Y(n_734) );
OR2x2_ASAP7_75t_L g750 ( .A(n_540), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_541), .B(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g577 ( .A(n_541), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g614 ( .A(n_541), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g639 ( .A(n_541), .B(n_605), .Y(n_639) );
OR2x2_ASAP7_75t_L g647 ( .A(n_541), .B(n_553), .Y(n_647) );
INVx2_ASAP7_75t_L g674 ( .A(n_541), .Y(n_674) );
INVx1_ASAP7_75t_L g692 ( .A(n_541), .Y(n_692) );
NOR2xp33_ASAP7_75t_R g725 ( .A(n_541), .B(n_566), .Y(n_725) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_575), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_550), .A2(n_617), .B1(n_620), .B2(n_623), .Y(n_616) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_564), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g631 ( .A(n_552), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g666 ( .A(n_552), .B(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g745 ( .A(n_552), .B(n_723), .Y(n_745) );
INVx3_ASAP7_75t_L g578 ( .A(n_553), .Y(n_578) );
AND2x4_ASAP7_75t_L g605 ( .A(n_553), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_553), .B(n_566), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_553), .B(n_627), .Y(n_672) );
AND2x2_ASAP7_75t_L g677 ( .A(n_553), .B(n_674), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_553), .B(n_565), .Y(n_714) );
INVx1_ASAP7_75t_L g784 ( .A(n_553), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_553), .B(n_702), .Y(n_795) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g576 ( .A(n_566), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_566), .B(n_578), .Y(n_595) );
INVx2_ASAP7_75t_L g606 ( .A(n_566), .Y(n_606) );
AND2x2_ASAP7_75t_L g632 ( .A(n_566), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_627), .Y(n_648) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_566), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_566), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g737 ( .A(n_566), .Y(n_737) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_576), .B(n_604), .Y(n_615) );
AOI221x1_ASAP7_75t_SL g709 ( .A1(n_577), .A2(n_710), .B1(n_713), .B2(n_715), .C(n_719), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_577), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g767 ( .A(n_577), .B(n_632), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_577), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g698 ( .A(n_578), .B(n_626), .Y(n_698) );
AND2x2_ASAP7_75t_L g736 ( .A(n_578), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_587), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_581), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g684 ( .A(n_581), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_581), .B(n_600), .Y(n_689) );
AND2x4_ASAP7_75t_L g718 ( .A(n_581), .B(n_619), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_581), .B(n_650), .Y(n_754) );
OR2x2_ASAP7_75t_L g772 ( .A(n_581), .B(n_703), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_581), .B(n_663), .Y(n_782) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g613 ( .A(n_582), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_587), .A2(n_646), .B1(n_649), .B2(n_651), .Y(n_645) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
INVx2_ASAP7_75t_L g601 ( .A(n_589), .Y(n_601) );
AND2x2_ASAP7_75t_L g740 ( .A(n_590), .B(n_600), .Y(n_740) );
AND2x2_ASAP7_75t_L g786 ( .A(n_590), .B(n_653), .Y(n_786) );
AND2x2_ASAP7_75t_L g791 ( .A(n_590), .B(n_642), .Y(n_791) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI32xp33_ASAP7_75t_L g760 ( .A1(n_592), .A2(n_662), .A3(n_742), .B1(n_761), .B2(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g628 ( .A(n_595), .Y(n_628) );
AOI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_602), .B(n_607), .C(n_616), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_599), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_600), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g780 ( .A(n_600), .Y(n_780) );
AND2x2_ASAP7_75t_L g690 ( .A(n_602), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_603), .B(n_605), .Y(n_602) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_603), .Y(n_790) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_604), .Y(n_659) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_604), .Y(n_759) );
INVx1_ASAP7_75t_L g656 ( .A(n_605), .Y(n_656) );
AND2x2_ASAP7_75t_L g722 ( .A(n_605), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_605), .B(n_733), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_614), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_609), .A2(n_689), .B(n_690), .Y(n_688) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g618 ( .A(n_613), .B(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g642 ( .A(n_613), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_618), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g749 ( .A(n_618), .Y(n_749) );
AND2x2_ASAP7_75t_L g779 ( .A(n_618), .B(n_780), .Y(n_779) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_619), .Y(n_756) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_621), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g696 ( .A(n_622), .Y(n_696) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g655 ( .A(n_626), .B(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_627), .Y(n_723) );
AND2x2_ASAP7_75t_L g732 ( .A(n_628), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_652), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_639), .B2(n_640), .C(n_645), .Y(n_630) );
INVx1_ASAP7_75t_L g751 ( .A(n_632), .Y(n_751) );
INVxp33_ASAP7_75t_SL g783 ( .A(n_632), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_634), .A2(n_730), .B(n_738), .Y(n_729) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_638), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g651 ( .A(n_639), .Y(n_651) );
AND2x2_ASAP7_75t_L g686 ( .A(n_639), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_639), .B(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_639), .A2(n_767), .B1(n_768), .B2(n_771), .Y(n_766) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g661 ( .A(n_642), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_642), .B(n_650), .Y(n_700) );
AND2x4_ASAP7_75t_L g717 ( .A(n_644), .B(n_663), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_644), .B(n_718), .Y(n_764) );
AND2x2_ASAP7_75t_L g776 ( .A(n_644), .B(n_728), .Y(n_776) );
NAND2xp33_ASAP7_75t_L g761 ( .A(n_646), .B(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_SL g704 ( .A(n_647), .Y(n_704) );
INVx1_ASAP7_75t_L g775 ( .A(n_648), .Y(n_775) );
INVx2_ASAP7_75t_SL g727 ( .A(n_650), .Y(n_727) );
AOI211xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_657), .C(n_675), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_664), .C(n_668), .Y(n_657) );
OR2x6_ASAP7_75t_SL g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g687 ( .A(n_659), .Y(n_687) );
INVx1_ASAP7_75t_SL g712 ( .A(n_662), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_662), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_667), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g753 ( .A1(n_671), .A2(n_754), .B1(n_755), .B2(n_757), .Y(n_753) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_685), .B(n_688), .C(n_693), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_705), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g785 ( .A1(n_704), .A2(n_786), .B1(n_787), .B2(n_791), .C1(n_792), .C2(n_794), .Y(n_785) );
INVx2_ASAP7_75t_L g720 ( .A(n_706), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_746), .C(n_765), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_729), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_717), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_718), .B(n_780), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_724), .B2(n_726), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVxp33_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_727), .B(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_735), .A2(n_739), .B1(n_741), .B2(n_744), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
OAI211xp5_ASAP7_75t_SL g746 ( .A1(n_747), .A2(n_750), .B(n_752), .C(n_760), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_773), .C(n_785), .Y(n_765) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_777), .B(n_784), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_781), .B(n_783), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
INVxp33_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_800), .B(n_809), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx1_ASAP7_75t_SL g838 ( .A(n_820), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_837), .B(n_839), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_827), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
AOI22x1_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B1(n_831), .B2(n_832), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g836 ( .A(n_834), .Y(n_836) );
endmodule