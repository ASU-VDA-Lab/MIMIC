module fake_aes_103_n_17 (n_1, n_2, n_4, n_3, n_5, n_0, n_17);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g6 ( .A(n_0), .Y(n_6) );
O2A1O1Ixp5_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_1), .B(n_0), .C(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
AO21x2_ASAP7_75t_L g10 ( .A1(n_6), .A2(n_3), .B(n_4), .Y(n_10) );
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_4), .B1(n_5), .B2(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
NAND4xp25_ASAP7_75t_L g14 ( .A(n_12), .B(n_7), .C(n_10), .D(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
XNOR2x1_ASAP7_75t_L g16 ( .A(n_15), .B(n_9), .Y(n_16) );
OAI21xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_14), .B(n_7), .Y(n_17) );
endmodule