module fake_jpeg_17705_n_171 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_45),
.B1(n_64),
.B2(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_45),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_58),
.B1(n_57),
.B2(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_98),
.B1(n_104),
.B2(n_115),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_62),
.B1(n_60),
.B2(n_56),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_49),
.B1(n_59),
.B2(n_61),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_117),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_80),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_63),
.B1(n_52),
.B2(n_47),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_1),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_110),
.B1(n_116),
.B2(n_93),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_113),
.B1(n_95),
.B2(n_4),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_2),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_105),
.B1(n_102),
.B2(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_139),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_97),
.B1(n_100),
.B2(n_46),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_5),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_3),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_120),
.B1(n_125),
.B2(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_142),
.B1(n_135),
.B2(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_124),
.B1(n_126),
.B2(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_121),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_119),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_132),
.B(n_137),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_5),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_143),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_150),
.B(n_153),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_22),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_6),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_156),
.C(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_8),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_151),
.B(n_28),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_27),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_25),
.B(n_42),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_21),
.B(n_40),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_20),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_29),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_18),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_30),
.C(n_39),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_16),
.C(n_38),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_15),
.C(n_36),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_14),
.Y(n_171)
);


endmodule