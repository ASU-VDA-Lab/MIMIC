module real_jpeg_1159_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_39),
.B1(n_61),
.B2(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_1),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_3),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_34),
.B1(n_37),
.B2(n_100),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_100),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_100),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_34),
.B1(n_37),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_34),
.B1(n_37),
.B2(n_54),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_6),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_321)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_8),
.B(n_28),
.C(n_30),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_27),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_8),
.B(n_47),
.C(n_50),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_197),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_8),
.B(n_93),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_8),
.B(n_79),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_8),
.A2(n_34),
.B1(n_37),
.B2(n_197),
.Y(n_262)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_122),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_11),
.A2(n_34),
.B1(n_37),
.B2(n_122),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_122),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_12),
.A2(n_34),
.B1(n_37),
.B2(n_56),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_12),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_13),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_42),
.B1(n_61),
.B2(n_62),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_15),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_34),
.B1(n_37),
.B2(n_161),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_161),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_327),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_314),
.B(n_326),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_137),
.B(n_311),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_125),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_101),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_22),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_22),
.B(n_101),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_22),
.B(n_126),
.Y(n_313)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.CI(n_82),
.CON(n_22),
.SN(n_22)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_24),
.B(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_25),
.A2(n_40),
.B1(n_41),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_25),
.A2(n_38),
.B1(n_40),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_25),
.A2(n_40),
.B1(n_76),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_25),
.A2(n_40),
.B1(n_170),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_25),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_25),
.A2(n_201),
.B(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_26),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_26),
.A2(n_27),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_27),
.B(n_158),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_30),
.B(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_34),
.A2(n_37),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_34),
.B(n_187),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_34),
.B(n_69),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_37),
.A2(n_62),
.A3(n_68),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_40),
.A2(n_118),
.B(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_40),
.A2(n_157),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_53),
.B2(n_55),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_49),
.B1(n_53),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_44),
.A2(n_182),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_44),
.A2(n_49),
.B1(n_180),
.B2(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_45),
.A2(n_79),
.B1(n_87),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_45),
.A2(n_79),
.B1(n_116),
.B2(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_45),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_45),
.B(n_183),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_49),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_49),
.A2(n_204),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_50),
.B(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_73),
.B2(n_81),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_59),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g136 ( 
.A(n_59),
.B(n_74),
.C(n_78),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_59),
.B(n_129),
.C(n_136),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_67),
.B2(n_72),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_67),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_62),
.A2(n_65),
.B(n_197),
.C(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_62),
.B(n_197),
.Y(n_198)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_67),
.B1(n_72),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_66),
.A2(n_121),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_66),
.A2(n_162),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_66),
.A2(n_162),
.B1(n_321),
.B2(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_67),
.A2(n_97),
.B(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_78),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_78),
.B(n_130),
.C(n_134),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_79),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B(n_96),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_85),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_89),
.B1(n_96),
.B2(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_93),
.B1(n_113),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_90),
.A2(n_197),
.B(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_91),
.A2(n_92),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_91),
.A2(n_92),
.B1(n_177),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_91),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_91),
.A2(n_92),
.B1(n_222),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_92),
.A2(n_176),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_92),
.B(n_191),
.Y(n_224)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_93),
.A2(n_190),
.B(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_117),
.C(n_119),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_110),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_111),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_119),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_124),
.B(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_125),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_131),
.Y(n_320)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_135),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_163),
.B(n_310),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_139),
.B(n_142),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_148),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_143),
.B(n_146),
.Y(n_308)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_148),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.C(n_159),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_149),
.A2(n_150),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_151),
.B(n_153),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_305),
.B(n_309),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_274),
.B(n_302),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_216),
.B(n_273),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_192),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_192),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.C(n_184),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_168),
.B(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_172),
.C(n_175),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_178),
.B(n_184),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_206),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_193),
.B(n_207),
.C(n_215),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_205),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_194),
.B(n_200),
.C(n_202),
.Y(n_287)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_213),
.Y(n_278)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_268),
.B(n_272),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_257),
.B(n_267),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_239),
.B(n_256),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_225),
.B1(n_231),
.B2(n_232),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_228),
.C(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_250),
.B(n_255),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_248),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.C(n_265),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_289),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_288),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_288),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_286),
.C(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.C(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_301),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_295),
.C(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);


endmodule