module real_jpeg_1736_n_17 (n_108, n_8, n_0, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_100, n_106, n_11, n_14, n_110, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_101, n_1, n_16, n_15, n_13, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_100;
input n_106;
input n_11;
input n_14;
input n_110;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_101;
input n_1;
input n_16;
input n_15;
input n_13;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.C(n_62),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_4),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_44),
.B(n_48),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_39),
.C(n_54),
.Y(n_38)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_35),
.B1(n_68),
.B2(n_71),
.Y(n_34)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_26),
.B1(n_97),
.B2(n_98),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_19),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_23),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_24),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI221xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_73),
.C(n_87),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_30),
.B(n_86),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_64),
.C(n_65),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_57),
.C(n_58),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.C(n_52),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_82),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_88),
.A3(n_89),
.B1(n_92),
.B2(n_93),
.C1(n_96),
.C2(n_110),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.C(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_100),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_101),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_102),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_103),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_104),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_105),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_106),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_107),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_108),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_109),
.Y(n_86)
);


endmodule