module fake_netlist_1_6421_n_721 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_721);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_721;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_26), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_63), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_20), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_22), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_24), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_32), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
NOR2xp67_ASAP7_75t_L g89 ( .A(n_61), .B(n_25), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_39), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_78), .Y(n_91) );
NOR2xp67_ASAP7_75t_L g92 ( .A(n_70), .B(n_45), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_57), .Y(n_93) );
BUFx10_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_6), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_41), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_55), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_67), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_40), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_5), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_1), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_1), .Y(n_102) );
BUFx8_ASAP7_75t_SL g103 ( .A(n_64), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_65), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_76), .B(n_51), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_46), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_54), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_60), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_49), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_28), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_29), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_44), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_79), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_43), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_8), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_34), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_87), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_118), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_119), .B(n_0), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_119), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_124), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_80), .B(n_0), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_108), .B(n_27), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_122), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_122), .Y(n_144) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_81), .A2(n_30), .B(n_74), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_83), .A2(n_23), .B(n_73), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_100), .B(n_2), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_84), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_101), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_103), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_105), .Y(n_153) );
OAI22x1_ASAP7_75t_R g154 ( .A1(n_95), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_104), .B(n_7), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_109), .B(n_9), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_94), .B(n_9), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_114), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_112), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_123), .B(n_10), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_101), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_101), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_98), .B(n_47), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_127), .B(n_11), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_85), .B(n_14), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_94), .B(n_15), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_168), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_130), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_168), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_133), .B(n_127), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_168), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_86), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g181 ( .A(n_157), .B(n_127), .C(n_86), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_158), .B(n_94), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_129), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_129), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_162), .B(n_117), .Y(n_188) );
BUFx8_ASAP7_75t_SL g189 ( .A(n_133), .Y(n_189) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_157), .B(n_85), .C(n_121), .Y(n_190) );
INVxp67_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_146), .B(n_170), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_146), .B(n_110), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_130), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_158), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
INVxp67_ASAP7_75t_SL g201 ( .A(n_172), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_151), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_170), .B(n_91), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g204 ( .A1(n_149), .A2(n_95), .B1(n_120), .B2(n_93), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_170), .B(n_107), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_140), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_152), .B(n_111), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_125), .B1(n_120), .B2(n_93), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_152), .B(n_116), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_160), .B(n_97), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_172), .B(n_113), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_160), .B(n_96), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_137), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_143), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_135), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_141), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_144), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_131), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_141), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_151), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_148), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_144), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_161), .B(n_125), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_161), .B(n_106), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_131), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_182), .B(n_164), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_201), .B(n_164), .Y(n_239) );
OAI221xp5_ASAP7_75t_L g240 ( .A1(n_235), .A2(n_171), .B1(n_156), .B2(n_139), .C(n_153), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_186), .B(n_141), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_230), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_211), .A2(n_99), .B1(n_159), .B2(n_153), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_225), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_188), .A2(n_141), .B1(n_167), .B2(n_134), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_183), .B(n_132), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
O2A1O1Ixp5_ASAP7_75t_L g248 ( .A1(n_185), .A2(n_130), .B(n_132), .C(n_142), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_227), .Y(n_250) );
BUFx6f_ASAP7_75t_SL g251 ( .A(n_188), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_183), .B(n_132), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_230), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_237), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_237), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_185), .B(n_144), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_99), .B1(n_138), .B2(n_142), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_231), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_231), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_185), .B(n_89), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_214), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_179), .B(n_136), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_185), .B(n_92), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_207), .Y(n_264) );
NOR3xp33_ASAP7_75t_L g265 ( .A(n_204), .B(n_136), .C(n_138), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_191), .B(n_136), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_217), .B(n_167), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_200), .B(n_145), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_216), .B(n_167), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_214), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_188), .A2(n_167), .B1(n_147), .B2(n_145), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_209), .B(n_167), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_216), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_186), .B(n_167), .Y(n_274) );
AND2x6_ASAP7_75t_SL g275 ( .A(n_189), .B(n_154), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_194), .B(n_167), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_207), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_200), .B(n_226), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_203), .B(n_147), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_198), .B(n_147), .Y(n_281) );
NOR2x2_ASAP7_75t_L g282 ( .A(n_198), .B(n_154), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_147), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_232), .B(n_169), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_192), .B(n_169), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_214), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_202), .B(n_15), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_218), .B(n_165), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_219), .Y(n_289) );
BUFx5_ASAP7_75t_L g290 ( .A(n_182), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_200), .B(n_166), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_218), .B(n_165), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_188), .A2(n_166), .B1(n_163), .B2(n_150), .Y(n_294) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_231), .B(n_163), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_193), .A2(n_166), .B1(n_163), .B2(n_150), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_233), .B(n_166), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_233), .B(n_166), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_233), .B(n_163), .Y(n_299) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_181), .A2(n_163), .B(n_150), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_193), .B(n_150), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_199), .B(n_150), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_199), .B(n_16), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_222), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_205), .B(n_17), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_205), .B(n_18), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_240), .A2(n_205), .B1(n_180), .B2(n_176), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_239), .B(n_188), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_241), .A2(n_226), .B(n_200), .Y(n_310) );
AO22x1_ASAP7_75t_L g311 ( .A1(n_257), .A2(n_202), .B1(n_188), .B2(n_226), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_246), .B(n_188), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_253), .A2(n_181), .B(n_173), .C(n_180), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_252), .B(n_190), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_266), .B(n_190), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_304), .A2(n_173), .B1(n_176), .B2(n_178), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_273), .B(n_177), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_254), .B(n_177), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_284), .B(n_213), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_257), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_281), .A2(n_212), .B1(n_178), .B2(n_226), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_280), .A2(n_182), .B(n_224), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_243), .A2(n_236), .B1(n_231), .B2(n_224), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_268), .A2(n_222), .B(n_196), .C(n_174), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_265), .B(n_231), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_238), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_241), .A2(n_174), .B(n_196), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_258), .B(n_210), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_269), .B(n_234), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_258), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_244), .B(n_234), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_258), .B(n_229), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_283), .B(n_229), .C(n_228), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_255), .B(n_228), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_262), .B(n_223), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_242), .A2(n_223), .B(n_221), .C(n_220), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_274), .A2(n_221), .B(n_220), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_274), .A2(n_272), .B(n_276), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_247), .B(n_215), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_278), .A2(n_215), .B(n_210), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g343 ( .A1(n_245), .A2(n_208), .B(n_197), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_249), .B(n_208), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_271), .A2(n_197), .B(n_195), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_303), .A2(n_195), .B(n_187), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_238), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_250), .Y(n_348) );
AO22x1_ASAP7_75t_L g349 ( .A1(n_282), .A2(n_187), .B1(n_184), .B2(n_175), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_270), .A2(n_184), .B(n_175), .C(n_31), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_251), .A2(n_19), .B1(n_21), .B2(n_37), .Y(n_351) );
AOI21x1_ASAP7_75t_L g352 ( .A1(n_303), .A2(n_305), .B(n_256), .Y(n_352) );
AND2x6_ASAP7_75t_L g353 ( .A(n_286), .B(n_42), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_264), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_277), .B(n_48), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_279), .B(n_75), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_275), .Y(n_357) );
BUFx8_ASAP7_75t_L g358 ( .A(n_251), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_238), .Y(n_359) );
A2O1A1Ixp33_ASAP7_75t_L g360 ( .A1(n_291), .A2(n_289), .B(n_248), .C(n_300), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_322), .B(n_287), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_267), .B(n_305), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_308), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_352), .A2(n_306), .B(n_300), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_345), .A2(n_302), .B(n_301), .Y(n_365) );
AO31x2_ASAP7_75t_L g366 ( .A1(n_360), .A2(n_296), .A3(n_298), .B(n_297), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g367 ( .A(n_325), .B(n_294), .C(n_260), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_329), .A2(n_292), .B(n_263), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_324), .A2(n_335), .B(n_345), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_320), .B(n_238), .Y(n_370) );
AO31x2_ASAP7_75t_L g371 ( .A1(n_313), .A2(n_296), .A3(n_299), .B(n_293), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_348), .A2(n_288), .B1(n_285), .B2(n_259), .Y(n_372) );
AOI211x1_ASAP7_75t_L g373 ( .A1(n_311), .A2(n_295), .B(n_52), .C(n_53), .Y(n_373) );
AOI21x1_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_356), .B(n_355), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g375 ( .A(n_359), .B(n_50), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_326), .A2(n_290), .B(n_58), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_315), .B(n_290), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_314), .B(n_290), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_290), .B(n_59), .Y(n_379) );
AOI221x1_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_324), .B1(n_343), .B2(n_309), .C(n_312), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_327), .B(n_290), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_319), .B(n_72), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_316), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_318), .B(n_56), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_333), .Y(n_386) );
AO32x2_ASAP7_75t_L g387 ( .A1(n_307), .A2(n_66), .A3(n_317), .B1(n_353), .B2(n_349), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_339), .B(n_334), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_347), .B(n_328), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_332), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_336), .A2(n_342), .B(n_330), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_338), .A2(n_331), .B(n_323), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_321), .A2(n_328), .B1(n_347), .B2(n_358), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_384), .Y(n_395) );
BUFx2_ASAP7_75t_SL g396 ( .A(n_390), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_379), .A2(n_350), .B(n_344), .Y(n_397) );
AOI21x1_ASAP7_75t_L g398 ( .A1(n_374), .A2(n_321), .B(n_353), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_337), .B(n_353), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_369), .A2(n_353), .B(n_332), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_332), .B(n_347), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_392), .B(n_358), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_386), .B(n_357), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_388), .A2(n_376), .B(n_362), .Y(n_404) );
AO31x2_ASAP7_75t_L g405 ( .A1(n_380), .A2(n_378), .A3(n_377), .B(n_372), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_365), .A2(n_391), .B(n_378), .Y(n_407) );
AO21x1_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_381), .B(n_361), .Y(n_408) );
AOI22x1_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_390), .B1(n_385), .B2(n_373), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_367), .B(n_393), .Y(n_410) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_393), .B(n_372), .Y(n_411) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_387), .A2(n_370), .B1(n_389), .B2(n_363), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_382), .A2(n_387), .B(n_366), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_366), .A2(n_387), .B(n_371), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_366), .A2(n_371), .B(n_375), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_363), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_379), .A2(n_374), .B(n_364), .Y(n_421) );
OAI21x1_ASAP7_75t_L g422 ( .A1(n_379), .A2(n_374), .B(n_364), .Y(n_422) );
OAI21x1_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_374), .B(n_364), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_417), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_420), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_406), .B(n_419), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_407), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_415), .B(n_414), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_408), .Y(n_429) );
OAI21x1_ASAP7_75t_L g430 ( .A1(n_421), .A2(n_422), .B(n_423), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_408), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_411), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_411), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_416), .B(n_412), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_418), .B(n_405), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_407), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_418), .B(n_405), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_415), .B(n_399), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_396), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_416), .B(n_412), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_403), .A2(n_402), .B1(n_412), .B2(n_409), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_412), .B(n_396), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_401), .Y(n_446) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_422), .B(n_421), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_405), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_405), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_423), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_409), .A2(n_397), .B(n_404), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_403), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
AND2x6_ASAP7_75t_L g457 ( .A(n_398), .B(n_399), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_403), .B(n_395), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_424), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_426), .B(n_413), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_455), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_429), .B(n_413), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_429), .B(n_413), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_427), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_459), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_431), .B(n_398), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_458), .B(n_397), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_439), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_458), .A2(n_404), .B1(n_444), .B2(n_428), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_431), .B(n_442), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_448), .B(n_451), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_434), .B(n_442), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_428), .B(n_456), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_428), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_428), .B(n_451), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_437), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_448), .B(n_456), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_435), .B(n_438), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_435), .B(n_438), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_440), .B(n_425), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_445), .B(n_446), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_440), .B(n_445), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_432), .A2(n_433), .B1(n_450), .B2(n_443), .C(n_441), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g497 ( .A1(n_454), .A2(n_450), .B(n_443), .C(n_433), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_449), .A2(n_452), .B1(n_446), .B2(n_443), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_443), .B(n_449), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_432), .B(n_452), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_452), .B(n_447), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_457), .Y(n_503) );
AO31x2_ASAP7_75t_L g504 ( .A1(n_453), .A2(n_447), .A3(n_457), .B(n_430), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_447), .B(n_453), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_430), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_457), .B(n_440), .Y(n_509) );
BUFx2_ASAP7_75t_R g510 ( .A(n_457), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_479), .B(n_457), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_500), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_474), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_464), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_500), .B(n_457), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_478), .B(n_457), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_461), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_495), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_479), .B(n_457), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_495), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_488), .B(n_490), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_476), .B(n_488), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_490), .B(n_476), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_482), .B(n_483), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_491), .B(n_462), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_485), .B(n_483), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_485), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_482), .B(n_492), .Y(n_533) );
INVx11_ASAP7_75t_L g534 ( .A(n_510), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_492), .B(n_466), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_463), .B(n_486), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_466), .B(n_473), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_473), .B(n_484), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_473), .B(n_484), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_495), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_477), .B(n_486), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_493), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_474), .B(n_481), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_478), .B(n_503), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_481), .B(n_487), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_487), .B(n_480), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_493), .B(n_489), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_502), .B(n_478), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_467), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_469), .B(n_467), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_509), .B(n_503), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_469), .B(n_468), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_509), .B(n_502), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_471), .B(n_499), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_468), .B(n_465), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_465), .B(n_499), .Y(n_563) );
NOR2x1p5_ASAP7_75t_L g564 ( .A(n_508), .B(n_505), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_499), .B(n_508), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_471), .B(n_506), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_535), .B(n_494), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_527), .B(n_498), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_516), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_526), .B(n_475), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_527), .B(n_505), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_565), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_526), .B(n_506), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_533), .B(n_472), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_564), .B(n_504), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_517), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_554), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_528), .B(n_504), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_565), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_528), .B(n_504), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_564), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_542), .B(n_504), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_513), .B(n_507), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_530), .B(n_504), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_543), .B(n_507), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_533), .B(n_507), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_517), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_513), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_543), .B(n_497), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_515), .B(n_546), .Y(n_591) );
NAND2xp67_ASAP7_75t_SL g592 ( .A(n_511), .B(n_523), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_535), .B(n_553), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_514), .B(n_518), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_551), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_520), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_512), .B(n_531), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_529), .B(n_550), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_513), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_551), .B(n_536), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_561), .B(n_562), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_550), .B(n_553), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_522), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_520), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_521), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_525), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_513), .B(n_541), .C(n_536), .D(n_515), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_532), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_532), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_561), .B(n_562), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_537), .B(n_559), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_563), .B(n_537), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_549), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_559), .B(n_511), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_593), .B(n_523), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_567), .B(n_538), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_567), .B(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_603), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_615), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_578), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_583), .B(n_539), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_578), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_572), .B(n_563), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_595), .B(n_560), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_594), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_593), .B(n_547), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_590), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_591), .B(n_512), .Y(n_636) );
NAND2x1_ASAP7_75t_SL g637 ( .A(n_600), .B(n_558), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_617), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_585), .B(n_539), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_604), .B(n_547), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_574), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_598), .B(n_534), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_591), .B(n_546), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_599), .B(n_545), .Y(n_645) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_600), .B(n_558), .Y(n_646) );
OR2x6_ASAP7_75t_L g647 ( .A(n_589), .B(n_556), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_573), .B(n_549), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_570), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_616), .B(n_545), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_573), .B(n_566), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_601), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_589), .B(n_552), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_546), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_597), .Y(n_657) );
AOI32xp33_ASAP7_75t_L g658 ( .A1(n_628), .A2(n_576), .A3(n_598), .B1(n_619), .B2(n_591), .Y(n_658) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_633), .A2(n_582), .B(n_571), .C(n_579), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_626), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g661 ( .A(n_637), .B(n_576), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_633), .B(n_581), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_647), .A2(n_611), .B1(n_582), .B2(n_556), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_634), .A2(n_576), .B(n_575), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_647), .A2(n_556), .B1(n_584), .B2(n_592), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_623), .B(n_587), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_647), .A2(n_534), .B1(n_584), .B2(n_558), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_648), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_653), .Y(n_669) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_653), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_621), .B(n_580), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_642), .A2(n_558), .B(n_580), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_643), .B(n_541), .Y(n_673) );
NAND2x1_ASAP7_75t_SL g674 ( .A(n_636), .B(n_546), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_656), .B(n_519), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_627), .B(n_639), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_648), .B(n_541), .C(n_586), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_632), .B(n_519), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_639), .A2(n_541), .B(n_614), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_657), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_635), .Y(n_681) );
OAI31xp33_ASAP7_75t_L g682 ( .A1(n_663), .A2(n_631), .A3(n_654), .B(n_638), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_667), .A2(n_646), .B1(n_654), .B2(n_641), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_658), .A2(n_644), .B1(n_621), .B2(n_622), .Y(n_684) );
OAI21xp33_ASAP7_75t_L g685 ( .A1(n_659), .A2(n_627), .B(n_622), .Y(n_685) );
AOI311xp33_ASAP7_75t_L g686 ( .A1(n_663), .A2(n_624), .A3(n_625), .B(n_649), .C(n_652), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_659), .A2(n_651), .B(n_620), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_662), .B(n_645), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_665), .A2(n_644), .B1(n_630), .B2(n_636), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_674), .A2(n_629), .B(n_650), .C(n_640), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_665), .A2(n_655), .B(n_618), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_661), .A2(n_651), .B(n_557), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_668), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g694 ( .A1(n_673), .A2(n_519), .B(n_613), .C(n_596), .Y(n_694) );
AOI321xp33_ASAP7_75t_L g695 ( .A1(n_664), .A2(n_607), .A3(n_610), .B1(n_609), .B2(n_608), .C(n_606), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_693), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_690), .B(n_676), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_683), .A2(n_672), .B(n_679), .C(n_670), .Y(n_698) );
OAI21xp33_ASAP7_75t_SL g699 ( .A1(n_682), .A2(n_670), .B(n_678), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_685), .B(n_660), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_683), .A2(n_677), .B(n_681), .Y(n_701) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_687), .A2(n_671), .A3(n_666), .B1(n_675), .B2(n_669), .C1(n_680), .C2(n_566), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g703 ( .A1(n_689), .A2(n_612), .B(n_605), .Y(n_703) );
NAND3x1_ASAP7_75t_L g704 ( .A(n_700), .B(n_686), .C(n_692), .Y(n_704) );
NOR3xp33_ASAP7_75t_SL g705 ( .A(n_699), .B(n_691), .C(n_684), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_701), .A2(n_694), .B(n_688), .C(n_695), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_698), .B(n_612), .C(n_605), .Y(n_707) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_702), .B(n_597), .C(n_555), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_705), .B(n_696), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_704), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_707), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_710), .B(n_697), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
OAI22xp33_ASAP7_75t_SL g715 ( .A1(n_714), .A2(n_713), .B1(n_709), .B2(n_712), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_706), .B(n_708), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_703), .B1(n_519), .B2(n_552), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_524), .B(n_540), .Y(n_718) );
OAI21x1_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_524), .B(n_540), .Y(n_719) );
AO21x2_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_540), .B(n_544), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_552), .B1(n_548), .B2(n_544), .Y(n_721) );
endmodule