module fake_netlist_5_155_n_1736 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1736);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1736;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_88),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_30),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_95),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_32),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_27),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_32),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_34),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_60),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_47),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_57),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_109),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_28),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_2),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_58),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_36),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_92),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_54),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_48),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_117),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_33),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_86),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_102),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_38),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_97),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_48),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_113),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_15),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_127),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_53),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_99),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_85),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_72),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_105),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_24),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_52),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_11),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_118),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_39),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_31),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_67),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_100),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_74),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_110),
.Y(n_247)
);

BUFx8_ASAP7_75t_SL g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_133),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_75),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_28),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_77),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_68),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_155),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_34),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_121),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_31),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_98),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_130),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_103),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_101),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_83),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_125),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_106),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_131),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_23),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_20),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_81),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_20),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_19),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_69),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_104),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_120),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_145),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_40),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_153),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_142),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_71),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_13),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_52),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_108),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_42),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_46),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_116),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_93),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_96),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_62),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_4),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_73),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_56),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_90),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_12),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_205),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_248),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_168),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_220),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_222),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_231),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_157),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_203),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_222),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_214),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_159),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_169),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_214),
.Y(n_329)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_169),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_171),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_160),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_171),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_179),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_165),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_179),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_180),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_180),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_203),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_156),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_166),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_208),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_208),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_163),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_206),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_161),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_237),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_172),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_173),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_178),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_290),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_181),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_280),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_200),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_164),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_294),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_186),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_187),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_158),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_327),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_221),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_333),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_329),
.A2(n_277),
.B1(n_286),
.B2(n_242),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_342),
.A2(n_308),
.B(n_297),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_270),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_311),
.A2(n_321),
.B1(n_357),
.B2(n_319),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_371),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_348),
.B(n_309),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_314),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_312),
.B(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

CKINVDCx11_ASAP7_75t_R g405 ( 
.A(n_374),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_315),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_188),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_315),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_354),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_317),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_356),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

OR2x6_ASAP7_75t_L g425 ( 
.A(n_330),
.B(n_221),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_359),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_375),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_318),
.Y(n_429)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_379),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_323),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_378),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_323),
.A2(n_162),
.B(n_161),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_339),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_324),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_339),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_340),
.B(n_190),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g442 ( 
.A(n_313),
.B(n_191),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_344),
.B(n_194),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_326),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_395),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_395),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_SL g456 ( 
.A(n_392),
.B(n_170),
.C(n_167),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_393),
.A2(n_212),
.B1(n_297),
.B2(n_308),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_279),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_411),
.Y(n_462)
);

BUFx6f_ASAP7_75t_SL g463 ( 
.A(n_425),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_346),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_393),
.A2(n_162),
.B1(n_232),
.B2(n_230),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_279),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_192),
.C(n_183),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_402),
.Y(n_480)
);

NOR2x1p5_ASAP7_75t_L g481 ( 
.A(n_427),
.B(n_212),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_404),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_393),
.A2(n_292),
.B1(n_350),
.B2(n_264),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_398),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_389),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_388),
.B(n_325),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_400),
.B(n_174),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_397),
.A2(n_292),
.B1(n_238),
.B2(n_197),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_287),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_195),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_400),
.B(n_174),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_420),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_400),
.B(n_174),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_397),
.A2(n_238),
.B1(n_192),
.B2(n_196),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_195),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_434),
.B(n_196),
.C(n_183),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_433),
.A2(n_243),
.B1(n_229),
.B2(n_310),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_410),
.B(n_209),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_425),
.B(n_330),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_423),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_198),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

NOR2x1p5_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_175),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_425),
.A2(n_227),
.B1(n_226),
.B2(n_306),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_417),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_410),
.B(n_209),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_388),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_433),
.A2(n_189),
.B1(n_185),
.B2(n_182),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_418),
.B(n_345),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_422),
.B(n_347),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_445),
.B(n_204),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_434),
.A2(n_230),
.B1(n_301),
.B2(n_291),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_410),
.B(n_258),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_424),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_434),
.A2(n_232),
.B1(n_235),
.B2(n_223),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_410),
.B(n_176),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_429),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_429),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_425),
.B(n_197),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_427),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_419),
.B(n_177),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_435),
.B(n_210),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_429),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_430),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_435),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_446),
.A2(n_269),
.B1(n_223),
.B2(n_219),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_440),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_439),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_443),
.B(n_207),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_440),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_444),
.B(n_211),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_419),
.B(n_209),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_419),
.B(n_426),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_447),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_430),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_430),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_412),
.B(n_347),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_419),
.B(n_428),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_431),
.B(n_250),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_430),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_430),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_412),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_403),
.A2(n_268),
.B(n_201),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_412),
.B(n_193),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_446),
.A2(n_235),
.B1(n_301),
.B2(n_291),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_412),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_440),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_442),
.B(n_250),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_399),
.B(n_207),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_440),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_413),
.A2(n_219),
.B1(n_217),
.B2(n_275),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_413),
.B(n_215),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_533),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_541),
.B(n_413),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_462),
.B(n_413),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_529),
.A2(n_498),
.B1(n_516),
.B2(n_550),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_499),
.B(n_199),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_529),
.A2(n_216),
.B1(n_225),
.B2(n_228),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_535),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_464),
.B(n_432),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_448),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_432),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_455),
.B(n_398),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_559),
.B(n_521),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_466),
.A2(n_245),
.B(n_244),
.C(n_254),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_536),
.B(n_432),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_535),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_530),
.B(n_195),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_458),
.B(n_471),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_202),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_530),
.B(n_195),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_503),
.B(n_213),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_530),
.B(n_195),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_506),
.B(n_218),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_498),
.B(n_261),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_539),
.A2(n_249),
.B1(n_233),
.B2(n_234),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_554),
.B(n_572),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_448),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_498),
.A2(n_217),
.B1(n_244),
.B2(n_245),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_432),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_473),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_473),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_468),
.A2(n_438),
.B(n_437),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_474),
.B(n_254),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_549),
.A2(n_262),
.B1(n_264),
.B2(n_269),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_448),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_516),
.B(n_491),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_516),
.B(n_351),
.Y(n_635)
);

BUFx5_ASAP7_75t_L g636 ( 
.A(n_585),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_551),
.B(n_241),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_450),
.A2(n_276),
.B(n_275),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_551),
.B(n_247),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_477),
.B(n_262),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_466),
.B(n_585),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_479),
.B(n_276),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_449),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_449),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_483),
.B(n_267),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_483),
.B(n_408),
.Y(n_647)
);

BUFx5_ASAP7_75t_L g648 ( 
.A(n_589),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_351),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_484),
.B(n_408),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_484),
.B(n_408),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_589),
.B(n_261),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_452),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_492),
.B(n_409),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_492),
.B(n_496),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_452),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_496),
.B(n_409),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_500),
.B(n_409),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_481),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_481),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_550),
.A2(n_285),
.B1(n_253),
.B2(n_255),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_500),
.B(n_414),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_453),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_456),
.B(n_224),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_567),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_502),
.B(n_414),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_524),
.B(n_236),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_453),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_459),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_459),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_469),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_476),
.A2(n_261),
.B1(n_382),
.B2(n_377),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_508),
.B(n_414),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_517),
.B(n_261),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_525),
.B(n_421),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_545),
.B(n_239),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_525),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_515),
.A2(n_274),
.B1(n_271),
.B2(n_272),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_527),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_552),
.B(n_240),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_518),
.B(n_252),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_469),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_526),
.B(n_256),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_520),
.B(n_250),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_531),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_421),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_485),
.B(n_451),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_550),
.A2(n_307),
.B1(n_305),
.B2(n_303),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_454),
.A2(n_438),
.B(n_437),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_538),
.B(n_421),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_550),
.A2(n_265),
.B1(n_283),
.B2(n_263),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_538),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_451),
.B(n_163),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_451),
.B(n_163),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_540),
.B(n_257),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_573),
.B(n_273),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_540),
.B(n_281),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_470),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_L g703 ( 
.A1(n_515),
.A2(n_532),
.B1(n_550),
.B2(n_461),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_438),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_546),
.B(n_261),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_562),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_562),
.B(n_437),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_476),
.A2(n_382),
.B1(n_377),
.B2(n_376),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_470),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_507),
.B(n_376),
.C(n_373),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_298),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_563),
.B(n_284),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_523),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_564),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_472),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_569),
.B(n_373),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_564),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_507),
.B(n_372),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_372),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_451),
.B(n_370),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_566),
.B(n_568),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_472),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_568),
.B(n_0),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_571),
.B(n_575),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_465),
.B(n_370),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_567),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_523),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_575),
.B(n_369),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_569),
.B(n_369),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_509),
.A2(n_368),
.B1(n_367),
.B2(n_366),
.C(n_363),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_512),
.A2(n_368),
.B1(n_367),
.B2(n_366),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_475),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_586),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_586),
.A2(n_363),
.B1(n_362),
.B2(n_361),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_497),
.A2(n_362),
.B1(n_361),
.B2(n_360),
.C(n_358),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_576),
.B(n_586),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_579),
.B(n_360),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_465),
.B(n_358),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_475),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_537),
.B(n_353),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_579),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_488),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_581),
.B(n_0),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_595),
.B(n_353),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_488),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_457),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_465),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_591),
.B(n_1),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_457),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_544),
.B(n_352),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_352),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_557),
.B(n_148),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_457),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_457),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_574),
.B(n_2),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_519),
.B(n_141),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_584),
.B(n_577),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_584),
.B(n_135),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_488),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_577),
.B(n_134),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_578),
.B(n_119),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_622),
.A2(n_463),
.B1(n_461),
.B2(n_580),
.Y(n_765)
);

AND2x6_ASAP7_75t_SL g766 ( 
.A(n_664),
.B(n_592),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_635),
.Y(n_767)
);

NOR2x1p5_ASAP7_75t_L g768 ( 
.A(n_607),
.B(n_465),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_678),
.A2(n_463),
.B1(n_461),
.B2(n_489),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_744),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_665),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_601),
.B(n_490),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_678),
.A2(n_512),
.B(n_532),
.C(n_561),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_693),
.A2(n_553),
.B(n_547),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_721),
.B(n_490),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_744),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_683),
.A2(n_463),
.B1(n_461),
.B2(n_501),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_634),
.B(n_519),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_665),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_490),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_612),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_635),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_624),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_726),
.B(n_490),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_612),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_717),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_741),
.B(n_511),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_505),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_634),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_613),
.A2(n_618),
.B(n_616),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_SL g793 ( 
.A1(n_638),
.A2(n_461),
.B(n_519),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_683),
.B(n_487),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_703),
.B(n_511),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_664),
.B(n_511),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_703),
.B(n_665),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_608),
.B(n_597),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_614),
.B(n_505),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_731),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_633),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_665),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_750),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_699),
.Y(n_804)
);

AND2x6_ASAP7_75t_L g805 ( 
.A(n_759),
.B(n_522),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_511),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_680),
.B(n_588),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_655),
.B(n_722),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_649),
.B(n_519),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_645),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_649),
.B(n_519),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_680),
.B(n_460),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_680),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_758),
.A2(n_510),
.B1(n_594),
.B2(n_592),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_643),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_596),
.B(n_598),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_758),
.A2(n_592),
.B1(n_578),
.B2(n_582),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_691),
.B(n_592),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_719),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_672),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_603),
.B(n_592),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_680),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_644),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_710),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_631),
.A2(n_582),
.B1(n_590),
.B2(n_583),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_697),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_653),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_667),
.B(n_615),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_631),
.A2(n_611),
.B1(n_746),
.B2(n_673),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_710),
.B(n_547),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_615),
.B(n_478),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_659),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_660),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_711),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_725),
.B(n_542),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_747),
.B(n_542),
.Y(n_837)
);

BUFx4f_ASAP7_75t_L g838 ( 
.A(n_759),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_710),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_676),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_710),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_750),
.B(n_505),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_728),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_714),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_729),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_679),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_687),
.A2(n_619),
.B(n_617),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_701),
.B(n_712),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_682),
.B(n_542),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_688),
.B(n_542),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_728),
.A2(n_534),
.B1(n_590),
.B2(n_583),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_701),
.B(n_712),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_689),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_696),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_728),
.A2(n_528),
.B1(n_570),
.B2(n_565),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_711),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_706),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_728),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_715),
.B(n_505),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_698),
.B(n_534),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_718),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_513),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_746),
.A2(n_528),
.B1(n_570),
.B2(n_565),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_733),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_707),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_745),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_684),
.B(n_480),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_641),
.B(n_547),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_673),
.A2(n_480),
.B1(n_560),
.B2(n_558),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_730),
.B(n_504),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_755),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_647),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_650),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_684),
.B(n_504),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_613),
.B(n_513),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_600),
.A2(n_495),
.B1(n_560),
.B2(n_558),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_651),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_736),
.B(n_513),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_681),
.A2(n_482),
.B1(n_556),
.B2(n_555),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_713),
.B(n_3),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_616),
.B(n_513),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_617),
.B(n_547),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_686),
.A2(n_486),
.B1(n_556),
.B2(n_555),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_630),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_751),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_713),
.B(n_3),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_686),
.B(n_482),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_654),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_751),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_619),
.B(n_4),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_720),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_700),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_700),
.B(n_486),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_761),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_SL g896 ( 
.A(n_661),
.B(n_493),
.C(n_495),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_657),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_618),
.B(n_548),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_640),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_740),
.A2(n_548),
.B1(n_543),
.B2(n_514),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_658),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_730),
.B(n_543),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_637),
.B(n_514),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_662),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_636),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_642),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_753),
.A2(n_493),
.B1(n_522),
.B2(n_593),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_724),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_666),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_674),
.Y(n_910)
);

AO22x1_ASAP7_75t_L g911 ( 
.A1(n_724),
.A2(n_593),
.B1(n_522),
.B2(n_10),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_739),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_663),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_737),
.B(n_604),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_677),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_748),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_646),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_668),
.Y(n_918)
);

NAND2x1_ASAP7_75t_L g919 ( 
.A(n_605),
.B(n_553),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_621),
.B(n_593),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_610),
.A2(n_553),
.B1(n_467),
.B2(n_115),
.Y(n_921)
);

OR2x2_ASAP7_75t_SL g922 ( 
.A(n_681),
.B(n_5),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_636),
.B(n_553),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_636),
.B(n_467),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_636),
.B(n_467),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_R g926 ( 
.A(n_754),
.B(n_111),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_669),
.Y(n_927)
);

BUFx5_ASAP7_75t_L g928 ( 
.A(n_749),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_743),
.A2(n_467),
.B1(n_10),
.B2(n_12),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_636),
.B(n_467),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_762),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_670),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_636),
.B(n_467),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_690),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_763),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_623),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_639),
.B(n_107),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_694),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_692),
.B(n_7),
.Y(n_939)
);

NAND2x1_ASAP7_75t_L g940 ( 
.A(n_632),
.B(n_94),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_648),
.B(n_752),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_641),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_648),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_732),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_648),
.B(n_78),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_648),
.B(n_7),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_648),
.B(n_14),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_671),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_648),
.B(n_14),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_602),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_905),
.A2(n_606),
.B(n_599),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_813),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_770),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_905),
.A2(n_760),
.B(n_757),
.Y(n_954)
);

OAI22x1_ASAP7_75t_L g955 ( 
.A1(n_828),
.A2(n_695),
.B1(n_620),
.B2(n_743),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_771),
.B(n_620),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_912),
.B(n_756),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_848),
.B(n_626),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_923),
.A2(n_764),
.B(n_704),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_774),
.A2(n_629),
.B(n_702),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_893),
.B(n_625),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_912),
.B(n_742),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_783),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_923),
.A2(n_709),
.B(n_735),
.Y(n_964)
);

AOI22x1_ASAP7_75t_L g965 ( 
.A1(n_852),
.A2(n_685),
.B1(n_723),
.B2(n_716),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_773),
.A2(n_734),
.B1(n_708),
.B2(n_738),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_778),
.B(n_609),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_808),
.A2(n_652),
.B(n_705),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_808),
.A2(n_652),
.B(n_705),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_847),
.A2(n_675),
.B(n_734),
.C(n_708),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_943),
.A2(n_675),
.B(n_66),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_776),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_798),
.B(n_16),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_813),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_789),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_943),
.A2(n_65),
.B(n_18),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_797),
.A2(n_794),
.B(n_795),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_942),
.B(n_16),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_788),
.A2(n_792),
.B(n_812),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_908),
.B(n_21),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_813),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_772),
.B(n_22),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_780),
.B(n_22),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_829),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_891),
.A2(n_887),
.B(n_881),
.C(n_806),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_839),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_781),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_942),
.B(n_26),
.Y(n_988)
);

BUFx8_ASAP7_75t_L g989 ( 
.A(n_804),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_781),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_829),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_796),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_873),
.B(n_39),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_788),
.A2(n_40),
.B(n_42),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_791),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_874),
.B(n_43),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_807),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_839),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_792),
.A2(n_49),
.B(n_50),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_771),
.A2(n_51),
.B(n_799),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_878),
.B(n_51),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_886),
.A2(n_856),
.B(n_835),
.C(n_890),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_786),
.Y(n_1003)
);

INVx3_ASAP7_75t_SL g1004 ( 
.A(n_803),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_914),
.B(n_872),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_945),
.A2(n_946),
.B(n_949),
.C(n_947),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_SL g1007 ( 
.A1(n_883),
.A2(n_777),
.B(n_765),
.C(n_769),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_801),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_838),
.A2(n_950),
.B1(n_818),
.B2(n_805),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_944),
.A2(n_937),
.B1(n_816),
.B2(n_892),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_826),
.B(n_821),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_810),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_937),
.A2(n_816),
.B1(n_790),
.B2(n_899),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_793),
.A2(n_838),
.B(n_814),
.C(n_885),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_785),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_815),
.Y(n_1016)
);

CKINVDCx8_ASAP7_75t_R g1017 ( 
.A(n_766),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_844),
.B(n_832),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_826),
.B(n_800),
.Y(n_1019)
);

CKINVDCx14_ASAP7_75t_R g1020 ( 
.A(n_842),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_839),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_819),
.B(n_861),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_778),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_820),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_906),
.B(n_889),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_917),
.B(n_775),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_898),
.A2(n_869),
.B(n_907),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_817),
.A2(n_904),
.B(n_897),
.C(n_910),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_784),
.B(n_787),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_771),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_821),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_823),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_827),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_771),
.A2(n_836),
.B(n_799),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_767),
.B(n_782),
.C(n_939),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_830),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_809),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_840),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_929),
.A2(n_860),
.B(n_853),
.C(n_846),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_809),
.B(n_811),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_802),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_913),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_SL g1043 ( 
.A1(n_854),
.A2(n_864),
.B(n_857),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_867),
.A2(n_894),
.B(n_875),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_845),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_811),
.B(n_802),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_822),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_768),
.B(n_833),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_836),
.A2(n_925),
.B(n_933),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_916),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_901),
.A2(n_938),
.B(n_934),
.C(n_909),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_922),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_834),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_927),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_824),
.B(n_841),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_915),
.B(n_865),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_929),
.A2(n_888),
.B(n_825),
.C(n_837),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_932),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_924),
.A2(n_933),
.B(n_925),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_841),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_849),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_870),
.B(n_837),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_SL g1064 ( 
.A(n_926),
.B(n_945),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_903),
.B(n_948),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_898),
.A2(n_869),
.B(n_907),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_924),
.A2(n_930),
.B(n_831),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_805),
.A2(n_903),
.B1(n_920),
.B2(n_779),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_916),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_SL g1070 ( 
.A(n_805),
.B(n_858),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_805),
.B(n_902),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_941),
.B(n_843),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_871),
.B(n_902),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_871),
.A2(n_921),
.B(n_877),
.C(n_876),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_930),
.A2(n_831),
.B(n_882),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_941),
.B(n_849),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_876),
.A2(n_882),
.B(n_868),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_850),
.B(n_862),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_866),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_948),
.B(n_936),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_825),
.A2(n_850),
.B(n_862),
.C(n_859),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_866),
.B(n_868),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_900),
.A2(n_880),
.B(n_884),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_928),
.B(n_911),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_948),
.B(n_936),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_948),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_863),
.B(n_896),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_919),
.A2(n_851),
.B(n_855),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_936),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_935),
.A2(n_872),
.B(n_895),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_872),
.B(n_895),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_895),
.B(n_935),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_936),
.B(n_935),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_951),
.A2(n_931),
.B(n_940),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1006),
.A2(n_931),
.B(n_879),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_990),
.B(n_928),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1020),
.Y(n_1097)
);

CKINVDCx11_ASAP7_75t_R g1098 ( 
.A(n_1004),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_958),
.B(n_928),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_928),
.B(n_931),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1010),
.A2(n_928),
.B1(n_931),
.B2(n_966),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_963),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1052),
.A2(n_982),
.B1(n_983),
.B2(n_977),
.Y(n_1103)
);

AOI221x1_ASAP7_75t_L g1104 ( 
.A1(n_999),
.A2(n_984),
.B1(n_991),
.B2(n_1000),
.C(n_955),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_975),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_987),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1014),
.A2(n_1074),
.A3(n_979),
.B(n_1077),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1067),
.A2(n_1075),
.B(n_1060),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_985),
.A2(n_1058),
.B(n_1039),
.C(n_1007),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1057),
.B(n_1051),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1003),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1008),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_964),
.A2(n_1049),
.B(n_1088),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_954),
.A2(n_1044),
.B(n_1034),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1045),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1025),
.B(n_1015),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_SL g1118 ( 
.A(n_1092),
.B(n_1018),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1057),
.B(n_1076),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1053),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1121)
);

AO21x1_ASAP7_75t_L g1122 ( 
.A1(n_1064),
.A2(n_1084),
.B(n_1083),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_966),
.A2(n_1013),
.B1(n_1028),
.B2(n_991),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_997),
.A2(n_980),
.B(n_992),
.Y(n_1124)
);

CKINVDCx6p67_ASAP7_75t_R g1125 ( 
.A(n_1048),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1063),
.B(n_957),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_959),
.A2(n_965),
.B(n_1090),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1070),
.A2(n_1083),
.B(n_1078),
.Y(n_1128)
);

AO22x1_ASAP7_75t_L g1129 ( 
.A1(n_984),
.A2(n_1019),
.B1(n_1026),
.B2(n_1005),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_957),
.B(n_1078),
.Y(n_1130)
);

OAI22x1_ASAP7_75t_L g1131 ( 
.A1(n_1035),
.A2(n_1009),
.B1(n_1011),
.B2(n_1068),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1040),
.B(n_1023),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1012),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1070),
.A2(n_968),
.B(n_969),
.Y(n_1134)
);

AO21x1_ASAP7_75t_L g1135 ( 
.A1(n_1084),
.A2(n_1087),
.B(n_973),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1072),
.B(n_962),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_SL g1137 ( 
.A1(n_961),
.A2(n_1027),
.B(n_1066),
.C(n_1065),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1081),
.A2(n_1027),
.B(n_1066),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_962),
.B(n_1073),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_1017),
.B(n_989),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1080),
.A2(n_1085),
.B(n_1091),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_971),
.A2(n_1071),
.B(n_1093),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_993),
.A2(n_996),
.B1(n_1001),
.B2(n_1024),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1082),
.A2(n_996),
.A3(n_993),
.B(n_1001),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1038),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1071),
.A2(n_956),
.B(n_970),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_956),
.A2(n_1056),
.B(n_1086),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1089),
.A2(n_1046),
.B(n_1043),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1055),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_994),
.A2(n_976),
.A3(n_988),
.B(n_978),
.Y(n_1150)
);

OAI22x1_ASAP7_75t_L g1151 ( 
.A1(n_1029),
.A2(n_988),
.B1(n_978),
.B2(n_1031),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_SL g1152 ( 
.A1(n_967),
.A2(n_1037),
.B1(n_1023),
.B2(n_1079),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1005),
.B(n_1061),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1002),
.B(n_1022),
.C(n_967),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_967),
.A2(n_1023),
.B1(n_1089),
.B2(n_1033),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1030),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1005),
.B(n_1061),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1016),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_989),
.B(n_953),
.C(n_972),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_1041),
.B(n_1047),
.C(n_1054),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1032),
.B(n_1036),
.Y(n_1161)
);

NAND3x1_ASAP7_75t_L g1162 ( 
.A(n_974),
.B(n_1050),
.C(n_1005),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_1050),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1042),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1030),
.B(n_952),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1059),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_974),
.A2(n_981),
.B(n_1050),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1069),
.B(n_952),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1030),
.A2(n_952),
.B(n_986),
.Y(n_1169)
);

INVx6_ASAP7_75t_SL g1170 ( 
.A(n_1021),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_986),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_986),
.A2(n_828),
.B1(n_848),
.B2(n_773),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_998),
.A2(n_905),
.B(n_951),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_998),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_SL g1175 ( 
.A1(n_998),
.A2(n_1014),
.B(n_905),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1021),
.B(n_912),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1021),
.A2(n_960),
.B(n_1067),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_990),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1030),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_963),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_990),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1030),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_963),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1025),
.B(n_828),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_990),
.B(n_781),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_990),
.B(n_828),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_979),
.A2(n_828),
.B(n_1027),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_985),
.A2(n_828),
.B(n_848),
.Y(n_1194)
);

AO22x2_ASAP7_75t_L g1195 ( 
.A1(n_984),
.A2(n_991),
.B1(n_795),
.B2(n_848),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_963),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_951),
.A2(n_905),
.B(n_1006),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1010),
.A2(n_828),
.B1(n_848),
.B2(n_773),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1040),
.B(n_1023),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_999),
.A2(n_828),
.B(n_982),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_951),
.A2(n_905),
.B(n_1006),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_958),
.B(n_912),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_951),
.A2(n_905),
.B(n_1006),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_951),
.A2(n_905),
.B(n_1006),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_977),
.A2(n_999),
.B(n_1039),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_958),
.B(n_912),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_985),
.A2(n_828),
.B(n_847),
.C(n_852),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1025),
.B(n_828),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_990),
.B(n_781),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_951),
.A2(n_905),
.B(n_1006),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1052),
.A2(n_828),
.B1(n_806),
.B2(n_795),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_963),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_990),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1034),
.A2(n_979),
.B(n_1049),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_977),
.A2(n_1014),
.A3(n_1074),
.B(n_979),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1030),
.B(n_771),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1027),
.A2(n_1066),
.B(n_1083),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_963),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1020),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1030),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_990),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_SL g1225 ( 
.A1(n_977),
.A2(n_999),
.B(n_1039),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_960),
.A2(n_1067),
.B(n_1075),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1040),
.B(n_1023),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1025),
.B(n_828),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_1007),
.A2(n_773),
.B(n_828),
.C(n_1014),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1010),
.A2(n_828),
.B1(n_848),
.B2(n_773),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_984),
.A2(n_991),
.B1(n_795),
.B2(n_848),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_958),
.B(n_912),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_958),
.B(n_912),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_958),
.B(n_912),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1010),
.A2(n_828),
.B1(n_806),
.B2(n_847),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1006),
.A2(n_905),
.B(n_951),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1191),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1204),
.A2(n_1212),
.B(n_1205),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1098),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1209),
.A2(n_1235),
.B(n_1194),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1122),
.A2(n_1135),
.A3(n_1200),
.B(n_1236),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1190),
.A2(n_1228),
.B1(n_1210),
.B2(n_1119),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1236),
.A2(n_1127),
.B(n_1100),
.Y(n_1245)
);

AOI222xp33_ASAP7_75t_L g1246 ( 
.A1(n_1124),
.A2(n_1230),
.B1(n_1198),
.B2(n_1193),
.C1(n_1123),
.C2(n_1231),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1193),
.A2(n_1134),
.B(n_1128),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1161),
.B(n_1117),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1229),
.A2(n_1119),
.B(n_1110),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1194),
.A2(n_1198),
.B(n_1230),
.C(n_1123),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1143),
.A2(n_1101),
.A3(n_1172),
.B(n_1151),
.Y(n_1251)
);

AOI222xp33_ASAP7_75t_L g1252 ( 
.A1(n_1195),
.A2(n_1231),
.B1(n_1213),
.B2(n_1192),
.C1(n_1143),
.C2(n_1172),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1101),
.A2(n_1095),
.A3(n_1131),
.B(n_1094),
.Y(n_1253)
);

AOI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_1195),
.A2(n_1103),
.B1(n_1206),
.B2(n_1225),
.C(n_1154),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1129),
.A2(n_1173),
.B(n_1216),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1137),
.A2(n_1146),
.B(n_1136),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1110),
.A2(n_1108),
.B(n_1175),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1178),
.A2(n_1201),
.B(n_1180),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1102),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1125),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1132),
.B(n_1199),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1112),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_1208),
.B(n_1226),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1211),
.B(n_1106),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1185),
.B(n_1181),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1140),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1183),
.A2(n_1222),
.B(n_1187),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1132),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1203),
.A2(n_1207),
.B1(n_1234),
.B2(n_1232),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1188),
.A2(n_1115),
.B(n_1114),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_1116),
.B(n_1215),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1142),
.A2(n_1148),
.B(n_1147),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1113),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1099),
.A2(n_1155),
.B(n_1153),
.Y(n_1274)
);

AND2x6_ASAP7_75t_L g1275 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1219),
.A2(n_1234),
.B1(n_1233),
.B2(n_1232),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1219),
.A2(n_1233),
.B1(n_1139),
.B2(n_1152),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1224),
.B(n_1139),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1121),
.A2(n_1130),
.B(n_1136),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1118),
.A2(n_1199),
.B1(n_1227),
.B2(n_1159),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1227),
.B(n_1145),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1126),
.B(n_1223),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1141),
.A2(n_1126),
.B(n_1160),
.Y(n_1283)
);

AND2x2_ASAP7_75t_SL g1284 ( 
.A(n_1120),
.B(n_1096),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1176),
.A2(n_1167),
.B(n_1166),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1163),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1149),
.A2(n_1164),
.B1(n_1158),
.B2(n_1220),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1182),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1162),
.A2(n_1169),
.B(n_1218),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1156),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1105),
.Y(n_1291)
);

CKINVDCx9p33_ASAP7_75t_R g1292 ( 
.A(n_1168),
.Y(n_1292)
);

AOI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1165),
.A2(n_1214),
.B(n_1196),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1218),
.A2(n_1184),
.B(n_1111),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_SL g1295 ( 
.A1(n_1133),
.A2(n_1189),
.B(n_1171),
.C(n_1174),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1168),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1182),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1144),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1156),
.Y(n_1299)
);

AND2x2_ASAP7_75t_SL g1300 ( 
.A(n_1217),
.B(n_1223),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1144),
.Y(n_1301)
);

AOI211xp5_ASAP7_75t_L g1302 ( 
.A1(n_1097),
.A2(n_1221),
.B(n_1150),
.C(n_1186),
.Y(n_1302)
);

OAI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_1150),
.B1(n_1144),
.B2(n_1217),
.C(n_1107),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1150),
.A2(n_1107),
.B(n_1170),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1170),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1107),
.B(n_828),
.C(n_780),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1175),
.B(n_1152),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1209),
.A2(n_1007),
.B(n_828),
.C(n_773),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1190),
.A2(n_828),
.B1(n_806),
.B2(n_848),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1236),
.A2(n_1202),
.B(n_1197),
.Y(n_1312)
);

BUFx2_ASAP7_75t_R g1313 ( 
.A(n_1097),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1120),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1095),
.A2(n_1202),
.B(n_1197),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1194),
.B(n_828),
.C(n_780),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1102),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1194),
.A2(n_828),
.B1(n_852),
.B2(n_848),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1102),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1162),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1122),
.A2(n_1135),
.A3(n_1200),
.B(n_1109),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1095),
.A2(n_1202),
.B(n_1197),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1191),
.B(n_1211),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1191),
.B(n_1211),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1191),
.B(n_1211),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1209),
.A2(n_828),
.B(n_852),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1194),
.A2(n_828),
.B1(n_852),
.B2(n_848),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1102),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1132),
.B(n_1199),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1102),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1138),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1162),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1138),
.A2(n_1193),
.B(n_1197),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1102),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1190),
.B(n_1210),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1122),
.A2(n_1135),
.A3(n_1200),
.B(n_1109),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1224),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1197),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1156),
.Y(n_1357)
);

AOI22x1_ASAP7_75t_L g1358 ( 
.A1(n_1213),
.A2(n_848),
.B1(n_852),
.B2(n_1131),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1244),
.B(n_1316),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1311),
.A2(n_1328),
.B1(n_1319),
.B2(n_1342),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1278),
.B(n_1248),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1281),
.B(n_1261),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1355),
.B(n_1286),
.Y(n_1363)
);

INVx4_ASAP7_75t_SL g1364 ( 
.A(n_1308),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1351),
.A2(n_1257),
.B(n_1247),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1291),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1268),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1318),
.A2(n_1330),
.B1(n_1336),
.B2(n_1325),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1343),
.B(n_1353),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1340),
.A2(n_1241),
.B(n_1322),
.C(n_1256),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1306),
.A2(n_1312),
.B(n_1249),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1345),
.A2(n_1326),
.B1(n_1341),
.B2(n_1284),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1326),
.A2(n_1341),
.B1(n_1284),
.B2(n_1280),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1339),
.B(n_1264),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1308),
.A2(n_1283),
.B(n_1250),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1269),
.B(n_1237),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1281),
.B(n_1346),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1296),
.B(n_1265),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1315),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1277),
.A2(n_1308),
.B1(n_1302),
.B2(n_1350),
.Y(n_1381)
);

INVx3_ASAP7_75t_SL g1382 ( 
.A(n_1305),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_SL g1383 ( 
.A1(n_1309),
.A2(n_1358),
.B(n_1246),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1329),
.B(n_1350),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1279),
.A2(n_1254),
.B(n_1239),
.C(n_1277),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1329),
.A2(n_1287),
.B1(n_1262),
.B2(n_1282),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1344),
.B(n_1276),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_L g1388 ( 
.A(n_1259),
.B(n_1273),
.Y(n_1388)
);

AOI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1309),
.A2(n_1292),
.B(n_1307),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1287),
.A2(n_1276),
.B1(n_1271),
.B2(n_1242),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1242),
.A2(n_1307),
.B1(n_1323),
.B2(n_1348),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1304),
.A2(n_1303),
.B(n_1285),
.C(n_1242),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1321),
.A2(n_1335),
.B(n_1323),
.C(n_1333),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1321),
.A2(n_1335),
.B(n_1333),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1274),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1347),
.B(n_1352),
.Y(n_1397)
);

O2A1O1Ixp5_ASAP7_75t_L g1398 ( 
.A1(n_1255),
.A2(n_1332),
.B(n_1317),
.C(n_1298),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1240),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1293),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1238),
.A2(n_1337),
.B(n_1320),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1321),
.A2(n_1348),
.B1(n_1335),
.B2(n_1333),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1310),
.A2(n_1337),
.B(n_1320),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1301),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1295),
.A2(n_1274),
.B1(n_1268),
.B2(n_1252),
.C(n_1240),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1314),
.A2(n_1349),
.B(n_1356),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1295),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1251),
.B(n_1331),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1294),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1312),
.A2(n_1348),
.B(n_1356),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1268),
.A2(n_1305),
.B1(n_1357),
.B2(n_1299),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1266),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1288),
.A2(n_1297),
.B(n_1267),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1275),
.B(n_1251),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1331),
.A2(n_1354),
.B(n_1253),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1314),
.A2(n_1349),
.B(n_1245),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1290),
.B(n_1288),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1297),
.A2(n_1267),
.B(n_1313),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1331),
.A2(n_1354),
.B(n_1253),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1300),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1245),
.A2(n_1270),
.B(n_1263),
.Y(n_1421)
);

NOR2xp67_ASAP7_75t_L g1422 ( 
.A(n_1260),
.B(n_1299),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1357),
.A2(n_1266),
.B1(n_1260),
.B2(n_1275),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1275),
.B(n_1354),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1275),
.B(n_1354),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1275),
.B(n_1331),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1357),
.B(n_1243),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1258),
.A2(n_1267),
.B(n_1253),
.C(n_1243),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1243),
.B(n_1253),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1258),
.A2(n_1289),
.B(n_1272),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1270),
.A2(n_1263),
.B1(n_828),
.B2(n_1311),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1311),
.A2(n_828),
.B(n_1194),
.C(n_1209),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1311),
.A2(n_828),
.B(n_806),
.C(n_1138),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1244),
.B(n_1316),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1278),
.B(n_1248),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1291),
.Y(n_1437)
);

O2A1O1Ixp5_ASAP7_75t_L g1438 ( 
.A1(n_1311),
.A2(n_1200),
.B(n_828),
.C(n_1351),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1278),
.B(n_1248),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1404),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1400),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1394),
.A2(n_1410),
.B(n_1372),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1377),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1360),
.B(n_1367),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1437),
.B(n_1359),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1379),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1407),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1366),
.A2(n_1394),
.B(n_1395),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1391),
.A2(n_1402),
.B(n_1385),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1421),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1433),
.A2(n_1432),
.B(n_1385),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1409),
.B(n_1425),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1396),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1396),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1398),
.A2(n_1438),
.B(n_1371),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1387),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1414),
.B(n_1424),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1429),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1433),
.A2(n_1392),
.B(n_1428),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1420),
.B(n_1426),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1430),
.B(n_1413),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1408),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1392),
.B(n_1427),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1438),
.A2(n_1371),
.B(n_1431),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1390),
.A2(n_1376),
.B(n_1388),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1416),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_1373),
.B(n_1381),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1401),
.A2(n_1403),
.B(n_1406),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1393),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1397),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1406),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1375),
.B(n_1439),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1361),
.B(n_1440),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1365),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1435),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1436),
.B(n_1362),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1364),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1464),
.B(n_1380),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1464),
.B(n_1405),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1462),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1451),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1458),
.Y(n_1483)
);

OR2x2_ASAP7_75t_SL g1484 ( 
.A(n_1465),
.B(n_1368),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1464),
.B(n_1364),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1463),
.B(n_1386),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1454),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1451),
.B(n_1364),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1454),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1441),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1445),
.B(n_1444),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1441),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1452),
.A2(n_1369),
.B1(n_1370),
.B2(n_1418),
.C(n_1423),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1462),
.B(n_1378),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1463),
.B(n_1368),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1455),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1453),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1468),
.A2(n_1383),
.B1(n_1389),
.B2(n_1384),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1469),
.A2(n_1419),
.B(n_1415),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1453),
.Y(n_1500)
);

BUFx10_ASAP7_75t_L g1501 ( 
.A(n_1491),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1490),
.Y(n_1502)
);

INVx5_ASAP7_75t_L g1503 ( 
.A(n_1494),
.Y(n_1503)
);

AOI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1480),
.A2(n_1445),
.B1(n_1444),
.B2(n_1468),
.C(n_1457),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1495),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1491),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1475),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1490),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1498),
.A2(n_1465),
.B(n_1457),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1499),
.A2(n_1469),
.B(n_1472),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1493),
.A2(n_1498),
.B1(n_1480),
.B2(n_1465),
.C(n_1422),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1480),
.A2(n_1468),
.B1(n_1466),
.B2(n_1460),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1478),
.B(n_1453),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1493),
.A2(n_1468),
.B1(n_1466),
.B2(n_1460),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1497),
.Y(n_1515)
);

OAI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1480),
.A2(n_1465),
.B1(n_1446),
.B2(n_1447),
.C(n_1476),
.Y(n_1516)
);

AOI222xp33_ASAP7_75t_L g1517 ( 
.A1(n_1479),
.A2(n_1476),
.B1(n_1475),
.B2(n_1447),
.C1(n_1446),
.C2(n_1399),
.Y(n_1517)
);

OAI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1486),
.A2(n_1465),
.B(n_1456),
.C(n_1443),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1486),
.A2(n_1465),
.B1(n_1473),
.B2(n_1462),
.C(n_1411),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1483),
.A2(n_1468),
.B1(n_1470),
.B2(n_1471),
.C(n_1460),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1495),
.Y(n_1521)
);

AOI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1483),
.A2(n_1471),
.B1(n_1470),
.B2(n_1460),
.C(n_1461),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1485),
.A2(n_1466),
.B1(n_1478),
.B2(n_1460),
.Y(n_1523)
);

OAI31xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1485),
.A2(n_1477),
.A3(n_1474),
.B(n_1461),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1485),
.A2(n_1466),
.B1(n_1473),
.B2(n_1453),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1482),
.A2(n_1472),
.B(n_1467),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_1459),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

AND2x6_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1384),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1479),
.B(n_1473),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1481),
.A2(n_1466),
.B1(n_1449),
.B2(n_1450),
.Y(n_1532)
);

AOI211xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1488),
.A2(n_1417),
.B(n_1363),
.C(n_1448),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1492),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1497),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_L g1536 ( 
.A(n_1495),
.B(n_1461),
.C(n_1442),
.D(n_1471),
.Y(n_1536)
);

NOR2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1536),
.B(n_1481),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1487),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1504),
.B(n_1489),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1497),
.Y(n_1541)
);

AND2x2_ASAP7_75t_SL g1542 ( 
.A(n_1512),
.B(n_1481),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

INVx6_ASAP7_75t_L g1544 ( 
.A(n_1503),
.Y(n_1544)
);

INVx4_ASAP7_75t_SL g1545 ( 
.A(n_1529),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1528),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1531),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1529),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1534),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1527),
.Y(n_1552)
);

AO21x1_ASAP7_75t_L g1553 ( 
.A1(n_1514),
.A2(n_1496),
.B(n_1492),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1527),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1510),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1529),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1505),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1521),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1506),
.B(n_1489),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1530),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1501),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1501),
.Y(n_1564)
);

NOR2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1515),
.B(n_1481),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1547),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1538),
.B(n_1540),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1549),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1544),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1539),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1543),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1548),
.B(n_1500),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1540),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1564),
.B(n_1382),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1548),
.B(n_1535),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1548),
.B(n_1535),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1543),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1532),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1563),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1553),
.A2(n_1518),
.B(n_1509),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1546),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1552),
.B(n_1522),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_1511),
.B1(n_1520),
.B2(n_1509),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1507),
.Y(n_1589)
);

NAND4xp75_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1456),
.C(n_1511),
.D(n_1443),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1545),
.B(n_1478),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1551),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1551),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1560),
.B(n_1559),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.B(n_1525),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1539),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1559),
.B(n_1484),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1575),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1588),
.A2(n_1519),
.B(n_1517),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1569),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1581),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1583),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1587),
.B(n_1597),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1561),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_L g1612 ( 
.A(n_1574),
.B(n_1563),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1568),
.B(n_1561),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1581),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1597),
.B(n_1562),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1597),
.B(n_1562),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1558),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1588),
.A2(n_1542),
.B1(n_1537),
.B2(n_1519),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1574),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1585),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1569),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1578),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1550),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1589),
.B(n_1558),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1550),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1566),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1577),
.B(n_1558),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1577),
.B(n_1557),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1592),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1556),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1566),
.B(n_1553),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1626),
.B(n_1598),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1636),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1630),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1584),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1619),
.A2(n_1542),
.B1(n_1584),
.B2(n_1609),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1567),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1611),
.B(n_1567),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1630),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1582),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1570),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

AND2x2_ASAP7_75t_SL g1651 ( 
.A(n_1623),
.B(n_1578),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1635),
.B(n_1591),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1602),
.B(n_1604),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1636),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1635),
.A2(n_1584),
.B1(n_1591),
.B2(n_1586),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1603),
.A2(n_1584),
.B1(n_1591),
.B2(n_1586),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1576),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1620),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1615),
.B(n_1576),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1605),
.B(n_1412),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1637),
.B(n_1613),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1653),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1641),
.A2(n_1590),
.B1(n_1615),
.B2(n_1599),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1653),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1659),
.Y(n_1667)
);

BUFx2_ASAP7_75t_SL g1668 ( 
.A(n_1653),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1640),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1610),
.C(n_1555),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1642),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1653),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1645),
.B(n_1616),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1659),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1651),
.A2(n_1599),
.B1(n_1591),
.B2(n_1572),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1651),
.A2(n_1599),
.B1(n_1591),
.B2(n_1572),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1661),
.A2(n_1601),
.B(n_1586),
.C(n_1572),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1651),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1647),
.A2(n_1601),
.B(n_1629),
.C(n_1632),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1679),
.A2(n_1649),
.B1(n_1646),
.B2(n_1645),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1669),
.Y(n_1683)
);

INVxp33_ASAP7_75t_L g1684 ( 
.A(n_1674),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1677),
.B(n_1646),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1679),
.B(n_1646),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1672),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1667),
.B(n_1647),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1675),
.B(n_1649),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1666),
.B(n_1642),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1664),
.A2(n_1649),
.B1(n_1652),
.B2(n_1660),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1686),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1688),
.A2(n_1656),
.B1(n_1657),
.B2(n_1680),
.C(n_1678),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1691),
.A2(n_1671),
.B(n_1662),
.C(n_1654),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1684),
.B(n_1690),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1681),
.B(n_1643),
.Y(n_1696)
);

AOI221x1_ASAP7_75t_L g1697 ( 
.A1(n_1687),
.A2(n_1668),
.B1(n_1673),
.B2(n_1665),
.C(n_1663),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1681),
.A2(n_1670),
.B(n_1654),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1682),
.A2(n_1652),
.B1(n_1660),
.B2(n_1658),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1685),
.A2(n_1660),
.B1(n_1658),
.B2(n_1670),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1688),
.B(n_1644),
.C(n_1639),
.D(n_1658),
.Y(n_1701)
);

OAI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1683),
.A2(n_1655),
.B(n_1638),
.C(n_1639),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1694),
.A2(n_1683),
.B1(n_1689),
.B2(n_1644),
.C(n_1655),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1693),
.A2(n_1643),
.B1(n_1655),
.B2(n_1638),
.C(n_1648),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1698),
.A2(n_1638),
.B1(n_1650),
.B2(n_1648),
.C(n_1617),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1692),
.A2(n_1650),
.B(n_1624),
.C(n_1634),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1696),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1707),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1703),
.B(n_1699),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1704),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1705),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1707),
.Y(n_1713)
);

OAI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1710),
.A2(n_1702),
.B(n_1697),
.C(n_1695),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1715)
);

OAI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1709),
.A2(n_1700),
.B(n_1653),
.C(n_1622),
.Y(n_1716)
);

OAI211xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1712),
.A2(n_1631),
.B(n_1622),
.C(n_1606),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1718),
.B(n_1711),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_R g1720 ( 
.A(n_1715),
.B(n_1382),
.Y(n_1720)
);

NAND3x1_ASAP7_75t_L g1721 ( 
.A(n_1714),
.B(n_1625),
.C(n_1621),
.Y(n_1721)
);

NAND4xp75_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1716),
.C(n_1717),
.D(n_1606),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1722),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1723),
.B(n_1720),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1633),
.B1(n_1719),
.B2(n_1570),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1725),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1600),
.B1(n_1573),
.B2(n_1569),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1573),
.B(n_1600),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1728),
.B(n_1596),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1727),
.A2(n_1596),
.B1(n_1573),
.B2(n_1600),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1729),
.A2(n_1596),
.B(n_1627),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1730),
.A2(n_1627),
.B1(n_1571),
.B2(n_1618),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1731),
.Y(n_1733)
);

AOI22x1_ASAP7_75t_L g1734 ( 
.A1(n_1732),
.A2(n_1571),
.B1(n_1601),
.B2(n_1593),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1733),
.A2(n_1579),
.B1(n_1580),
.B2(n_1594),
.Y(n_1735)
);

OAI31xp33_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1734),
.A3(n_1594),
.B(n_1580),
.Y(n_1736)
);


endmodule