module real_aes_8349_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_1), .A2(n_157), .B(n_160), .C(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_2), .A2(n_186), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g486 ( .A(n_3), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_4), .B(n_216), .Y(n_215) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_5), .A2(n_186), .B(n_470), .Y(n_469) );
AND2x6_ASAP7_75t_L g157 ( .A(n_6), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g253 ( .A(n_7), .Y(n_253) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_8), .B(n_41), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_9), .A2(n_185), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_10), .B(n_169), .Y(n_242) );
INVx1_ASAP7_75t_L g474 ( .A(n_11), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_12), .B(n_210), .Y(n_509) );
INVx1_ASAP7_75t_L g149 ( .A(n_13), .Y(n_149) );
INVx1_ASAP7_75t_L g521 ( .A(n_14), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_15), .A2(n_78), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_15), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_16), .A2(n_194), .B(n_275), .C(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_17), .B(n_216), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_18), .B(n_452), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_19), .B(n_186), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_20), .B(n_200), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_21), .A2(n_210), .B(n_261), .C(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_22), .B(n_216), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_23), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_24), .A2(n_196), .B(n_277), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_25), .B(n_169), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_26), .Y(n_151) );
INVx1_ASAP7_75t_L g223 ( .A(n_27), .Y(n_223) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_28), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_29), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_30), .B(n_169), .Y(n_487) );
INVx1_ASAP7_75t_L g192 ( .A(n_31), .Y(n_192) );
INVx1_ASAP7_75t_L g464 ( .A(n_32), .Y(n_464) );
INVx2_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_34), .A2(n_128), .B1(n_131), .B2(n_725), .C1(n_726), .C2(n_728), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_35), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_36), .A2(n_210), .B(n_211), .C(n_213), .Y(n_209) );
INVxp67_ASAP7_75t_L g195 ( .A(n_37), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g208 ( .A(n_38), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_39), .A2(n_160), .B(n_222), .C(n_226), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_40), .A2(n_157), .B(n_160), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g463 ( .A(n_42), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_43), .A2(n_171), .B(n_251), .C(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_44), .B(n_169), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_45), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_46), .Y(n_188) );
INVx1_ASAP7_75t_L g259 ( .A(n_47), .Y(n_259) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_48), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_49), .A2(n_59), .B1(n_737), .B2(n_738), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_49), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_50), .B(n_186), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_51), .A2(n_160), .B1(n_263), .B2(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_52), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_53), .Y(n_483) );
CKINVDCx14_ASAP7_75t_R g249 ( .A(n_54), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_55), .A2(n_213), .B(n_251), .C(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_56), .Y(n_126) );
INVx1_ASAP7_75t_L g471 ( .A(n_57), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_58), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_59), .Y(n_738) );
INVx1_ASAP7_75t_L g158 ( .A(n_60), .Y(n_158) );
INVx1_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
INVx1_ASAP7_75t_SL g212 ( .A(n_62), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_63), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_64), .B(n_216), .Y(n_265) );
INVx1_ASAP7_75t_L g164 ( .A(n_65), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_SL g451 ( .A1(n_66), .A2(n_213), .B(n_452), .C(n_453), .Y(n_451) );
INVxp67_ASAP7_75t_L g454 ( .A(n_67), .Y(n_454) );
INVx1_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_69), .A2(n_186), .B(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_70), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_71), .A2(n_186), .B(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_72), .Y(n_467) );
INVx1_ASAP7_75t_L g527 ( .A(n_73), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_74), .A2(n_185), .B(n_187), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_75), .Y(n_220) );
INVx1_ASAP7_75t_L g273 ( .A(n_76), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_77), .A2(n_102), .B1(n_113), .B2(n_741), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_78), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_79), .A2(n_157), .B(n_160), .C(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_80), .A2(n_186), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g276 ( .A(n_81), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_82), .B(n_193), .Y(n_498) );
INVx2_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g241 ( .A(n_84), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_85), .B(n_452), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_86), .A2(n_157), .B(n_160), .C(n_485), .Y(n_484) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_87), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g122 ( .A(n_87), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g439 ( .A(n_87), .B(n_124), .Y(n_439) );
INVx2_ASAP7_75t_L g724 ( .A(n_87), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_88), .A2(n_160), .B(n_163), .C(n_173), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_89), .B(n_178), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_90), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_91), .A2(n_157), .B(n_160), .C(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_92), .Y(n_513) );
INVx1_ASAP7_75t_L g450 ( .A(n_93), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_94), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_95), .B(n_193), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_96), .B(n_144), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_97), .B(n_144), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g262 ( .A(n_99), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_100), .A2(n_186), .B(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_SL g741 ( .A(n_105), .Y(n_741) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g124 ( .A(n_109), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_127), .B1(n_731), .B2(n_733), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g732 ( .A(n_117), .Y(n_732) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_119), .A2(n_734), .B(n_739), .Y(n_733) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_126), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g740 ( .A(n_122), .Y(n_740) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_123), .B(n_724), .Y(n_730) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g723 ( .A(n_124), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_128), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_439), .B1(n_440), .B2(n_721), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_132), .A2(n_133), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_133), .A2(n_439), .B1(n_721), .B2(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_373), .Y(n_133) );
NAND5xp2_ASAP7_75t_L g134 ( .A(n_135), .B(n_302), .C(n_332), .D(n_353), .E(n_359), .Y(n_134) );
AOI221xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_232), .B1(n_266), .B2(n_268), .C(n_279), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_229), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_201), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_SL g353 ( .A1(n_140), .A2(n_217), .B(n_354), .C(n_357), .Y(n_353) );
AND2x2_ASAP7_75t_L g423 ( .A(n_140), .B(n_218), .Y(n_423) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_179), .Y(n_140) );
AND2x2_ASAP7_75t_L g281 ( .A(n_141), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g285 ( .A(n_141), .B(n_282), .Y(n_285) );
OR2x2_ASAP7_75t_L g311 ( .A(n_141), .B(n_218), .Y(n_311) );
AND2x2_ASAP7_75t_L g313 ( .A(n_141), .B(n_204), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_141), .B(n_203), .Y(n_331) );
INVx1_ASAP7_75t_L g364 ( .A(n_141), .Y(n_364) );
INVx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
BUFx2_ASAP7_75t_L g231 ( .A(n_142), .Y(n_231) );
AND2x2_ASAP7_75t_L g267 ( .A(n_142), .B(n_204), .Y(n_267) );
AND2x2_ASAP7_75t_L g420 ( .A(n_142), .B(n_218), .Y(n_420) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_150), .B(n_175), .Y(n_142) );
INVx3_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_143), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_143), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g500 ( .A(n_143), .B(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_144), .A2(n_448), .B(n_455), .Y(n_447) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_146), .B(n_147), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_159), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_152), .A2(n_178), .B(n_220), .C(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_239), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_152), .A2(n_174), .B1(n_461), .B2(n_465), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_152), .A2(n_483), .B(n_484), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_152), .A2(n_527), .B(n_528), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
AND2x4_ASAP7_75t_L g186 ( .A(n_153), .B(n_157), .Y(n_186) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx1_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g264 ( .A(n_155), .Y(n_264) );
INVx1_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx3_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx1_ASAP7_75t_L g452 ( .A(n_156), .Y(n_452) );
INVx4_ASAP7_75t_SL g174 ( .A(n_157), .Y(n_174) );
BUFx3_ASAP7_75t_L g226 ( .A(n_157), .Y(n_226) );
INVx5_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
AND2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
BUFx3_ASAP7_75t_L g172 ( .A(n_161), .Y(n_172) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_168), .C(n_170), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_165), .A2(n_170), .B(n_241), .C(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_166), .A2(n_167), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
INVx4_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx2_ASAP7_75t_L g251 ( .A(n_169), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_170), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_170), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g187 ( .A1(n_174), .A2(n_188), .B(n_189), .C(n_190), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_174), .A2(n_189), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_174), .A2(n_189), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_174), .A2(n_189), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_174), .A2(n_189), .B(n_273), .C(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_174), .A2(n_189), .B(n_450), .C(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_174), .A2(n_189), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_174), .A2(n_189), .B(n_518), .C(n_519), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g200 ( .A(n_177), .Y(n_200) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_177), .A2(n_505), .B(n_512), .Y(n_504) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g236 ( .A(n_178), .Y(n_236) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_178), .A2(n_247), .B(n_254), .Y(n_246) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_178), .A2(n_516), .B(n_522), .Y(n_515) );
AND2x2_ASAP7_75t_L g301 ( .A(n_179), .B(n_202), .Y(n_301) );
OR2x2_ASAP7_75t_L g305 ( .A(n_179), .B(n_218), .Y(n_305) );
AND2x2_ASAP7_75t_L g330 ( .A(n_179), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g377 ( .A(n_179), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_179), .B(n_339), .Y(n_425) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_198), .Y(n_179) );
INVx1_ASAP7_75t_L g283 ( .A(n_180), .Y(n_283) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_180), .A2(n_526), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_SL g494 ( .A1(n_181), .A2(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_182), .A2(n_460), .B(n_466), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_182), .B(n_467), .Y(n_466) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_182), .A2(n_482), .B(n_489), .Y(n_481) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_184), .A2(n_199), .B(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_191), .B(n_197), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_195), .B2(n_196), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_193), .A2(n_223), .B(n_224), .C(n_225), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_193), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
INVx5_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_194), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_194), .B(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_194), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_196), .B(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_196), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g225 ( .A(n_197), .Y(n_225) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OAI322xp33_ASAP7_75t_L g426 ( .A1(n_201), .A2(n_362), .A3(n_385), .B1(n_406), .B2(n_427), .C1(n_429), .C2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_202), .B(n_282), .Y(n_429) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g230 ( .A(n_203), .B(n_231), .Y(n_230) );
AND2x4_ASAP7_75t_L g298 ( .A(n_203), .B(n_218), .Y(n_298) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g339 ( .A(n_204), .B(n_218), .Y(n_339) );
AND2x2_ASAP7_75t_L g383 ( .A(n_204), .B(n_217), .Y(n_383) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_204) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_205), .A2(n_257), .B(n_265), .Y(n_256) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_205), .A2(n_271), .B(n_278), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_210), .B(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_214), .Y(n_510) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_216), .A2(n_469), .B(n_475), .Y(n_468) );
AND2x2_ASAP7_75t_L g266 ( .A(n_217), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g284 ( .A(n_217), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_217), .B(n_313), .Y(n_437) );
INVx3_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g229 ( .A(n_218), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_218), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g351 ( .A(n_218), .B(n_282), .Y(n_351) );
AND2x2_ASAP7_75t_L g378 ( .A(n_218), .B(n_313), .Y(n_378) );
OR2x2_ASAP7_75t_L g434 ( .A(n_218), .B(n_285), .Y(n_434) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
INVx1_ASAP7_75t_SL g320 ( .A(n_229), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_230), .B(n_351), .Y(n_352) );
AND2x2_ASAP7_75t_L g386 ( .A(n_230), .B(n_376), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_230), .B(n_309), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_230), .B(n_431), .Y(n_430) );
OAI31xp33_ASAP7_75t_L g404 ( .A1(n_232), .A2(n_266), .A3(n_405), .B(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_245), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_233), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g387 ( .A(n_233), .B(n_322), .Y(n_387) );
OR2x2_ASAP7_75t_L g394 ( .A(n_233), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g406 ( .A(n_233), .B(n_295), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g340 ( .A(n_234), .B(n_341), .Y(n_340) );
BUFx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g268 ( .A(n_235), .B(n_269), .Y(n_268) );
INVx4_ASAP7_75t_L g289 ( .A(n_235), .Y(n_289) );
AND2x2_ASAP7_75t_L g326 ( .A(n_235), .B(n_270), .Y(n_326) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_243), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_236), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_236), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_236), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g325 ( .A(n_245), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g395 ( .A(n_245), .Y(n_395) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_246), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_256), .Y(n_295) );
INVx2_ASAP7_75t_L g315 ( .A(n_246), .Y(n_315) );
AND2x2_ASAP7_75t_L g329 ( .A(n_246), .B(n_256), .Y(n_329) );
AND2x2_ASAP7_75t_L g336 ( .A(n_246), .B(n_292), .Y(n_336) );
BUFx3_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_246), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g291 ( .A(n_255), .Y(n_291) );
AND2x2_ASAP7_75t_L g299 ( .A(n_255), .B(n_289), .Y(n_299) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g269 ( .A(n_256), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_256), .Y(n_323) );
INVx2_ASAP7_75t_L g488 ( .A(n_263), .Y(n_488) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_SL g306 ( .A(n_267), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_267), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_267), .B(n_376), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_268), .B(n_346), .Y(n_399) );
INVx1_ASAP7_75t_SL g433 ( .A(n_268), .Y(n_433) );
INVx1_ASAP7_75t_SL g341 ( .A(n_269), .Y(n_341) );
INVx1_ASAP7_75t_SL g292 ( .A(n_270), .Y(n_292) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_270), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_289), .Y(n_314) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_289), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_270), .B(n_318), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B(n_286), .C(n_297), .Y(n_279) );
AOI31xp33_ASAP7_75t_L g396 ( .A1(n_280), .A2(n_397), .A3(n_398), .B(n_399), .Y(n_396) );
AND2x2_ASAP7_75t_L g369 ( .A(n_281), .B(n_298), .Y(n_369) );
BUFx3_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_282), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g345 ( .A(n_282), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_282), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g300 ( .A(n_285), .Y(n_300) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_285), .A2(n_410), .B1(n_413), .B2(n_414), .C1(n_415), .C2(n_416), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
INVx1_ASAP7_75t_L g415 ( .A(n_287), .Y(n_415) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_289), .B(n_292), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_289), .B(n_315), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_289), .B(n_290), .Y(n_385) );
INVx1_ASAP7_75t_L g436 ( .A(n_289), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_290), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g438 ( .A(n_290), .Y(n_438) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_292), .Y(n_361) );
AOI32xp33_ASAP7_75t_L g297 ( .A1(n_293), .A2(n_298), .A3(n_299), .B1(n_300), .B2(n_301), .Y(n_297) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_295), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_295), .Y(n_372) );
OR2x2_ASAP7_75t_L g413 ( .A(n_295), .B(n_314), .Y(n_413) );
INVx1_ASAP7_75t_L g349 ( .A(n_296), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_298), .B(n_309), .Y(n_334) );
INVx3_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
AOI322xp5_ASAP7_75t_L g359 ( .A1(n_298), .A2(n_343), .A3(n_360), .B1(n_362), .B2(n_365), .C1(n_369), .C2(n_370), .Y(n_359) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g412 ( .A(n_299), .Y(n_412) );
A2O1A1O1Ixp25_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_315), .D(n_316), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_303), .B(n_346), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_305), .A2(n_317), .B1(n_320), .B2(n_321), .C(n_324), .Y(n_316) );
INVx1_ASAP7_75t_SL g431 ( .A(n_305), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_314), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_309), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_311), .A2(n_395), .B1(n_402), .B2(n_403), .C(n_404), .Y(n_401) );
OAI222xp33_ASAP7_75t_L g432 ( .A1(n_312), .A2(n_433), .B1(n_434), .B2(n_435), .C1(n_437), .C2(n_438), .Y(n_432) );
AND2x2_ASAP7_75t_L g390 ( .A(n_313), .B(n_376), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_313), .A2(n_328), .B(n_375), .Y(n_402) );
INVx1_ASAP7_75t_L g416 ( .A(n_313), .Y(n_416) );
INVx2_ASAP7_75t_SL g319 ( .A(n_314), .Y(n_319) );
AND2x2_ASAP7_75t_L g322 ( .A(n_315), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_SL g356 ( .A(n_318), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_318), .B(n_328), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_319), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_319), .B(n_329), .Y(n_358) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_327), .B(n_330), .Y(n_324) );
INVx1_ASAP7_75t_SL g342 ( .A(n_326), .Y(n_342) );
AND2x2_ASAP7_75t_L g389 ( .A(n_326), .B(n_372), .Y(n_389) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g428 ( .A(n_328), .B(n_346), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_329), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g414 ( .A(n_330), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_344), .C(n_347), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B1(n_342), .B2(n_343), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_341), .A2(n_348), .B1(n_350), .B2(n_352), .Y(n_347) );
OR2x2_ASAP7_75t_L g418 ( .A(n_342), .B(n_346), .Y(n_418) );
OR2x2_ASAP7_75t_L g421 ( .A(n_342), .B(n_356), .Y(n_421) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_363), .A2(n_418), .B1(n_419), .B2(n_421), .C(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND3xp33_ASAP7_75t_SL g373 ( .A(n_374), .B(n_388), .C(n_400), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_379), .B1(n_381), .B2(n_384), .C1(n_386), .C2(n_387), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_376), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g398 ( .A(n_378), .Y(n_398) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_391), .B2(n_393), .C(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g403 ( .A(n_389), .Y(n_403) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
NOR5xp2_ASAP7_75t_L g400 ( .A(n_401), .B(n_409), .C(n_417), .D(n_426), .E(n_432), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g727 ( .A(n_440), .Y(n_727) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_441), .B(n_658), .Y(n_440) );
NOR4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_588), .C(n_619), .D(n_638), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_546), .C(n_561), .D(n_579), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_491), .B1(n_523), .B2(n_534), .C1(n_539), .C2(n_541), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_476), .Y(n_444) );
INVx1_ASAP7_75t_L g602 ( .A(n_445), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_456), .Y(n_445) );
AND2x2_ASAP7_75t_L g477 ( .A(n_446), .B(n_468), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_446), .B(n_480), .Y(n_631) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g538 ( .A(n_447), .B(n_458), .Y(n_538) );
AND2x2_ASAP7_75t_L g547 ( .A(n_447), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g573 ( .A(n_447), .Y(n_573) );
AND2x2_ASAP7_75t_L g594 ( .A(n_447), .B(n_458), .Y(n_594) );
BUFx2_ASAP7_75t_L g617 ( .A(n_447), .Y(n_617) );
AND2x2_ASAP7_75t_L g641 ( .A(n_447), .B(n_459), .Y(n_641) );
AND2x2_ASAP7_75t_L g705 ( .A(n_447), .B(n_468), .Y(n_705) );
AND2x2_ASAP7_75t_L g606 ( .A(n_456), .B(n_537), .Y(n_606) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_457), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
OR2x2_ASAP7_75t_L g566 ( .A(n_458), .B(n_481), .Y(n_566) );
AND2x2_ASAP7_75t_L g578 ( .A(n_458), .B(n_537), .Y(n_578) );
BUFx2_ASAP7_75t_L g710 ( .A(n_458), .Y(n_710) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g479 ( .A(n_459), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g560 ( .A(n_459), .B(n_481), .Y(n_560) );
AND2x2_ASAP7_75t_L g613 ( .A(n_459), .B(n_468), .Y(n_613) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_459), .Y(n_649) );
AND2x2_ASAP7_75t_L g536 ( .A(n_468), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_SL g548 ( .A(n_468), .Y(n_548) );
INVx2_ASAP7_75t_L g559 ( .A(n_468), .Y(n_559) );
BUFx2_ASAP7_75t_L g583 ( .A(n_468), .Y(n_583) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_468), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AOI332xp33_ASAP7_75t_L g561 ( .A1(n_477), .A2(n_562), .A3(n_566), .B1(n_567), .B2(n_571), .B3(n_574), .C1(n_575), .C2(n_577), .Y(n_561) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_477), .B(n_537), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_477), .B(n_551), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_SL g579 ( .A1(n_478), .A2(n_580), .B(n_583), .C(n_584), .Y(n_579) );
AND2x2_ASAP7_75t_L g718 ( .A(n_478), .B(n_559), .Y(n_718) );
INVx3_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g615 ( .A(n_479), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g620 ( .A(n_479), .B(n_617), .Y(n_620) );
INVx1_ASAP7_75t_L g551 ( .A(n_480), .Y(n_551) );
AND2x2_ASAP7_75t_L g654 ( .A(n_480), .B(n_613), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_480), .B(n_594), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_480), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_480), .B(n_572), .Y(n_680) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g537 ( .A(n_481), .Y(n_537) );
OAI31xp33_ASAP7_75t_L g719 ( .A1(n_491), .A2(n_640), .A3(n_647), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
AND2x2_ASAP7_75t_L g523 ( .A(n_492), .B(n_524), .Y(n_523) );
NAND2x1_ASAP7_75t_SL g542 ( .A(n_492), .B(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_492), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_492), .B(n_545), .Y(n_634) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_493), .A2(n_547), .B(n_549), .C(n_552), .Y(n_546) );
OR2x2_ASAP7_75t_L g563 ( .A(n_493), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g576 ( .A(n_493), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_493), .B(n_525), .Y(n_582) );
INVx2_ASAP7_75t_L g600 ( .A(n_493), .Y(n_600) );
AND2x2_ASAP7_75t_L g611 ( .A(n_493), .B(n_565), .Y(n_611) );
AND2x2_ASAP7_75t_L g643 ( .A(n_493), .B(n_601), .Y(n_643) );
AND2x2_ASAP7_75t_L g647 ( .A(n_493), .B(n_570), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_493), .B(n_502), .Y(n_652) );
AND2x2_ASAP7_75t_L g686 ( .A(n_493), .B(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_493), .B(n_589), .Y(n_720) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_502), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g628 ( .A(n_502), .Y(n_628) );
AND2x2_ASAP7_75t_L g690 ( .A(n_502), .B(n_611), .Y(n_690) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
OR2x2_ASAP7_75t_L g544 ( .A(n_503), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g554 ( .A(n_503), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_503), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g662 ( .A(n_503), .Y(n_662) );
AND2x2_ASAP7_75t_L g679 ( .A(n_503), .B(n_525), .Y(n_679) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g570 ( .A(n_504), .B(n_514), .Y(n_570) );
AND2x2_ASAP7_75t_L g599 ( .A(n_504), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g610 ( .A(n_504), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_504), .B(n_565), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g545 ( .A(n_515), .Y(n_545) );
AND2x2_ASAP7_75t_L g601 ( .A(n_515), .B(n_565), .Y(n_601) );
INVx1_ASAP7_75t_L g703 ( .A(n_523), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_524), .Y(n_707) );
INVx2_ASAP7_75t_L g565 ( .A(n_525), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_536), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_536), .B(n_641), .Y(n_699) );
OR2x2_ASAP7_75t_L g540 ( .A(n_537), .B(n_538), .Y(n_540) );
INVx1_ASAP7_75t_SL g592 ( .A(n_537), .Y(n_592) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_543), .A2(n_596), .B1(n_598), .B2(n_602), .C(n_603), .Y(n_595) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g623 ( .A(n_544), .B(n_587), .Y(n_623) );
INVx2_ASAP7_75t_L g555 ( .A(n_545), .Y(n_555) );
INVx1_ASAP7_75t_L g581 ( .A(n_545), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_545), .B(n_565), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_545), .B(n_568), .Y(n_675) );
INVx1_ASAP7_75t_L g683 ( .A(n_545), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_547), .B(n_551), .Y(n_597) );
AND2x4_ASAP7_75t_L g572 ( .A(n_548), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g685 ( .A(n_551), .B(n_641), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_554), .B(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_L g693 ( .A(n_555), .Y(n_693) );
INVxp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g593 ( .A(n_559), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g665 ( .A(n_559), .B(n_641), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_559), .B(n_578), .Y(n_671) );
AOI322xp5_ASAP7_75t_L g625 ( .A1(n_560), .A2(n_594), .A3(n_601), .B1(n_626), .B2(n_629), .C1(n_630), .C2(n_632), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_560), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g691 ( .A(n_563), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g637 ( .A(n_564), .Y(n_637) );
INVx2_ASAP7_75t_L g568 ( .A(n_565), .Y(n_568) );
INVx1_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_566), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g663 ( .A(n_568), .B(n_576), .Y(n_663) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g575 ( .A(n_570), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g618 ( .A(n_570), .B(n_611), .Y(n_618) );
AND2x2_ASAP7_75t_L g622 ( .A(n_570), .B(n_582), .Y(n_622) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_571), .A2(n_633), .B(n_635), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_571), .A2(n_703), .B1(n_704), .B2(n_706), .Y(n_702) );
INVx3_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g577 ( .A(n_572), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_572), .B(n_592), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_574), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g714 ( .A(n_581), .Y(n_714) );
INVx4_ASAP7_75t_L g587 ( .A(n_582), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_582), .B(n_609), .Y(n_657) );
INVx1_ASAP7_75t_SL g669 ( .A(n_583), .Y(n_669) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_587), .B(n_683), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_590), .B(n_595), .C(n_612), .Y(n_588) );
OAI221xp5_ASAP7_75t_SL g708 ( .A1(n_590), .A2(n_628), .B1(n_707), .B2(n_709), .C(n_711), .Y(n_708) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_592), .B(n_705), .Y(n_704) );
OAI31xp33_ASAP7_75t_L g684 ( .A1(n_593), .A2(n_670), .A3(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g624 ( .A(n_594), .Y(n_624) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g674 ( .A(n_599), .Y(n_674) );
AND2x2_ASAP7_75t_L g687 ( .A(n_601), .B(n_610), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_611), .B(n_714), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_618), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_621), .B1(n_623), .B2(n_624), .C(n_625), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_620), .A2(n_689), .B(n_691), .C(n_694), .Y(n_688) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_623), .B(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g650 ( .A(n_631), .Y(n_650) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g636 ( .A(n_634), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_634), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B(n_644), .C(n_653), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_642), .A2(n_652), .B1(n_716), .B2(n_717), .C(n_719), .Y(n_715) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_648), .B2(n_651), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_SL g716 ( .A(n_655), .Y(n_716) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_688), .C(n_708), .D(n_715), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_664), .B(n_666), .C(n_684), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B(n_672), .C(n_676), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g695 ( .A(n_673), .Y(n_695) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OR2x2_ASAP7_75t_L g706 ( .A(n_674), .B(n_707), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_700), .C(n_702), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_705), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule