module fake_jpeg_7192_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_15),
.B1(n_26),
.B2(n_13),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_26),
.Y(n_45)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_2),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_18),
.B(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_13),
.Y(n_66)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_15),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_26),
.B1(n_13),
.B2(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_27),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_54),
.B1(n_58),
.B2(n_30),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_29),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_34),
.Y(n_79)
);

OAI22x1_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_48),
.B1(n_30),
.B2(n_38),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_75),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_43),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_56),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_81),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_55),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_75),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_80),
.B1(n_52),
.B2(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_99),
.B1(n_103),
.B2(n_106),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_54),
.B1(n_58),
.B2(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_60),
.B1(n_63),
.B2(n_42),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_65),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_41),
.B1(n_19),
.B2(n_27),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_98),
.C(n_99),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_84),
.B(n_86),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_92),
.B1(n_93),
.B2(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_41),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_20),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_121),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_104),
.C(n_110),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_111),
.B(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_108),
.B1(n_118),
.B2(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_9),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_14),
.C(n_23),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_4),
.Y(n_134)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_124),
.B1(n_126),
.B2(n_10),
.C(n_3),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_128),
.C(n_4),
.Y(n_135)
);

AOI21x1_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_29),
.B(n_34),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_34),
.C(n_135),
.Y(n_139)
);


endmodule