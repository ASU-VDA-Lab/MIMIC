module fake_jpeg_11706_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_54),
.B(n_59),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_55),
.A2(n_38),
.B1(n_50),
.B2(n_20),
.Y(n_156)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_0),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_61),
.Y(n_134)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_65),
.B(n_74),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_49),
.C(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_72),
.Y(n_150)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_17),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g160 ( 
.A(n_76),
.Y(n_160)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_83),
.Y(n_138)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_3),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_29),
.B(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_96),
.Y(n_109)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_5),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_100),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_19),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_102),
.Y(n_151)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_111),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_106),
.B(n_87),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_44),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_27),
.B1(n_51),
.B2(n_36),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_121),
.B1(n_125),
.B2(n_47),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_27),
.B1(n_51),
.B2(n_36),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_120),
.A2(n_60),
.B1(n_75),
.B2(n_72),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_27),
.B1(n_51),
.B2(n_36),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_48),
.B1(n_46),
.B2(n_42),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_28),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_20),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_155),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_48),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_46),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_109),
.B1(n_104),
.B2(n_129),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_66),
.B(n_38),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_66),
.Y(n_175)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_134),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_162),
.B(n_180),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_114),
.B1(n_98),
.B2(n_93),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_163),
.A2(n_174),
.B1(n_182),
.B2(n_119),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_106),
.A2(n_64),
.B1(n_84),
.B2(n_92),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_195),
.Y(n_229)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_40),
.B(n_43),
.C(n_28),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_166),
.B(n_175),
.Y(n_225)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_170),
.A2(n_214),
.B(n_135),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_111),
.B(n_58),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_171),
.B(n_192),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_97),
.B1(n_95),
.B2(n_53),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_88),
.B1(n_79),
.B2(n_68),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_179),
.A2(n_200),
.B1(n_147),
.B2(n_123),
.Y(n_235)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_108),
.A2(n_69),
.B1(n_40),
.B2(n_43),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_184),
.B1(n_196),
.B2(n_198),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_141),
.A2(n_56),
.B1(n_62),
.B2(n_20),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_209),
.C(n_135),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_193),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_134),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_118),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_133),
.A2(n_50),
.B1(n_47),
.B2(n_90),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_126),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_203),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_133),
.A2(n_47),
.B1(n_78),
.B2(n_35),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_138),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_206),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_113),
.A2(n_35),
.B1(n_30),
.B2(n_80),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_138),
.A2(n_35),
.B1(n_30),
.B2(n_33),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_113),
.B(n_5),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_208),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_150),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_138),
.A2(n_33),
.B1(n_19),
.B2(n_9),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_107),
.B(n_5),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_117),
.B(n_5),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_130),
.B(n_142),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_140),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_33),
.B1(n_19),
.B2(n_10),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_142),
.CI(n_149),
.CON(n_219),
.SN(n_219)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_219),
.B(n_255),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_238),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_144),
.B1(n_159),
.B2(n_145),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_224),
.A2(n_228),
.B1(n_235),
.B2(n_243),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_144),
.B1(n_145),
.B2(n_135),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_231),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_180),
.A2(n_149),
.B1(n_147),
.B2(n_123),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_239),
.B1(n_248),
.B2(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_171),
.A2(n_122),
.B1(n_124),
.B2(n_136),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_124),
.B1(n_136),
.B2(n_131),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_131),
.C(n_128),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_211),
.Y(n_283)
);

BUFx24_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_128),
.B1(n_116),
.B2(n_126),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_116),
.B1(n_33),
.B2(n_19),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_249),
.A2(n_252),
.B1(n_194),
.B2(n_162),
.Y(n_297)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_185),
.A2(n_33),
.B1(n_19),
.B2(n_126),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_177),
.B(n_157),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_170),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_205),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_164),
.A2(n_157),
.B1(n_9),
.B2(n_10),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_173),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_177),
.B(n_172),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_264),
.A2(n_250),
.B(n_216),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_266),
.B(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_268),
.B(n_285),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_229),
.A2(n_164),
.B1(n_201),
.B2(n_208),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_269),
.A2(n_281),
.B1(n_297),
.B2(n_239),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_272),
.B(n_280),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_164),
.B1(n_201),
.B2(n_209),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_273),
.A2(n_274),
.B1(n_287),
.B2(n_254),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_201),
.B1(n_210),
.B2(n_178),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_236),
.C(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_289),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_195),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_235),
.A2(n_214),
.B1(n_166),
.B2(n_213),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_306),
.Y(n_335)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_241),
.B(n_168),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_167),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_291),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_232),
.B1(n_262),
.B2(n_238),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_247),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_221),
.B(n_231),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_300),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_191),
.Y(n_295)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_237),
.B1(n_246),
.B2(n_233),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_302),
.Y(n_333)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_257),
.B(n_203),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_176),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_219),
.B(n_161),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_304),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_230),
.B(n_190),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g305 ( 
.A1(n_223),
.A2(n_181),
.B(n_197),
.C(n_178),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g341 ( 
.A(n_305),
.B(n_246),
.C(n_233),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_219),
.B(n_165),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g319 ( 
.A(n_307),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_165),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_215),
.C(n_242),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_276),
.A2(n_227),
.B1(n_218),
.B2(n_259),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_270),
.B(n_306),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_312),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_270),
.A2(n_252),
.B(n_256),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_315),
.B(n_341),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_287),
.A2(n_240),
.B1(n_243),
.B2(n_248),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_320),
.B1(n_325),
.B2(n_337),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_293),
.A2(n_256),
.B(n_234),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_330),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_299),
.A2(n_307),
.B1(n_289),
.B2(n_282),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_309),
.B1(n_278),
.B2(n_319),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_266),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_332),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_217),
.B1(n_189),
.B2(n_187),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_234),
.B(n_237),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_331),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_300),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_275),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_271),
.A2(n_217),
.B1(n_189),
.B2(n_187),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_347),
.B(n_308),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_292),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_283),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_350),
.C(n_356),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_268),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_351),
.A2(n_353),
.B1(n_378),
.B2(n_337),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_280),
.B1(n_291),
.B2(n_273),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_352),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_338),
.A2(n_269),
.B1(n_265),
.B2(n_302),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_354),
.B(n_336),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_346),
.A2(n_265),
.B1(n_296),
.B2(n_286),
.Y(n_357)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_365),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_293),
.B1(n_281),
.B2(n_294),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_326),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_327),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_288),
.C(n_297),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_SL g405 ( 
.A(n_371),
.B(n_341),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_277),
.Y(n_372)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_277),
.B1(n_294),
.B2(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_295),
.B1(n_284),
.B2(n_215),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_344),
.B(n_311),
.Y(n_414)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_379),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_333),
.A2(n_222),
.B1(n_215),
.B2(n_226),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_382),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_342),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_372),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_397),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_389),
.C(n_391),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_390),
.A2(n_362),
.B1(n_361),
.B2(n_379),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_355),
.B(n_327),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_347),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_395),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_314),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_317),
.C(n_328),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_410),
.C(n_360),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_333),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_413),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_353),
.A2(n_325),
.B1(n_340),
.B2(n_334),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_403),
.A2(n_409),
.B1(n_381),
.B2(n_365),
.Y(n_415)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_407),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_405),
.B(n_413),
.Y(n_440)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_382),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_310),
.B(n_312),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_414),
.B(n_376),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_359),
.A2(n_340),
.B1(n_331),
.B2(n_321),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_368),
.B(n_329),
.C(n_323),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_360),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_380),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_344),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_415),
.A2(n_436),
.B1(n_398),
.B2(n_394),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_418),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_375),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_368),
.Y(n_419)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_409),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_402),
.Y(n_447)
);

AOI31xp33_ASAP7_75t_L g423 ( 
.A1(n_387),
.A2(n_359),
.A3(n_370),
.B(n_381),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_423),
.B(n_435),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_395),
.C(n_396),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_426),
.C(n_437),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_370),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_432),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_367),
.C(n_374),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_377),
.Y(n_427)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_383),
.Y(n_428)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_429),
.A2(n_434),
.B(n_439),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_430),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_363),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_363),
.B(n_311),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_406),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_362),
.C(n_361),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_345),
.B(n_322),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_SL g459 ( 
.A(n_440),
.B(n_322),
.C(n_307),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_394),
.C(n_385),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_447),
.Y(n_467)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_400),
.B(n_386),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_428),
.B(n_440),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_385),
.B1(n_412),
.B2(n_400),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_455),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_434),
.A2(n_403),
.B1(n_390),
.B2(n_412),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_453),
.B1(n_454),
.B2(n_433),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_426),
.A2(n_405),
.B1(n_386),
.B2(n_404),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_421),
.A2(n_432),
.B1(n_437),
.B2(n_417),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_319),
.B1(n_397),
.B2(n_345),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_319),
.B1(n_378),
.B2(n_323),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_460),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_459),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_419),
.A2(n_284),
.B1(n_222),
.B2(n_322),
.Y(n_460)
);

NOR3xp33_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_419),
.C(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_465),
.Y(n_481)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_463),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_439),
.B(n_427),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_464),
.A2(n_468),
.B(n_469),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_443),
.B(n_424),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_431),
.C(n_418),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_450),
.C(n_444),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_441),
.A2(n_433),
.B(n_431),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_470),
.A2(n_472),
.B1(n_476),
.B2(n_478),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_451),
.A2(n_222),
.B1(n_226),
.B2(n_261),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_442),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_461),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_453),
.A2(n_261),
.B1(n_12),
.B2(n_13),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_261),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_460),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_471),
.A2(n_452),
.B1(n_461),
.B2(n_442),
.Y(n_479)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_456),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_487),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_485),
.Y(n_496)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_456),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_477),
.C(n_454),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_490),
.B(n_493),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_464),
.A2(n_441),
.B(n_449),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_492),
.B(n_473),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_445),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_463),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_502),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_499),
.B(n_486),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_475),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g503 ( 
.A1(n_490),
.A2(n_468),
.B(n_476),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_505),
.B(n_488),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_472),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_491),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_483),
.A2(n_459),
.B(n_478),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_484),
.C(n_489),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_508),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_501),
.C(n_493),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_509),
.B(n_512),
.Y(n_518)
);

XOR2x2_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_483),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_510),
.A2(n_511),
.B(n_513),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_479),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_506),
.A2(n_497),
.B(n_505),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_516),
.B(n_517),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_500),
.C(n_494),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_518),
.Y(n_519)
);

AOI322xp5_ASAP7_75t_L g523 ( 
.A1(n_519),
.A2(n_491),
.A3(n_480),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_13),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_514),
.A2(n_503),
.B(n_487),
.Y(n_521)
);

OAI321xp33_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_12),
.A3(n_14),
.B1(n_16),
.B2(n_506),
.C(n_416),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_522),
.Y(n_525)
);


endmodule