module fake_netlist_5_174_n_2075 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2075);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2075;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1243;
wire n_1016;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_22),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_49),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_102),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_87),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_146),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_71),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_41),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_113),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_8),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_196),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_98),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_93),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_124),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_48),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_17),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_74),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_165),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_89),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_163),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_148),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_16),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_31),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_108),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_185),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_52),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_180),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_179),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_82),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_169),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_65),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_30),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_48),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_15),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_122),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_123),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_156),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_110),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_41),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_167),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_195),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_126),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_137),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_17),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_173),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_58),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_50),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_83),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_120),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_40),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_12),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_79),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_91),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_14),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_164),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_84),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_25),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_129),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_56),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_115),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_103),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_7),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_67),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_88),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_121),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_162),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_86),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_51),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_32),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_78),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_73),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_23),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_23),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_136),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_12),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_77),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_181),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_39),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_16),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_67),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_139),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_32),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_11),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_62),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_2),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_21),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_170),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_50),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_74),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_54),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_138),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_43),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_35),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_24),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_174),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_178),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_97),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_184),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_0),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_111),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_10),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_65),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_79),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_70),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_147),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_26),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_60),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_133),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_72),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_166),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_47),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_1),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_62),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_134),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_34),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_149),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_5),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_85),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_101),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_43),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_38),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_189),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_49),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_140),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_39),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_21),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_60),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_14),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_20),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_192),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_68),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_119),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_64),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_234),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_229),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_313),
.B(n_3),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_229),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_246),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_293),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_313),
.B(n_3),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_197),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_200),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_229),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_198),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_229),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_219),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_253),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_203),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_6),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_219),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_272),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_206),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_225),
.B(n_6),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_229),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_229),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_235),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_208),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_201),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_229),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_229),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_202),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_235),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_209),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_283),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_229),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_285),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_317),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_291),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_207),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_276),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_225),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_291),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_276),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_281),
.B(n_7),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_211),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_310),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_212),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_220),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_213),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_198),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_291),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_199),
.B(n_9),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_221),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_214),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_291),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_216),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_217),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_291),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_222),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_291),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_226),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_233),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_281),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_281),
.B(n_11),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_236),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_230),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_281),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_271),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_237),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_243),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_249),
.B(n_13),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_244),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_271),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_267),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_271),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_245),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_309),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_247),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_204),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_248),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_309),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_199),
.B(n_18),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_254),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_256),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_258),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_265),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_266),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_275),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_309),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_277),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_204),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_279),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_304),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_240),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_331),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_205),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_280),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_210),
.B(n_215),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_331),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_286),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_429),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_401),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_393),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_398),
.B(n_375),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_398),
.B(n_375),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_402),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_408),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_397),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_295),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_412),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_417),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_407),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_423),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_436),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_411),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_448),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_451),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_453),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_466),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_454),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_466),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_457),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_439),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g540 ( 
.A1(n_395),
.A2(n_278),
.B1(n_336),
.B2(n_351),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_403),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_461),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_267),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_424),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_331),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_405),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_470),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_414),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_472),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_415),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_455),
.B(n_459),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_426),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_400),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_419),
.B(n_267),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_475),
.B(n_478),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_413),
.B(n_391),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_425),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_425),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_479),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_526),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_480),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_566),
.A2(n_511),
.B1(n_561),
.B2(n_543),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_493),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_498),
.B(n_278),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_553),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_460),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_541),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_511),
.B(n_484),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_465),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_521),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_546),
.B(n_489),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_561),
.B(n_409),
.C(n_399),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_493),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_521),
.B(n_416),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_527),
.B(n_418),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_492),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_548),
.B(n_416),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_554),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_493),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_526),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_554),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_548),
.A2(n_422),
.B1(n_431),
.B2(n_437),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_558),
.B(n_465),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_526),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_531),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_556),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_503),
.Y(n_610)
);

INVxp67_ASAP7_75t_SL g611 ( 
.A(n_543),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_557),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_502),
.B(n_410),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_553),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_506),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_507),
.B(n_422),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_485),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_543),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_560),
.B(n_432),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_498),
.A2(n_351),
.B1(n_336),
.B2(n_224),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_549),
.B(n_431),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_563),
.B(n_432),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_531),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_549),
.B(n_435),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

AO22x2_ASAP7_75t_L g628 ( 
.A1(n_500),
.A2(n_224),
.B1(n_227),
.B2(n_205),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_564),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_565),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_503),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_531),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_508),
.B(n_438),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_502),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_531),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_531),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_568),
.B(n_432),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_568),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_497),
.A2(n_252),
.B1(n_380),
.B2(n_463),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_565),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_551),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_531),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_549),
.B(n_456),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_543),
.B(n_432),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_514),
.B(n_440),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_551),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_516),
.B(n_486),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_513),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_510),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_456),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_531),
.B(n_296),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_494),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_535),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_513),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_504),
.B(n_467),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_496),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_538),
.B(n_486),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_515),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_496),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_540),
.B(n_467),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_540),
.B(n_469),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_515),
.Y(n_669)
);

OA22x2_ASAP7_75t_L g670 ( 
.A1(n_540),
.A2(n_273),
.B1(n_274),
.B2(n_227),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_562),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_499),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_538),
.B(n_474),
.C(n_443),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_515),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_500),
.A2(n_449),
.B1(n_462),
.B2(n_445),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_469),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_499),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_539),
.A2(n_468),
.B1(n_476),
.B2(n_464),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_535),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_504),
.B(n_473),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_535),
.B(n_303),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_501),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_SL g686 ( 
.A(n_539),
.B(n_232),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_544),
.A2(n_210),
.B1(n_323),
.B2(n_312),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_535),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_504),
.B(n_473),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_523),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_523),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_505),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_562),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_530),
.B(n_481),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_532),
.B(n_481),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_509),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_517),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_509),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_520),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_535),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_532),
.B(n_491),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_535),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_518),
.B(n_477),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_547),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_547),
.B(n_301),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_572),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_547),
.B(n_303),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_519),
.B(n_482),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_547),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_404),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_570),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_570),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_524),
.B(n_375),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_547),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_528),
.A2(n_427),
.B1(n_428),
.B2(n_242),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_572),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_547),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_533),
.B(n_215),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_550),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_550),
.B(n_318),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_550),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_605),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_575),
.B(n_529),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_576),
.B(n_534),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_611),
.B(n_619),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_580),
.B(n_585),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_586),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_626),
.B(n_550),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_622),
.A2(n_512),
.B1(n_542),
.B2(n_555),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_622),
.A2(n_571),
.B1(n_537),
.B2(n_552),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_662),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_626),
.B(n_550),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_578),
.B(n_628),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_573),
.A2(n_332),
.B(n_364),
.C(n_223),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_586),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_626),
.A2(n_562),
.B1(n_332),
.B2(n_218),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_683),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_582),
.B(n_595),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_683),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_647),
.A2(n_562),
.B1(n_223),
.B2(n_228),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_658),
.A2(n_569),
.B(n_550),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_580),
.B(n_441),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_683),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_667),
.B(n_218),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_647),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_689),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_647),
.A2(n_562),
.B1(n_231),
.B2(n_238),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_585),
.B(n_471),
.Y(n_754)
);

NOR2x1p5_ASAP7_75t_L g755 ( 
.A(n_630),
.B(n_250),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_604),
.B(n_483),
.Y(n_756)
);

BUFx8_ASAP7_75t_L g757 ( 
.A(n_634),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_606),
.B(n_550),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_630),
.B(n_321),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_689),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_606),
.B(n_569),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_579),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_597),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_689),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_656),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_578),
.A2(n_312),
.B1(n_290),
.B2(n_289),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_573),
.B(n_569),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_589),
.B(n_512),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_604),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_594),
.B(n_522),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_676),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_584),
.B(n_569),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_667),
.A2(n_562),
.B1(n_228),
.B2(n_335),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_642),
.B(n_324),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_634),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_584),
.B(n_569),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_693),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_602),
.B(n_569),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_545),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_590),
.B(n_559),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_656),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_656),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_708),
.A2(n_569),
.B(n_536),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_602),
.B(n_570),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_668),
.A2(n_562),
.B1(n_231),
.B2(n_339),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_609),
.B(n_570),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_724),
.A2(n_536),
.B(n_533),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_609),
.B(n_570),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_612),
.B(n_617),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_664),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_612),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_693),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_631),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_617),
.B(n_570),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_625),
.B(n_570),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_625),
.B(n_562),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_583),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_578),
.A2(n_345),
.B1(n_349),
.B2(n_353),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_627),
.B(n_533),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_627),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_642),
.B(n_648),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_629),
.B(n_533),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_668),
.A2(n_289),
.B1(n_377),
.B2(n_364),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_655),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_655),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_581),
.B(n_536),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_598),
.B(n_638),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_631),
.B(n_359),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_613),
.B(n_292),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_699),
.B(n_536),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_697),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_620),
.B(n_367),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_700),
.B(n_567),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_713),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_705),
.B(n_567),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_613),
.B(n_463),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_657),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_623),
.B(n_369),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_657),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_697),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_637),
.B(n_373),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_698),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_659),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_659),
.B(n_567),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_673),
.B(n_488),
.C(n_257),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_698),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_618),
.B(n_378),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_578),
.A2(n_381),
.B1(n_383),
.B2(n_260),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_663),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_663),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_666),
.B(n_567),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_666),
.B(n_238),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_628),
.A2(n_261),
.B1(n_260),
.B2(n_259),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_722),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_672),
.B(n_251),
.Y(n_836)
);

INVxp33_ASAP7_75t_SL g837 ( 
.A(n_641),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_687),
.B(n_251),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_678),
.B(n_259),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_628),
.A2(n_261),
.B1(n_290),
.B2(n_308),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_675),
.B(n_308),
.Y(n_842)
);

AND2x6_ASAP7_75t_SL g843 ( 
.A(n_616),
.B(n_273),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_628),
.A2(n_339),
.B1(n_335),
.B2(n_354),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_722),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_605),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_621),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_678),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_621),
.A2(n_323),
.B1(n_355),
.B2(n_356),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_682),
.B(n_685),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_722),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_593),
.B(n_319),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_682),
.B(n_685),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_692),
.B(n_358),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_692),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_709),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_676),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_664),
.B(n_255),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_645),
.A2(n_358),
.B(n_377),
.C(n_239),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_645),
.A2(n_239),
.B(n_362),
.C(n_387),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_709),
.Y(n_861)
);

BUFx5_ASAP7_75t_L g862 ( 
.A(n_684),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_614),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_603),
.B(n_262),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_725),
.B(n_491),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_725),
.B(n_263),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_713),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_712),
.B(n_264),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_719),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_688),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_716),
.B(n_268),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_713),
.B(n_269),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_719),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_721),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_712),
.B(n_270),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_723),
.B(n_282),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_677),
.B(n_274),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_577),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_605),
.B(n_686),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_688),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_577),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_621),
.A2(n_392),
.B1(n_390),
.B2(n_284),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_294),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_686),
.B(n_299),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_621),
.A2(n_240),
.B1(n_241),
.B2(n_388),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_717),
.B(n_300),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_591),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_717),
.B(n_302),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_679),
.B(n_718),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_592),
.B(n_305),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_713),
.B(n_677),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_670),
.A2(n_362),
.B1(n_387),
.B2(n_287),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_651),
.B(n_306),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_592),
.B(n_307),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_670),
.A2(n_342),
.B1(n_386),
.B2(n_385),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_633),
.B(n_287),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_591),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_804),
.B(n_649),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_863),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_736),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_751),
.B(n_592),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_751),
.B(n_600),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_729),
.B(n_600),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_824),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_762),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_863),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_727),
.B(n_650),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_765),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_730),
.B(n_704),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_732),
.A2(n_654),
.B(n_650),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_797),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_852),
.A2(n_333),
.B1(n_334),
.B2(n_315),
.C(n_298),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_775),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_771),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_738),
.A2(n_654),
.B(n_707),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_711),
.C(n_314),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_726),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_765),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_804),
.B(n_311),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_730),
.B(n_791),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_824),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_741),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_757),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_793),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_737),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_791),
.B(n_639),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_800),
.B(n_643),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_737),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_743),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_800),
.B(n_805),
.Y(n_932)
);

CKINVDCx11_ASAP7_75t_R g933 ( 
.A(n_726),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_757),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_763),
.B(n_790),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_830),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_805),
.B(n_644),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_818),
.B(n_600),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_743),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_744),
.B(n_670),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_897),
.B(n_608),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_818),
.B(n_608),
.Y(n_942)
);

AOI22x1_ASAP7_75t_L g943 ( 
.A1(n_830),
.A2(n_660),
.B1(n_706),
.B2(n_608),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_781),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_745),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_752),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_SL g947 ( 
.A(n_806),
.B(n_322),
.C(n_320),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_820),
.B(n_632),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_820),
.A2(n_601),
.B(n_599),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_839),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_793),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_797),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_831),
.B(n_632),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_781),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_752),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_771),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_782),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_782),
.B(n_632),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_892),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_739),
.B(n_695),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_846),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_745),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_741),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_846),
.Y(n_964)
);

NOR2x1_ASAP7_75t_L g965 ( 
.A(n_755),
.B(n_646),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_897),
.B(n_646),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_839),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_831),
.B(n_646),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_848),
.B(n_660),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_760),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_748),
.B(n_754),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_760),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_SL g973 ( 
.A(n_871),
.B(n_326),
.C(n_325),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_848),
.B(n_660),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_777),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_768),
.B(n_706),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_777),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_771),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_806),
.B(n_240),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_834),
.B(n_706),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_757),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_748),
.B(n_695),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_857),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_792),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_764),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_823),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_857),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_764),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_735),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_810),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_735),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_750),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_750),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_823),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_827),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_745),
.B(n_596),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_750),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_835),
.B(n_845),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_792),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_812),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_857),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_812),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_858),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_870),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_749),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_749),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_870),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_821),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_842),
.A2(n_684),
.B1(n_710),
.B2(n_691),
.Y(n_1009)
);

BUFx10_ASAP7_75t_L g1010 ( 
.A(n_770),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_841),
.B(n_583),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_870),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_837),
.A2(n_327),
.B1(n_328),
.B2(n_384),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_835),
.B(n_596),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_815),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_821),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_728),
.A2(n_715),
.B1(n_714),
.B2(n_696),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_815),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_855),
.B(n_696),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_855),
.B(n_702),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_892),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_SL g1023 ( 
.A(n_827),
.B(n_348),
.C(n_329),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_856),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_869),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_842),
.B(n_801),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_754),
.B(n_702),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_869),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_881),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_808),
.A2(n_715),
.B1(n_714),
.B2(n_574),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_734),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_845),
.B(n_596),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_873),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_769),
.B(n_574),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_731),
.B(n_574),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_731),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_837),
.A2(n_780),
.B1(n_779),
.B2(n_872),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_844),
.A2(n_684),
.B1(n_710),
.B2(n_599),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_873),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_856),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_851),
.B(n_596),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_L g1042 ( 
.A(n_867),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_808),
.B(n_588),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_733),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_881),
.Y(n_1045)
);

AND2x6_ASAP7_75t_L g1046 ( 
.A(n_756),
.B(n_583),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_847),
.A2(n_374),
.B(n_297),
.C(n_298),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_861),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_877),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_756),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_739),
.Y(n_1051)
);

BUFx8_ASAP7_75t_L g1052 ( 
.A(n_867),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_851),
.B(n_596),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_789),
.B(n_583),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_878),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_739),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_SL g1057 ( 
.A(n_739),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_808),
.B(n_671),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_849),
.A2(n_684),
.B1(n_710),
.B2(n_615),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_843),
.B(n_330),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_758),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_796),
.B(n_671),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_861),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_877),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_886),
.A2(n_684),
.B1(n_710),
.B2(n_615),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_878),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_874),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_874),
.Y(n_1068)
);

AO22x1_ASAP7_75t_L g1069 ( 
.A1(n_766),
.A2(n_347),
.B1(n_368),
.B2(n_376),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_877),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_817),
.Y(n_1071)
);

OR2x4_ASAP7_75t_L g1072 ( 
.A(n_817),
.B(n_288),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_761),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_891),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_850),
.B(n_583),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_880),
.B(n_588),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_862),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_798),
.Y(n_1078)
);

CKINVDCx6p67_ASAP7_75t_R g1079 ( 
.A(n_759),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_853),
.B(n_588),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_879),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_838),
.B(n_680),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_866),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_868),
.B(n_680),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_879),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_807),
.Y(n_1086)
);

AOI211xp5_ASAP7_75t_L g1087 ( 
.A1(n_826),
.A2(n_379),
.B(n_346),
.C(n_344),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_882),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_882),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_862),
.B(n_671),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_862),
.B(n_671),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_L g1092 ( 
.A(n_1003),
.B(n_774),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_913),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_962),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_943),
.A2(n_787),
.B(n_783),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_938),
.A2(n_747),
.B(n_767),
.Y(n_1096)
);

BUFx4f_ASAP7_75t_SL g1097 ( 
.A(n_925),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_913),
.Y(n_1098)
);

OA22x2_ASAP7_75t_L g1099 ( 
.A1(n_1044),
.A2(n_990),
.B1(n_883),
.B2(n_1013),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_982),
.B(n_803),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1027),
.B(n_833),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_942),
.A2(n_776),
.B(n_772),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_948),
.A2(n_778),
.B(n_784),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1026),
.B(n_918),
.C(n_1087),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_911),
.B(n_864),
.Y(n_1105)
);

NOR2xp67_ASAP7_75t_L g1106 ( 
.A(n_973),
.B(n_829),
.Y(n_1106)
);

AND3x4_ASAP7_75t_L g1107 ( 
.A(n_947),
.B(n_894),
.C(n_885),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_922),
.A2(n_854),
.B1(n_836),
.B2(n_840),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_913),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_953),
.A2(n_788),
.B(n_786),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_968),
.A2(n_795),
.B(n_794),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_913),
.A2(n_1077),
.B(n_917),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_913),
.A2(n_802),
.B(n_799),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_969),
.A2(n_898),
.B(n_888),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_906),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1077),
.A2(n_832),
.B(n_825),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_906),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_901),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_971),
.B(n_828),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_974),
.A2(n_898),
.B(n_888),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_SL g1121 ( 
.A(n_900),
.B(n_895),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_905),
.A2(n_740),
.B(n_876),
.C(n_889),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1077),
.A2(n_814),
.B(n_811),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_912),
.A2(n_816),
.B(n_887),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1061),
.A2(n_909),
.B(n_1054),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1007),
.A2(n_865),
.B(n_884),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_924),
.B(n_809),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1070),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_935),
.B(n_875),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1075),
.A2(n_680),
.B(n_742),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_923),
.Y(n_1131)
);

OA22x2_ASAP7_75t_L g1132 ( 
.A1(n_1044),
.A2(n_896),
.B1(n_288),
.B2(n_297),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1007),
.A2(n_669),
.B(n_601),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_1026),
.A2(n_813),
.B(n_819),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1083),
.B(n_893),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_959),
.A2(n_1022),
.B1(n_1050),
.B2(n_993),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_976),
.B(n_822),
.Y(n_1137)
);

OA22x2_ASAP7_75t_L g1138 ( 
.A1(n_1078),
.A2(n_361),
.B1(n_388),
.B2(n_374),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1007),
.A2(n_665),
.B(n_640),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_908),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1012),
.A2(n_665),
.B(n_640),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1071),
.B(n_773),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_923),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_976),
.B(n_785),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_932),
.A2(n_960),
.B1(n_1021),
.B2(n_1020),
.Y(n_1145)
);

INVx6_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_936),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1074),
.B(n_941),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_941),
.A2(n_859),
.A3(n_860),
.B(n_661),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1001),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_933),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_966),
.B(n_746),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_966),
.B(n_753),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1070),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_940),
.A2(n_652),
.B(n_653),
.Y(n_1156)
);

AOI31xp67_ASAP7_75t_L g1157 ( 
.A1(n_905),
.A2(n_674),
.A3(n_652),
.B(n_681),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_960),
.A2(n_587),
.B1(n_720),
.B2(n_607),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_940),
.B(n_653),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1004),
.A2(n_607),
.B(n_720),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_992),
.B(n_661),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_907),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1037),
.A2(n_340),
.B(n_338),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_997),
.B(n_1049),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_1046),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1064),
.B(n_669),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_914),
.A2(n_350),
.B(n_372),
.C(n_371),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1047),
.A2(n_350),
.B(n_372),
.C(n_371),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_674),
.B(n_681),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_962),
.Y(n_1170)
);

CKINVDCx11_ASAP7_75t_R g1171 ( 
.A(n_933),
.Y(n_1171)
);

AND3x4_ASAP7_75t_L g1172 ( 
.A(n_1023),
.B(n_240),
.C(n_241),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_900),
.B(n_587),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1004),
.A2(n_587),
.B(n_720),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_960),
.A2(n_334),
.B1(n_315),
.B2(n_366),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1078),
.A2(n_357),
.B1(n_365),
.B2(n_337),
.C(n_341),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1062),
.A2(n_1018),
.B(n_1080),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1012),
.A2(n_690),
.B(n_691),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_903),
.A2(n_904),
.B(n_1063),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_998),
.A2(n_929),
.B(n_928),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_935),
.B(n_241),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1047),
.A2(n_366),
.B(n_333),
.C(n_363),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1062),
.A2(n_690),
.B(n_710),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_950),
.A2(n_363),
.A3(n_361),
.B(n_862),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_903),
.A2(n_862),
.B(n_720),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_967),
.A2(n_862),
.A3(n_710),
.B(n_684),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_904),
.A2(n_862),
.B(n_720),
.Y(n_1187)
);

INVx6_ASAP7_75t_SL g1188 ( 
.A(n_960),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_962),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1004),
.A2(n_624),
.B(n_703),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_924),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_956),
.B(n_862),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1070),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1029),
.A2(n_703),
.B(n_701),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_945),
.A2(n_1029),
.B1(n_956),
.B2(n_1045),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1010),
.B(n_241),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1080),
.A2(n_996),
.B(n_967),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_902),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_925),
.B(n_587),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_945),
.A2(n_703),
.B1(n_701),
.B2(n_587),
.Y(n_1200)
);

AOI22x1_ASAP7_75t_L g1201 ( 
.A1(n_975),
.A2(n_703),
.B1(n_701),
.B2(n_636),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_900),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_934),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_915),
.B(n_343),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1029),
.A2(n_701),
.B(n_607),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_952),
.B(n_607),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_937),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_956),
.B(n_607),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_956),
.A2(n_624),
.B(n_635),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1001),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_636),
.B(n_635),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_958),
.A2(n_636),
.B(n_635),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_SL g1213 ( 
.A1(n_952),
.A2(n_81),
.B(n_188),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_952),
.B(n_636),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_927),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_930),
.B(n_624),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_SL g1217 ( 
.A(n_951),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_956),
.A2(n_624),
.B(n_635),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1045),
.B(n_624),
.Y(n_1219)
);

NOR4xp25_ASAP7_75t_L g1220 ( 
.A(n_931),
.B(n_370),
.C(n_360),
.D(n_352),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_958),
.A2(n_636),
.B(n_635),
.Y(n_1221)
);

OAI22x1_ASAP7_75t_L g1222 ( 
.A1(n_1031),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1045),
.A2(n_694),
.B(n_671),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1001),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_975),
.A2(n_694),
.B(n_176),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_977),
.A2(n_694),
.B(n_175),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_926),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1045),
.B(n_694),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_977),
.A2(n_694),
.B(n_172),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_984),
.A2(n_160),
.B(n_158),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1043),
.A2(n_152),
.B(n_151),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_939),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_L g1233 ( 
.A(n_1079),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_986),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1031),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_984),
.A2(n_150),
.B(n_144),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_999),
.A2(n_143),
.B(n_135),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_999),
.A2(n_127),
.B(n_125),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_946),
.B(n_29),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_955),
.B(n_33),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_994),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1045),
.A2(n_117),
.B(n_116),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1024),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1024),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1080),
.A2(n_106),
.B(n_105),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1015),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1040),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1025),
.A2(n_1028),
.B(n_1039),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1000),
.A2(n_104),
.B(n_99),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1000),
.A2(n_95),
.B(n_94),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1051),
.B(n_90),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_970),
.B(n_35),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_916),
.A2(n_978),
.B(n_983),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_972),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1002),
.A2(n_36),
.B(n_37),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1115),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1198),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1162),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1115),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1129),
.A2(n_1057),
.B1(n_1070),
.B2(n_1034),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1212),
.A2(n_1221),
.B(n_1120),
.Y(n_1262)
);

OAI211xp5_ASAP7_75t_L g1263 ( 
.A1(n_1176),
.A2(n_1060),
.B(n_921),
.C(n_899),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1171),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1114),
.A2(n_998),
.B(n_1002),
.Y(n_1265)
);

INVxp67_ASAP7_75t_SL g1266 ( 
.A(n_1162),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1095),
.A2(n_1017),
.B(n_1008),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1163),
.A2(n_979),
.B1(n_1069),
.B2(n_1060),
.C(n_921),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1225),
.A2(n_1229),
.B(n_1226),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1112),
.A2(n_949),
.B(n_1030),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1101),
.B(n_985),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1099),
.A2(n_1057),
.B1(n_1079),
.B2(n_1010),
.Y(n_1272)
);

AOI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1112),
.A2(n_1084),
.B(n_1076),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1125),
.A2(n_1035),
.B(n_1084),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1211),
.A2(n_1040),
.B(n_1067),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1129),
.B(n_988),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1125),
.A2(n_1035),
.B(n_1084),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1099),
.A2(n_1010),
.B1(n_899),
.B2(n_986),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1096),
.A2(n_1048),
.B(n_1085),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1215),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1232),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1254),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1126),
.A2(n_1048),
.B(n_1085),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1133),
.A2(n_1067),
.B(n_1081),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1139),
.A2(n_1081),
.B(n_1055),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1117),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1148),
.B(n_1019),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1124),
.A2(n_1084),
.B(n_987),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1141),
.A2(n_1033),
.B(n_1066),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1124),
.A2(n_1122),
.B(n_1103),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1143),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1147),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1104),
.A2(n_1057),
.B1(n_1034),
.B2(n_1036),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1100),
.B(n_1034),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1144),
.A2(n_991),
.B(n_1006),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1105),
.B(n_995),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1171),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1181),
.A2(n_995),
.B1(n_961),
.B2(n_964),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1169),
.A2(n_1088),
.B(n_1068),
.Y(n_1300)
);

AOI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_1076),
.B(n_1053),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1137),
.A2(n_1005),
.B(n_989),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1136),
.A2(n_961),
.B1(n_964),
.B2(n_1072),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1105),
.A2(n_1043),
.B1(n_1042),
.B2(n_945),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1234),
.A2(n_1072),
.B1(n_981),
.B2(n_963),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1178),
.A2(n_1041),
.B(n_1014),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1185),
.A2(n_1041),
.B(n_1014),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1142),
.A2(n_919),
.B1(n_1042),
.B2(n_944),
.Y(n_1308)
);

AOI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1145),
.A2(n_1076),
.B(n_1053),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1195),
.A2(n_1076),
.B(n_965),
.Y(n_1310)
);

AO21x1_ASAP7_75t_L g1311 ( 
.A1(n_1108),
.A2(n_996),
.B(n_1082),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1152),
.A2(n_1009),
.B(n_1065),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1155),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1151),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1243),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1244),
.Y(n_1317)
);

BUFx2_ASAP7_75t_R g1318 ( 
.A(n_1118),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1187),
.A2(n_1091),
.B(n_1090),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1106),
.A2(n_1086),
.B(n_1043),
.C(n_1082),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1167),
.A2(n_919),
.B1(n_1086),
.B2(n_1082),
.C(n_1073),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1118),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1244),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1097),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1135),
.B(n_1073),
.Y(n_1325)
);

AOI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1119),
.A2(n_910),
.B(n_920),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1153),
.A2(n_1058),
.B(n_980),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1247),
.Y(n_1328)
);

INVx6_ASAP7_75t_L g1329 ( 
.A(n_1128),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_1091),
.B(n_1090),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1093),
.A2(n_1058),
.B(n_1073),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1247),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1165),
.B(n_1093),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_SL g1334 ( 
.A1(n_1168),
.A2(n_1011),
.B(n_980),
.C(n_1046),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1165),
.A2(n_910),
.B1(n_920),
.B2(n_944),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1102),
.A2(n_1032),
.B(n_1038),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1165),
.A2(n_910),
.B1(n_920),
.B2(n_944),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1110),
.A2(n_1032),
.B(n_1059),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1111),
.A2(n_1201),
.B(n_1230),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1203),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1248),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1098),
.A2(n_1073),
.B(n_1016),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1092),
.B(n_910),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1159),
.B(n_949),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1097),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1246),
.B(n_920),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1132),
.A2(n_980),
.B1(n_954),
.B2(n_957),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_SL g1348 ( 
.A1(n_1134),
.A2(n_1177),
.B(n_1121),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1167),
.A2(n_957),
.B1(n_954),
.B2(n_944),
.C(n_1089),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1113),
.A2(n_1046),
.B(n_1011),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1132),
.A2(n_980),
.B1(n_954),
.B2(n_957),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1236),
.A2(n_1046),
.B(n_980),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1140),
.Y(n_1353)
);

BUFx8_ASAP7_75t_L g1354 ( 
.A(n_1217),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1184),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1184),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1113),
.A2(n_1046),
.B(n_1011),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1184),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1237),
.A2(n_1011),
.B(n_1089),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1241),
.B(n_957),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1107),
.A2(n_954),
.B1(n_1011),
.B2(n_1052),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1227),
.B(n_1052),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1238),
.A2(n_1089),
.B(n_1016),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1204),
.B(n_1089),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1168),
.A2(n_1016),
.A3(n_1001),
.B(n_42),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1098),
.A2(n_1016),
.B(n_38),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1249),
.A2(n_37),
.B(n_42),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1191),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1175),
.B(n_44),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1175),
.B(n_44),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1127),
.B(n_80),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1122),
.A2(n_1255),
.B(n_1156),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1250),
.A2(n_1116),
.B(n_1123),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1197),
.A2(n_45),
.B(n_46),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_SL g1375 ( 
.A(n_1233),
.B(n_45),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1213),
.A2(n_46),
.B(n_52),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1165),
.B(n_53),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1109),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1116),
.A2(n_54),
.B(n_55),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1123),
.A2(n_55),
.B(n_56),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1130),
.A2(n_57),
.B(n_58),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1220),
.B(n_59),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1127),
.B(n_59),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1233),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1239),
.B(n_61),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1196),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1146),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1160),
.A2(n_61),
.B(n_63),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1240),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1204),
.B(n_66),
.C(n_68),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1217),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1160),
.A2(n_66),
.B(n_70),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1164),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1108),
.B(n_72),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1130),
.A2(n_1253),
.B(n_1183),
.Y(n_1395)
);

BUFx8_ASAP7_75t_L g1396 ( 
.A(n_1150),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1245),
.A2(n_1242),
.B(n_1252),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1161),
.B(n_80),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1253),
.A2(n_73),
.B(n_75),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1166),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1150),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1146),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1182),
.A2(n_75),
.A3(n_76),
.B(n_77),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1184),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1174),
.A2(n_1190),
.B(n_1205),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1150),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1109),
.B(n_1128),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1216),
.B(n_1149),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1146),
.A2(n_1138),
.B1(n_1251),
.B2(n_1193),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1182),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1150),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1210),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1138),
.A2(n_1251),
.B1(n_1193),
.B2(n_1154),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1251),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1245),
.A2(n_1190),
.B(n_1174),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1194),
.A2(n_1205),
.B(n_1209),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1094),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1242),
.B(n_1231),
.C(n_1199),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1107),
.B(n_1154),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1210),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1202),
.B(n_1094),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1208),
.A2(n_1219),
.B(n_1192),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1172),
.B(n_1188),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1369),
.A2(n_1235),
.B1(n_1222),
.B2(n_1172),
.Y(n_1424)
);

AOI222xp33_ASAP7_75t_L g1425 ( 
.A1(n_1369),
.A2(n_1158),
.B1(n_1219),
.B2(n_1208),
.C1(n_1192),
.C2(n_1202),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1370),
.A2(n_1188),
.B1(n_1199),
.B2(n_1170),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1271),
.B(n_1224),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1297),
.B(n_1224),
.Y(n_1428)
);

NAND2x1_ASAP7_75t_L g1429 ( 
.A(n_1378),
.B(n_1189),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1370),
.A2(n_1199),
.B1(n_1170),
.B2(n_1189),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1368),
.Y(n_1431)
);

AOI21xp33_ASAP7_75t_L g1432 ( 
.A1(n_1394),
.A2(n_1200),
.B(n_1224),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1299),
.A2(n_1173),
.B1(n_1214),
.B2(n_1206),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1375),
.A2(n_1210),
.B1(n_1224),
.B2(n_1173),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1399),
.A2(n_1194),
.B(n_1209),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1318),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1272),
.A2(n_1386),
.B1(n_1278),
.B2(n_1364),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1368),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1268),
.A2(n_1206),
.B1(n_1214),
.B2(n_1218),
.C(n_1228),
.Y(n_1439)
);

AOI211xp5_ASAP7_75t_L g1440 ( 
.A1(n_1263),
.A2(n_1207),
.B(n_1218),
.C(n_1228),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1269),
.A2(n_1223),
.B(n_1157),
.Y(n_1441)
);

CKINVDCx6p67_ASAP7_75t_R g1442 ( 
.A(n_1264),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1298),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1258),
.B(n_1149),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1258),
.B(n_1149),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_1345),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1258),
.B(n_1149),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1287),
.B(n_1207),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1298),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1280),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1366),
.B(n_1223),
.Y(n_1451)
);

AOI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1390),
.A2(n_1186),
.B1(n_1207),
.B2(n_1303),
.C(n_1382),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1305),
.A2(n_1186),
.B1(n_1409),
.B2(n_1402),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1385),
.A2(n_1186),
.B1(n_1389),
.B2(n_1287),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1382),
.A2(n_1186),
.B1(n_1414),
.B2(n_1419),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1274),
.A2(n_1277),
.B(n_1348),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1281),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1313),
.A2(n_1349),
.B(n_1276),
.C(n_1321),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1350),
.A2(n_1357),
.B(n_1273),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1294),
.A2(n_1361),
.B1(n_1266),
.B2(n_1261),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1264),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1385),
.A2(n_1413),
.B1(n_1295),
.B2(n_1311),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1393),
.B(n_1400),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1259),
.B(n_1346),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1295),
.A2(n_1311),
.B1(n_1374),
.B2(n_1410),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1269),
.A2(n_1416),
.B(n_1262),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1259),
.B(n_1346),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_1371),
.B1(n_1383),
.B2(n_1423),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1325),
.B(n_1360),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1377),
.B(n_1418),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1406),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1340),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1343),
.A2(n_1347),
.B1(n_1351),
.B2(n_1308),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1322),
.B(n_1353),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1396),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1374),
.A2(n_1398),
.B1(n_1296),
.B2(n_1381),
.Y(n_1476)
);

AOI222xp33_ASAP7_75t_L g1477 ( 
.A1(n_1282),
.A2(n_1327),
.B1(n_1302),
.B2(n_1362),
.C1(n_1340),
.C2(n_1314),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1381),
.A2(n_1376),
.B1(n_1397),
.B2(n_1377),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1304),
.B(n_1320),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1286),
.B(n_1289),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1292),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1384),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1329),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1256),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1324),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1293),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1345),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1329),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1387),
.B(n_1402),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1260),
.B(n_1312),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1329),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1384),
.A2(n_1354),
.B1(n_1348),
.B2(n_1387),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1288),
.A2(n_1339),
.B(n_1373),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_SL g1496 ( 
.A(n_1324),
.B(n_1391),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1381),
.A2(n_1344),
.B1(n_1395),
.B2(n_1408),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1344),
.A2(n_1391),
.B1(n_1408),
.B2(n_1332),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1316),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1317),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1395),
.A2(n_1379),
.B1(n_1380),
.B2(n_1392),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_SL g1502 ( 
.A1(n_1335),
.A2(n_1337),
.B(n_1404),
.C(n_1422),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1354),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1323),
.B(n_1328),
.Y(n_1505)
);

INVx4_ASAP7_75t_SL g1506 ( 
.A(n_1403),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1396),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1401),
.B(n_1420),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1396),
.Y(n_1509)
);

INVx5_ASAP7_75t_L g1510 ( 
.A(n_1406),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1421),
.A2(n_1333),
.B1(n_1407),
.B2(n_1331),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1341),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1406),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1395),
.A2(n_1415),
.B(n_1373),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1416),
.A2(n_1262),
.B(n_1405),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1365),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1315),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1405),
.A2(n_1283),
.B(n_1363),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1315),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1417),
.A2(n_1356),
.B1(n_1355),
.B2(n_1358),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1388),
.A2(n_1392),
.B1(n_1380),
.B2(n_1379),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1388),
.A2(n_1367),
.B(n_1352),
.C(n_1359),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1407),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1333),
.A2(n_1309),
.B1(n_1378),
.B2(n_1342),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_R g1526 ( 
.A(n_1378),
.B(n_1310),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1290),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1403),
.B(n_1365),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1270),
.A2(n_1356),
.B1(n_1355),
.B2(n_1358),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1267),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1283),
.A2(n_1363),
.B(n_1339),
.Y(n_1531)
);

CKINVDCx11_ASAP7_75t_R g1532 ( 
.A(n_1403),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1365),
.B(n_1334),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_L g1534 ( 
.A(n_1334),
.B(n_1415),
.C(n_1291),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1365),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1352),
.B(n_1290),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1301),
.B(n_1338),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1365),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1403),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1279),
.Y(n_1540)
);

OAI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1367),
.A2(n_1372),
.B(n_1415),
.C(n_1291),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1270),
.A2(n_1372),
.B1(n_1291),
.B2(n_1265),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1267),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1403),
.Y(n_1544)
);

CKINVDCx16_ASAP7_75t_R g1545 ( 
.A(n_1270),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1372),
.A2(n_1359),
.B1(n_1338),
.B2(n_1336),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1265),
.A2(n_1279),
.B1(n_1300),
.B2(n_1285),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1285),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1307),
.B(n_1336),
.C(n_1306),
.Y(n_1549)
);

NAND2xp33_ASAP7_75t_R g1550 ( 
.A(n_1307),
.B(n_1330),
.Y(n_1550)
);

AOI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1300),
.A2(n_1306),
.B(n_1330),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1284),
.B(n_1319),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1284),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1319),
.A2(n_1003),
.B(n_727),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1275),
.B(n_911),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1275),
.A2(n_1003),
.B(n_727),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1257),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1278),
.A2(n_1044),
.B1(n_1299),
.B2(n_1031),
.Y(n_1558)
);

CKINVDCx8_ASAP7_75t_R g1559 ( 
.A(n_1345),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1256),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1276),
.B(n_911),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1257),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1257),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_SL g1564 ( 
.A(n_1268),
.B(n_727),
.C(n_675),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1369),
.A2(n_842),
.B1(n_1370),
.B2(n_1399),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1399),
.A2(n_1003),
.B(n_727),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1297),
.A2(n_1044),
.B1(n_675),
.B2(n_1003),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_R g1568 ( 
.A(n_1297),
.B(n_899),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1324),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1271),
.B(n_911),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1276),
.B(n_911),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1298),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1368),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1269),
.A2(n_1416),
.B(n_1262),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1375),
.A2(n_1037),
.B1(n_1044),
.B2(n_842),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1399),
.A2(n_1129),
.B(n_1313),
.C(n_1026),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1378),
.B(n_1165),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1271),
.B(n_911),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1384),
.B(n_899),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1274),
.A2(n_729),
.B(n_1112),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1271),
.B(n_911),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1575),
.A2(n_1565),
.B1(n_1424),
.B2(n_1567),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1438),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1564),
.A2(n_1568),
.B1(n_1566),
.B2(n_1437),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1565),
.A2(n_1424),
.B1(n_1558),
.B2(n_1477),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1460),
.A2(n_1453),
.B1(n_1470),
.B2(n_1494),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1459),
.A2(n_1537),
.B(n_1525),
.Y(n_1588)
);

AO21x1_ASAP7_75t_L g1589 ( 
.A1(n_1434),
.A2(n_1473),
.B(n_1440),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1576),
.B(n_1452),
.C(n_1468),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1576),
.A2(n_1428),
.B1(n_1426),
.B2(n_1570),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1470),
.A2(n_1494),
.B1(n_1428),
.B2(n_1507),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1580),
.A2(n_1458),
.B(n_1556),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1426),
.A2(n_1581),
.B1(n_1578),
.B2(n_1462),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1532),
.A2(n_1468),
.B1(n_1462),
.B2(n_1470),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1464),
.B(n_1467),
.Y(n_1596)
);

OAI221xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1458),
.A2(n_1465),
.B1(n_1478),
.B2(n_1476),
.C(n_1434),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1491),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1438),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1485),
.Y(n_1600)
);

CKINVDCx11_ASAP7_75t_R g1601 ( 
.A(n_1559),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1554),
.A2(n_1515),
.B(n_1502),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1532),
.A2(n_1463),
.B1(n_1479),
.B2(n_1425),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_SL g1604 ( 
.A(n_1572),
.B(n_1482),
.C(n_1443),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1479),
.A2(n_1489),
.B1(n_1562),
.B2(n_1450),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1489),
.A2(n_1457),
.B1(n_1557),
.B2(n_1563),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1461),
.A2(n_1476),
.B1(n_1455),
.B2(n_1442),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1461),
.A2(n_1485),
.B1(n_1496),
.B2(n_1474),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1481),
.A2(n_1486),
.B1(n_1454),
.B2(n_1555),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1475),
.A2(n_1507),
.B1(n_1504),
.B2(n_1435),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1454),
.A2(n_1444),
.B1(n_1445),
.B2(n_1447),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1504),
.A2(n_1579),
.B1(n_1444),
.B2(n_1447),
.C1(n_1445),
.C2(n_1528),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1502),
.A2(n_1456),
.B(n_1537),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1427),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1432),
.A2(n_1439),
.B(n_1511),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1568),
.A2(n_1492),
.B1(n_1569),
.B2(n_1436),
.Y(n_1616)
);

AO21x1_ASAP7_75t_L g1617 ( 
.A1(n_1498),
.A2(n_1533),
.B(n_1433),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1465),
.A2(n_1498),
.B1(n_1544),
.B2(n_1539),
.C(n_1478),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1480),
.Y(n_1619)
);

AOI322xp5_ASAP7_75t_L g1620 ( 
.A1(n_1545),
.A2(n_1430),
.A3(n_1517),
.B1(n_1535),
.B2(n_1538),
.C1(n_1497),
.C2(n_1449),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1509),
.A2(n_1472),
.B1(n_1573),
.B2(n_1518),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1475),
.A2(n_1500),
.B1(n_1499),
.B2(n_1509),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1520),
.A2(n_1431),
.B1(n_1451),
.B2(n_1506),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1491),
.A2(n_1483),
.B1(n_1488),
.B2(n_1495),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1505),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1451),
.A2(n_1506),
.B1(n_1560),
.B2(n_1484),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1506),
.A2(n_1456),
.B1(n_1503),
.B2(n_1522),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1501),
.A2(n_1523),
.B1(n_1524),
.B2(n_1488),
.C(n_1495),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1501),
.A2(n_1523),
.B1(n_1483),
.B2(n_1497),
.C(n_1529),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1490),
.B(n_1508),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1487),
.A2(n_1577),
.B1(n_1529),
.B2(n_1510),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1508),
.B(n_1514),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1577),
.A2(n_1510),
.B1(n_1429),
.B2(n_1514),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1512),
.B(n_1471),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1548),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1521),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1446),
.A2(n_1526),
.B1(n_1512),
.B2(n_1527),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1521),
.A2(n_1534),
.B1(n_1526),
.B2(n_1542),
.C(n_1541),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1510),
.B(n_1471),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1446),
.A2(n_1471),
.B1(n_1536),
.B2(n_1510),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1542),
.A2(n_1551),
.B1(n_1540),
.B2(n_1549),
.C(n_1547),
.Y(n_1642)
);

AOI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1550),
.A2(n_1552),
.B(n_1546),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1471),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1553),
.A2(n_1530),
.B1(n_1543),
.B2(n_1493),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1493),
.B(n_1519),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1547),
.A2(n_1441),
.B1(n_1516),
.B2(n_1466),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1574),
.A2(n_1531),
.B1(n_1564),
.B2(n_842),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1564),
.A2(n_770),
.B1(n_727),
.B2(n_1268),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1575),
.A2(n_1044),
.B1(n_1565),
.B2(n_1299),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1564),
.A2(n_770),
.B1(n_727),
.B2(n_1268),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1575),
.A2(n_1564),
.B(n_1268),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1474),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1575),
.A2(n_1044),
.B1(n_1565),
.B2(n_1299),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1566),
.A2(n_727),
.B1(n_1575),
.B2(n_1268),
.C(n_1564),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1461),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1564),
.A2(n_561),
.B1(n_1163),
.B2(n_1566),
.C(n_673),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1567),
.A2(n_1375),
.B1(n_1044),
.B2(n_979),
.Y(n_1662)
);

OAI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1575),
.A2(n_1424),
.B(n_561),
.C(n_500),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1564),
.A2(n_1268),
.B(n_727),
.C(n_1163),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1564),
.A2(n_561),
.B1(n_1163),
.B2(n_1566),
.C(n_673),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1513),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1464),
.B(n_1467),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1566),
.A2(n_727),
.B1(n_1575),
.B2(n_1268),
.C(n_1564),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1564),
.A2(n_561),
.B1(n_1163),
.B2(n_1566),
.C(n_673),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1448),
.B(n_1469),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1469),
.B(n_1570),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1675)
);

AOI21xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1567),
.A2(n_649),
.B(n_633),
.Y(n_1676)
);

NAND4xp25_ASAP7_75t_L g1677 ( 
.A(n_1424),
.B(n_914),
.C(n_673),
.D(n_590),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1424),
.B(n_914),
.C(n_673),
.D(n_590),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1444),
.B(n_1445),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1564),
.A2(n_561),
.B1(n_1163),
.B2(n_1566),
.C(n_673),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1448),
.B(n_1469),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1448),
.B(n_1469),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1575),
.A2(n_1044),
.B1(n_1565),
.B2(n_1299),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1510),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1469),
.B(n_1570),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_SL g1690 ( 
.A1(n_1566),
.A2(n_1037),
.B1(n_1375),
.B2(n_1044),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1561),
.B(n_1571),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1566),
.B(n_727),
.C(n_1268),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1513),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1469),
.B(n_1570),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1531),
.A2(n_1574),
.B(n_1466),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1696)
);

OAI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1575),
.A2(n_1424),
.B(n_561),
.C(n_500),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1566),
.A2(n_1037),
.B1(n_1375),
.B2(n_1044),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1470),
.B(n_1479),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1531),
.A2(n_1574),
.B(n_1466),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1567),
.A2(n_1375),
.B1(n_1044),
.B2(n_979),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1564),
.A2(n_842),
.B1(n_1575),
.B2(n_1565),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1636),
.Y(n_1704)
);

CKINVDCx6p67_ASAP7_75t_R g1705 ( 
.A(n_1700),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1672),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1645),
.B(n_1646),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1645),
.B(n_1646),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1611),
.B(n_1609),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1611),
.B(n_1609),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1683),
.B(n_1685),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1666),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1695),
.B(n_1701),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1614),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1643),
.B(n_1628),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1628),
.B(n_1642),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1583),
.A2(n_1586),
.B1(n_1655),
.B2(n_1657),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1588),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1700),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1590),
.B(n_1613),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1656),
.B(n_1670),
.Y(n_1722)
);

BUFx2_ASAP7_75t_SL g1723 ( 
.A(n_1589),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1637),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1602),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_L g1727 ( 
.A(n_1615),
.B(n_1692),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1647),
.B(n_1593),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1595),
.B(n_1648),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1648),
.B(n_1639),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1630),
.Y(n_1731)
);

OA21x2_ASAP7_75t_L g1732 ( 
.A1(n_1617),
.A2(n_1627),
.B(n_1607),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1585),
.B(n_1629),
.Y(n_1734)
);

AOI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1632),
.A2(n_1591),
.B(n_1594),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1619),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1626),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1631),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1596),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1586),
.A2(n_1703),
.B1(n_1699),
.B2(n_1657),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1664),
.B(n_1659),
.C(n_1665),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1596),
.Y(n_1742)
);

NAND2x1_ASAP7_75t_L g1743 ( 
.A(n_1688),
.B(n_1624),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1587),
.B(n_1620),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1668),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1641),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1603),
.B(n_1605),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1597),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1603),
.B(n_1605),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1606),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1606),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1644),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1612),
.B(n_1592),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1584),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1633),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1582),
.B(n_1691),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1638),
.B(n_1653),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1634),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1635),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1741),
.A2(n_1652),
.B1(n_1718),
.B2(n_1651),
.C(n_1649),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1706),
.B(n_1669),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1667),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1706),
.B(n_1711),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1722),
.A2(n_1703),
.B1(n_1699),
.B2(n_1696),
.Y(n_1764)
);

NAND3xp33_ASAP7_75t_SL g1765 ( 
.A(n_1741),
.B(n_1676),
.C(n_1671),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1704),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1741),
.A2(n_1697),
.B1(n_1663),
.B2(n_1650),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_R g1768 ( 
.A(n_1735),
.B(n_1600),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1722),
.A2(n_1682),
.B(n_1686),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1718),
.A2(n_1740),
.B1(n_1679),
.B2(n_1675),
.C(n_1674),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1752),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1754),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1725),
.B(n_1622),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1723),
.A2(n_1690),
.B1(n_1698),
.B2(n_1679),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1713),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1712),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1738),
.Y(n_1779)
);

AO221x1_ASAP7_75t_L g1780 ( 
.A1(n_1731),
.A2(n_1702),
.B1(n_1662),
.B2(n_1687),
.C(n_1654),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1727),
.A2(n_1696),
.B1(n_1675),
.B2(n_1674),
.C(n_1661),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1712),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1752),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1744),
.A2(n_1686),
.B1(n_1684),
.B2(n_1655),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1738),
.Y(n_1785)
);

OAI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1743),
.A2(n_1623),
.B(n_1598),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1740),
.A2(n_1661),
.B1(n_1660),
.B2(n_1684),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1711),
.B(n_1694),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1721),
.A2(n_1660),
.B(n_1673),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1754),
.Y(n_1790)
);

AOI221x1_ASAP7_75t_L g1791 ( 
.A1(n_1723),
.A2(n_1678),
.B1(n_1677),
.B2(n_1689),
.C(n_1598),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1715),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1744),
.A2(n_1610),
.B1(n_1658),
.B2(n_1604),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1719),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1616),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1744),
.A2(n_1608),
.B1(n_1621),
.B2(n_1658),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1725),
.B(n_1719),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1755),
.B(n_1599),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1742),
.B(n_1599),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1744),
.A2(n_1608),
.B1(n_1625),
.B2(n_1622),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1714),
.B(n_1640),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1713),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1754),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1742),
.B(n_1601),
.Y(n_1805)
);

AO21x2_ASAP7_75t_L g1806 ( 
.A1(n_1721),
.A2(n_1713),
.B(n_1730),
.Y(n_1806)
);

NAND4xp25_ASAP7_75t_L g1807 ( 
.A(n_1727),
.B(n_1748),
.C(n_1734),
.D(n_1721),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1742),
.B(n_1745),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1734),
.A2(n_1748),
.B1(n_1723),
.B2(n_1727),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1721),
.B(n_1734),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1752),
.Y(n_1811)
);

OAI33xp33_ASAP7_75t_L g1812 ( 
.A1(n_1748),
.A2(n_1731),
.A3(n_1724),
.B1(n_1757),
.B2(n_1750),
.B3(n_1751),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1731),
.A2(n_1735),
.B1(n_1726),
.B2(n_1730),
.C(n_1753),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1806),
.B(n_1707),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1766),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1763),
.B(n_1736),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1778),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1778),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1806),
.B(n_1707),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1810),
.B(n_1720),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1806),
.B(n_1707),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1779),
.B(n_1736),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1797),
.B(n_1707),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1782),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1797),
.B(n_1708),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1772),
.B(n_1728),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_R g1827 ( 
.A(n_1765),
.B(n_1735),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1797),
.B(n_1708),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1797),
.B(n_1708),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1808),
.B(n_1708),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1810),
.B(n_1737),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1783),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1798),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1780),
.A2(n_1726),
.B1(n_1747),
.B2(n_1749),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1773),
.B(n_1728),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1773),
.B(n_1794),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1794),
.B(n_1728),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1789),
.B(n_1737),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1807),
.B(n_1758),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1789),
.B(n_1737),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1798),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1777),
.Y(n_1842)
);

AND2x4_ASAP7_75t_SL g1843 ( 
.A(n_1775),
.B(n_1705),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1789),
.B(n_1737),
.Y(n_1844)
);

AND2x2_ASAP7_75t_SL g1845 ( 
.A(n_1789),
.B(n_1732),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1811),
.B(n_1752),
.Y(n_1846)
);

AND2x2_ASAP7_75t_SL g1847 ( 
.A(n_1784),
.B(n_1732),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1819),
.B(n_1821),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1823),
.B(n_1762),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1826),
.B(n_1761),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1817),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1852)
);

NAND2x1p5_ASAP7_75t_L g1853 ( 
.A(n_1820),
.B(n_1786),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1815),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1823),
.B(n_1762),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1817),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1818),
.Y(n_1858)
);

INVxp33_ASAP7_75t_L g1859 ( 
.A(n_1827),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1825),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1760),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1839),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1826),
.B(n_1761),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1770),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1831),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1775),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1833),
.B(n_1807),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1821),
.B(n_1770),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1815),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1825),
.B(n_1775),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1821),
.B(n_1730),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1826),
.B(n_1755),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1775),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1833),
.B(n_1755),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1825),
.B(n_1799),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_SL g1876 ( 
.A(n_1827),
.B(n_1769),
.C(n_1767),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1818),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1828),
.B(n_1799),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1818),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1841),
.B(n_1792),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1814),
.B(n_1730),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1824),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1841),
.B(n_1792),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1828),
.B(n_1829),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1815),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1828),
.B(n_1802),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1824),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_SL g1888 ( 
.A(n_1820),
.B(n_1814),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1838),
.B(n_1801),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1824),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1854),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1890),
.Y(n_1892)
);

BUFx4f_ASAP7_75t_L g1893 ( 
.A(n_1853),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1854),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1888),
.B(n_1866),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1853),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1888),
.B(n_1866),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1890),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1870),
.B(n_1828),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1861),
.B(n_1813),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1851),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1859),
.B(n_1768),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1876),
.B(n_1785),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_SL g1904 ( 
.A(n_1876),
.B(n_1809),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_R g1905 ( 
.A(n_1867),
.B(n_1732),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1854),
.Y(n_1906)
);

OAI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1862),
.A2(n_1847),
.B(n_1834),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1889),
.B(n_1838),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1889),
.B(n_1840),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1862),
.B(n_1847),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1881),
.B(n_1776),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1887),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1829),
.Y(n_1913)
);

NAND2xp33_ASAP7_75t_R g1914 ( 
.A(n_1881),
.B(n_1732),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1887),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1871),
.A2(n_1847),
.B1(n_1776),
.B2(n_1834),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1851),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1871),
.B(n_1864),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1852),
.B(n_1847),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1869),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1856),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1860),
.B(n_1829),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1852),
.A2(n_1780),
.B1(n_1781),
.B2(n_1787),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1869),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1864),
.B(n_1840),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1849),
.B(n_1795),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1853),
.B(n_1845),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1874),
.B(n_1812),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1873),
.B(n_1796),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_R g1930 ( 
.A(n_1873),
.B(n_1732),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1868),
.B(n_1844),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1869),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1868),
.B(n_1844),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1849),
.B(n_1814),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1856),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1916),
.A2(n_1784),
.B(n_1793),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1923),
.A2(n_1764),
.B1(n_1771),
.B2(n_1845),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1911),
.A2(n_1907),
.B1(n_1900),
.B2(n_1904),
.C(n_1910),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1902),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1895),
.B(n_1875),
.Y(n_1940)
);

AOI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1911),
.A2(n_1814),
.B1(n_1848),
.B2(n_1865),
.C(n_1717),
.Y(n_1941)
);

OAI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1905),
.A2(n_1791),
.B1(n_1800),
.B2(n_1753),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_L g1943 ( 
.A(n_1914),
.B(n_1791),
.C(n_1845),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1895),
.B(n_1875),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1903),
.A2(n_1845),
.B(n_1726),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1922),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1927),
.A2(n_1848),
.B1(n_1865),
.B2(n_1717),
.C(n_1716),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1897),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1921),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1922),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1893),
.A2(n_1800),
.B1(n_1753),
.B2(n_1717),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1922),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1921),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1926),
.B(n_1855),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1893),
.A2(n_1753),
.B1(n_1717),
.B2(n_1716),
.Y(n_1955)
);

OAI22x1_ASAP7_75t_L g1956 ( 
.A1(n_1929),
.A2(n_1805),
.B1(n_1884),
.B2(n_1860),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1930),
.A2(n_1928),
.B1(n_1897),
.B2(n_1716),
.Y(n_1957)
);

OAI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1919),
.A2(n_1716),
.B(n_1726),
.Y(n_1958)
);

AO22x2_ASAP7_75t_L g1959 ( 
.A1(n_1892),
.A2(n_1842),
.B1(n_1882),
.B2(n_1858),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1899),
.Y(n_1960)
);

AOI222xp33_ASAP7_75t_L g1961 ( 
.A1(n_1893),
.A2(n_1749),
.B1(n_1747),
.B2(n_1729),
.C1(n_1710),
.C2(n_1709),
.Y(n_1961)
);

OAI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1896),
.A2(n_1732),
.B1(n_1720),
.B2(n_1705),
.Y(n_1962)
);

AOI211xp5_ASAP7_75t_L g1963 ( 
.A1(n_1896),
.A2(n_1749),
.B(n_1747),
.C(n_1729),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1918),
.B(n_1855),
.Y(n_1964)
);

OAI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1918),
.A2(n_1732),
.B1(n_1720),
.B2(n_1705),
.Y(n_1965)
);

XNOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1899),
.B(n_1805),
.Y(n_1966)
);

AOI21xp33_ASAP7_75t_L g1967 ( 
.A1(n_1908),
.A2(n_1804),
.B(n_1758),
.Y(n_1967)
);

INVxp67_ASAP7_75t_L g1968 ( 
.A(n_1935),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1913),
.B(n_1878),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1908),
.A2(n_1831),
.B(n_1747),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1898),
.A2(n_1749),
.B(n_1901),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1909),
.B(n_1878),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1949),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1937),
.A2(n_1758),
.B1(n_1729),
.B2(n_1709),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1949),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1942),
.A2(n_1909),
.B(n_1933),
.C(n_1931),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1953),
.Y(n_1977)
);

NAND4xp25_ASAP7_75t_SL g1978 ( 
.A(n_1938),
.B(n_1934),
.C(n_1931),
.D(n_1925),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1948),
.B(n_1913),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1940),
.B(n_1884),
.Y(n_1980)
);

OAI221xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1936),
.A2(n_1933),
.B1(n_1925),
.B2(n_1729),
.C(n_1709),
.Y(n_1981)
);

OAI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1942),
.A2(n_1720),
.B1(n_1705),
.B2(n_1746),
.Y(n_1982)
);

AND2x4_ASAP7_75t_SL g1983 ( 
.A(n_1946),
.B(n_1756),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1941),
.A2(n_1710),
.B1(n_1709),
.B2(n_1733),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1939),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1956),
.B(n_1874),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1961),
.B(n_1829),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1944),
.B(n_1886),
.Y(n_1988)
);

OAI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1957),
.A2(n_1943),
.B(n_1947),
.C(n_1945),
.Y(n_1989)
);

NAND3xp33_ASAP7_75t_L g1990 ( 
.A(n_1963),
.B(n_1935),
.C(n_1915),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1958),
.B(n_1850),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1955),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1968),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1951),
.A2(n_1733),
.B(n_1710),
.C(n_1786),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1954),
.B(n_1966),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1968),
.Y(n_1996)
);

AOI322xp5_ASAP7_75t_L g1997 ( 
.A1(n_1965),
.A2(n_1710),
.A3(n_1837),
.B1(n_1835),
.B2(n_1830),
.C1(n_1733),
.C2(n_1886),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1950),
.B(n_1830),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1959),
.Y(n_1999)
);

OAI22x1_ASAP7_75t_L g2000 ( 
.A1(n_1952),
.A2(n_1912),
.B1(n_1917),
.B2(n_1774),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1975),
.Y(n_2001)
);

NOR3xp33_ASAP7_75t_SL g2002 ( 
.A(n_1978),
.B(n_1965),
.C(n_1962),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1975),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1973),
.Y(n_2004)
);

AOI322xp5_ASAP7_75t_L g2005 ( 
.A1(n_1992),
.A2(n_1962),
.A3(n_1972),
.B1(n_1967),
.B2(n_1964),
.C1(n_1960),
.C2(n_1733),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1985),
.B(n_1972),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1992),
.B(n_1970),
.Y(n_2007)
);

NOR2x1_ASAP7_75t_L g2008 ( 
.A(n_1993),
.B(n_1971),
.Y(n_2008)
);

OR3x1_ASAP7_75t_L g2009 ( 
.A(n_1999),
.B(n_1877),
.C(n_1857),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1979),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1980),
.B(n_1969),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1998),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1982),
.B(n_1976),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1996),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1988),
.B(n_1959),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1996),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_SL g2017 ( 
.A(n_1989),
.B(n_1774),
.C(n_1759),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1977),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1983),
.B(n_1959),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1974),
.B(n_1756),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2010),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_L g2022 ( 
.A1(n_2008),
.A2(n_1982),
.B(n_2000),
.Y(n_2022)
);

NAND3xp33_ASAP7_75t_L g2023 ( 
.A(n_2003),
.B(n_2016),
.C(n_2014),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_2010),
.Y(n_2024)
);

INVx4_ASAP7_75t_L g2025 ( 
.A(n_2014),
.Y(n_2025)
);

NOR2x1p5_ASAP7_75t_L g2026 ( 
.A(n_2006),
.B(n_1995),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2016),
.B(n_1984),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2001),
.B(n_2011),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_2017),
.B(n_1994),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_2019),
.Y(n_2030)
);

NAND5xp2_ASAP7_75t_L g2031 ( 
.A(n_2002),
.B(n_1981),
.C(n_1997),
.D(n_1987),
.E(n_1994),
.Y(n_2031)
);

OAI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2022),
.A2(n_2013),
.B(n_2008),
.C(n_2005),
.Y(n_2032)
);

NAND2xp33_ASAP7_75t_SL g2033 ( 
.A(n_2026),
.B(n_2007),
.Y(n_2033)
);

NOR4xp25_ASAP7_75t_L g2034 ( 
.A(n_2023),
.B(n_2001),
.C(n_2004),
.D(n_2018),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2030),
.B(n_2004),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_L g2036 ( 
.A(n_2023),
.B(n_2018),
.C(n_1986),
.Y(n_2036)
);

AOI321xp33_ASAP7_75t_L g2037 ( 
.A1(n_2029),
.A2(n_2012),
.A3(n_2015),
.B1(n_2011),
.B2(n_2019),
.C(n_2005),
.Y(n_2037)
);

AOI21xp33_ASAP7_75t_L g2038 ( 
.A1(n_2028),
.A2(n_2012),
.B(n_1990),
.Y(n_2038)
);

OAI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_2027),
.A2(n_1991),
.B1(n_2020),
.B2(n_2015),
.C(n_2009),
.Y(n_2039)
);

OAI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2025),
.A2(n_2009),
.B(n_1932),
.Y(n_2040)
);

NOR4xp25_ASAP7_75t_SL g2041 ( 
.A(n_2030),
.B(n_1879),
.C(n_1857),
.D(n_1858),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_2033),
.B(n_2025),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2036),
.B(n_2024),
.Y(n_2043)
);

OAI211xp5_ASAP7_75t_SL g2044 ( 
.A1(n_2032),
.A2(n_2021),
.B(n_2031),
.C(n_1932),
.Y(n_2044)
);

O2A1O1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_2034),
.A2(n_1924),
.B(n_1920),
.C(n_1906),
.Y(n_2045)
);

AOI221x1_ASAP7_75t_L g2046 ( 
.A1(n_2035),
.A2(n_1924),
.B1(n_1920),
.B2(n_1891),
.C(n_1906),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2038),
.B(n_1756),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_2044),
.B(n_2039),
.Y(n_2048)
);

O2A1O1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_2042),
.A2(n_2040),
.B(n_2037),
.C(n_2041),
.Y(n_2049)
);

NAND4xp75_ASAP7_75t_L g2050 ( 
.A(n_2043),
.B(n_1894),
.C(n_1891),
.D(n_1835),
.Y(n_2050)
);

NAND3x1_ASAP7_75t_L g2051 ( 
.A(n_2047),
.B(n_1882),
.C(n_1879),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2045),
.Y(n_2052)
);

OR5x1_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_1894),
.C(n_1885),
.D(n_1842),
.E(n_1877),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2047),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2048),
.B(n_1850),
.Y(n_2055)
);

OAI211xp5_ASAP7_75t_L g2056 ( 
.A1(n_2049),
.A2(n_1743),
.B(n_1863),
.C(n_1832),
.Y(n_2056)
);

OAI221xp5_ASAP7_75t_L g2057 ( 
.A1(n_2052),
.A2(n_1743),
.B1(n_1863),
.B2(n_1842),
.C(n_1746),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2054),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2050),
.B(n_1880),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2051),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2055),
.B(n_1830),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2058),
.B(n_1830),
.Y(n_2062)
);

XNOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2060),
.B(n_2053),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_2056),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2062),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2065),
.A2(n_2064),
.B1(n_2057),
.B2(n_2059),
.C(n_2061),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2066),
.A2(n_2064),
.B1(n_2063),
.B2(n_1842),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2066),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2067),
.A2(n_1883),
.B(n_1880),
.Y(n_2069)
);

AOI222xp33_ASAP7_75t_L g2070 ( 
.A1(n_2068),
.A2(n_1885),
.B1(n_1832),
.B2(n_1746),
.C1(n_1836),
.C2(n_1822),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2069),
.A2(n_1885),
.B1(n_1883),
.B2(n_1872),
.Y(n_2071)
);

OAI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2070),
.A2(n_1872),
.B1(n_1822),
.B2(n_1816),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_2071),
.A2(n_1746),
.B1(n_1790),
.B2(n_1803),
.Y(n_2073)
);

OAI221xp5_ASAP7_75t_R g2074 ( 
.A1(n_2073),
.A2(n_2072),
.B1(n_1843),
.B2(n_1836),
.C(n_1846),
.Y(n_2074)
);

AOI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_2074),
.A2(n_1757),
.B(n_1837),
.C(n_1835),
.Y(n_2075)
);


endmodule