module real_jpeg_24516_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_348, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_348;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_47),
.B1(n_58),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx8_ASAP7_75t_SL g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_5),
.A2(n_66),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_84),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_128),
.B1(n_151),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_33),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_59),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_116),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_116),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_47),
.B1(n_58),
.B2(n_116),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_42),
.B1(n_58),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_42),
.B1(n_70),
.B2(n_71),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_235)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_10),
.A2(n_70),
.B1(n_71),
.B2(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_125),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_10),
.A2(n_81),
.B1(n_125),
.B2(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_70),
.B1(n_71),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_133),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_133),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_11),
.A2(n_58),
.B1(n_133),
.B2(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_50),
.B1(n_70),
.B2(n_71),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_50),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_14),
.A2(n_37),
.B1(n_70),
.B2(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_14),
.A2(n_37),
.B1(n_219),
.B2(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_15),
.Y(n_131)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_15),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_100),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_98),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_19),
.B(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_75),
.B2(n_86),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_62),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_22),
.A2(n_23),
.B1(n_62),
.B2(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_25),
.A2(n_39),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_26),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_26),
.A2(n_38),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_27),
.A2(n_29),
.A3(n_33),
.B1(n_171),
.B2(n_180),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_28),
.B(n_31),
.Y(n_180)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_29),
.A2(n_68),
.B(n_112),
.C(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_32),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_32),
.A2(n_97),
.B(n_172),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_33),
.B(n_55),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_34),
.B(n_112),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_34),
.A2(n_46),
.A3(n_54),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_39),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_39),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_39),
.A2(n_84),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_39),
.A2(n_84),
.B1(n_195),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_39),
.A2(n_84),
.B1(n_95),
.B2(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_84),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_43),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_53),
.B(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_47),
.A2(n_112),
.B(n_218),
.Y(n_237)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_48),
.Y(n_219)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_60),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_51),
.A2(n_59),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_51),
.A2(n_59),
.B1(n_238),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_52),
.A2(n_53),
.B1(n_250),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_52),
.A2(n_266),
.B(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_52),
.A2(n_79),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_58),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_59),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_62),
.A2(n_63),
.B1(n_94),
.B2(n_334),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_91),
.C(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_73),
.B(n_74),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_64),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_64),
.A2(n_73),
.B1(n_115),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_64),
.A2(n_73),
.B1(n_124),
.B2(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_64),
.A2(n_74),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_64),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_69),
.B(n_112),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_69),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_69),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_69),
.A2(n_113),
.B1(n_257),
.B2(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_70),
.B(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_73),
.B(n_74),
.Y(n_208)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_81),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.C(n_93),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_91),
.A2(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_91),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_93),
.B(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_94),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_329),
.A3(n_340),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_100)
);

AOI311xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_280),
.A3(n_320),
.B(n_323),
.C(n_324),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_240),
.C(n_275),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_212),
.B(n_239),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_188),
.B(n_211),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_164),
.B(n_187),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_138),
.B(n_163),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_108),
.B(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_117),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_110),
.B1(n_117),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_112),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_113),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_113),
.A2(n_273),
.B(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_126),
.C(n_127),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B(n_134),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_137),
.B1(n_142),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_128),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_128),
.A2(n_183),
.B(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_128),
.A2(n_182),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_129),
.B(n_184),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_136),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_131),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_131),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_134),
.B(n_202),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_147),
.B(n_162),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_145),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_152),
.B(n_161),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_165),
.B(n_166),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_178),
.B1(n_185),
.B2(n_186),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_177),
.C(n_185),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_203),
.B2(n_204),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_206),
.C(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_198),
.C(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_208),
.B(n_258),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_214),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_229),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_216),
.B(n_228),
.C(n_229),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_224),
.Y(n_245)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_233),
.C(n_236),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_241),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_260),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_242),
.B(n_260),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_252),
.C(n_253),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_244),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_247),
.C(n_248),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_253),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_256),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_260),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_270),
.CI(n_274),
.CON(n_260),
.SN(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_269),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_277),
.Y(n_326)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_281),
.A2(n_321),
.B(n_325),
.C(n_328),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_302),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_282),
.B(n_322),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_290),
.CI(n_301),
.CON(n_282),
.SN(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_289),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_287),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_289),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_310),
.B(n_314),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_300),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_294),
.C(n_298),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_296),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_299),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_319),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_309),
.B1(n_317),
.B2(n_318),
.Y(n_303)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_307),
.B(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_331),
.B1(n_336),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_317),
.C(n_319),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_338),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_338),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.C(n_337),
.Y(n_330)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_331),
.Y(n_344)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);


endmodule