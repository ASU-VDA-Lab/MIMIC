module fake_jpeg_14479_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_49),
.B(n_55),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_60),
.B1(n_46),
.B2(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_34),
.B1(n_30),
.B2(n_20),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_44),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_64),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_46),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_20),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_36),
.B1(n_21),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_23),
.B1(n_22),
.B2(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_74),
.A2(n_91),
.B1(n_109),
.B2(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_86),
.Y(n_119)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_0),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_101),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_44),
.B1(n_39),
.B2(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_96),
.Y(n_140)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_0),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_22),
.B(n_27),
.C(n_28),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_106),
.B(n_53),
.C(n_66),
.Y(n_133)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_8),
.Y(n_143)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_58),
.B1(n_23),
.B2(n_35),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_70),
.C(n_66),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_126),
.Y(n_147)
);

OAI22x1_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_53),
.B1(n_66),
.B2(n_58),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_135),
.B1(n_104),
.B2(n_110),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_5),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_143),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_83),
.B1(n_106),
.B2(n_99),
.Y(n_135)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_7),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_88),
.B(n_79),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_149),
.B(n_171),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_151),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_80),
.B(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_165),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_106),
.B1(n_109),
.B2(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_155),
.B1(n_161),
.B2(n_166),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_106),
.B1(n_95),
.B2(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_89),
.B1(n_75),
.B2(n_98),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_174),
.Y(n_199)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_75),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_78),
.B1(n_103),
.B2(n_112),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_84),
.B1(n_100),
.B2(n_93),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_124),
.B1(n_132),
.B2(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_128),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_136),
.B1(n_124),
.B2(n_144),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_118),
.A2(n_9),
.B(n_10),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_9),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2x1_ASAP7_75t_SL g175 ( 
.A(n_116),
.B(n_12),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_141),
.B(n_126),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_12),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_184),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_128),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_129),
.A3(n_132),
.B1(n_130),
.B2(n_115),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_130),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_200),
.B(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_115),
.B1(n_137),
.B2(n_14),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_12),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_204),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_15),
.B1(n_16),
.B2(n_152),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_154),
.C(n_149),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_169),
.C(n_158),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_215),
.C(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_148),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_217),
.Y(n_242)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_177),
.C(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_227),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_184),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_161),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_230),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_180),
.A2(n_176),
.B(n_167),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_232),
.B(n_175),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_180),
.A2(n_176),
.B(n_162),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_203),
.B1(n_196),
.B2(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_198),
.B1(n_201),
.B2(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_196),
.B1(n_177),
.B2(n_178),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_246),
.B1(n_249),
.B2(n_221),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_233),
.B1(n_211),
.B2(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_198),
.B1(n_197),
.B2(n_204),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_175),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_225),
.A2(n_198),
.B1(n_166),
.B2(n_185),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_231),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_150),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_205),
.B1(n_206),
.B2(n_181),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_222),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_232),
.B(n_248),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_227),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_221),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_283),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_237),
.C(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_233),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_247),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_267),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_239),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_228),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_249),
.C(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_257),
.C(n_259),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_271),
.B(n_268),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_294),
.B(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_257),
.B1(n_269),
.B2(n_236),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_284),
.B1(n_209),
.B2(n_273),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_259),
.C(n_261),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_270),
.C(n_250),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_273),
.C(n_263),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_281),
.B(n_279),
.C(n_285),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_291),
.B1(n_295),
.B2(n_287),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_243),
.B(n_245),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_212),
.B(n_229),
.Y(n_309)
);

OAI221xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_309),
.B1(n_308),
.B2(n_226),
.C(n_220),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_287),
.B(n_212),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_300),
.A3(n_255),
.B1(n_298),
.B2(n_214),
.C1(n_218),
.C2(n_224),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_312),
.B1(n_206),
.B2(n_172),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_219),
.B(n_216),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_314),
.Y(n_316)
);

OAI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_315),
.A3(n_214),
.B1(n_159),
.B2(n_190),
.C(n_164),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule