module fake_jpeg_5848_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_41),
.B1(n_31),
.B2(n_34),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_29),
.B(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_15),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_40),
.B1(n_39),
.B2(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_50),
.B1(n_61),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_39),
.B1(n_21),
.B2(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_63),
.B1(n_61),
.B2(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_75),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_76),
.B(n_84),
.C(n_42),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_22),
.B1(n_24),
.B2(n_29),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_29),
.B1(n_32),
.B2(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_52),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_100),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_108),
.B1(n_81),
.B2(n_76),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_99),
.B1(n_74),
.B2(n_64),
.Y(n_121)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_97),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_53),
.C(n_42),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_46),
.B1(n_58),
.B2(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_48),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_56),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_104),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_42),
.C(n_45),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_51),
.C(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_80),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_93),
.Y(n_151)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_70),
.B1(n_82),
.B2(n_75),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_126),
.B1(n_132),
.B2(n_92),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_70),
.B1(n_87),
.B2(n_94),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_122),
.B1(n_91),
.B2(n_108),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_131),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_105),
.B(n_88),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_81),
.B1(n_67),
.B2(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_67),
.B1(n_72),
.B2(n_71),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_123),
.B1(n_117),
.B2(n_17),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_146),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_127),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_156),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_95),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_145),
.C(n_114),
.Y(n_170)
);

AO21x2_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_103),
.B(n_102),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_133),
.B1(n_124),
.B2(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_93),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_158),
.B1(n_132),
.B2(n_121),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_104),
.C(n_103),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_153),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_152),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_110),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_90),
.B1(n_54),
.B2(n_60),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_183),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_133),
.B1(n_119),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_135),
.B1(n_155),
.B2(n_158),
.Y(n_204)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_174),
.B1(n_180),
.B2(n_181),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_116),
.B1(n_126),
.B2(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_154),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_119),
.C(n_110),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_113),
.A3(n_123),
.B1(n_85),
.B2(n_51),
.C1(n_54),
.C2(n_29),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_54),
.B1(n_17),
.B2(n_30),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_140),
.C(n_142),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_30),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_54),
.C(n_18),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_135),
.C(n_156),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_146),
.B1(n_150),
.B2(n_152),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_192),
.B(n_20),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_193),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_197),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_150),
.B1(n_152),
.B2(n_144),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_134),
.B1(n_137),
.B2(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_183),
.B1(n_23),
.B2(n_18),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_134),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_208),
.B1(n_210),
.B2(n_168),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_147),
.C(n_14),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_147),
.B1(n_17),
.B2(n_30),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_18),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_18),
.B(n_23),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_182),
.C(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_177),
.C(n_169),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_186),
.C(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_172),
.C(n_179),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_219),
.C(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_179),
.C(n_176),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_233),
.B1(n_196),
.B2(n_188),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_18),
.C(n_23),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_23),
.C(n_17),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_210),
.C(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_187),
.B(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_0),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_208),
.B1(n_192),
.B2(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_243),
.B(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_245),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_213),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_246),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_238),
.C(n_215),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_231),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_205),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_219),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_13),
.B(n_12),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_1),
.B(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_230),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_3),
.C(n_4),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_220),
.B(n_226),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_261),
.B(n_268),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_223),
.C(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_247),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_228),
.B(n_221),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_11),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_12),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_267),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_11),
.C(n_2),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_11),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_255),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_243),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_276),
.B(n_278),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_234),
.B(n_248),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_283),
.C(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_296),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_262),
.C(n_5),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_4),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_10),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_286),
.B(n_289),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_299),
.B(n_304),
.Y(n_308)
);

AOI221xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_285),
.B1(n_272),
.B2(n_283),
.C(n_275),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

OA21x2_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_6),
.B(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_295),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_8),
.B(n_9),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_310),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_8),
.C(n_9),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_299),
.C1(n_309),
.C2(n_313),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.C(n_10),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_311),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_10),
.Y(n_317)
);


endmodule