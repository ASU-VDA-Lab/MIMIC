module real_aes_7853_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_1), .A2(n_137), .B(n_141), .C(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_2), .A2(n_173), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g461 ( .A(n_3), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_4), .B(n_213), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g488 ( .A1(n_5), .A2(n_173), .B(n_489), .Y(n_488) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g196 ( .A(n_7), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_8), .B(n_40), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_9), .A2(n_172), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_10), .B(n_149), .Y(n_240) );
INVx1_ASAP7_75t_L g493 ( .A(n_11), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_12), .B(n_207), .Y(n_516) );
INVx1_ASAP7_75t_L g157 ( .A(n_13), .Y(n_157) );
INVx1_ASAP7_75t_L g538 ( .A(n_14), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_15), .A2(n_147), .B(n_221), .C(n_223), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_16), .B(n_213), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_17), .B(n_472), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_18), .B(n_173), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_19), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_20), .A2(n_207), .B(n_208), .C(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_21), .B(n_213), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_22), .B(n_149), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_23), .A2(n_181), .B(n_223), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_24), .B(n_149), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_25), .Y(n_253) );
INVx1_ASAP7_75t_L g145 ( .A(n_26), .Y(n_145) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_27), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_28), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_29), .B(n_149), .Y(n_462) );
INVx1_ASAP7_75t_L g179 ( .A(n_30), .Y(n_179) );
INVx1_ASAP7_75t_L g483 ( .A(n_31), .Y(n_483) );
INVx2_ASAP7_75t_L g135 ( .A(n_32), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_33), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_34), .A2(n_207), .B(n_266), .C(n_268), .Y(n_265) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_35), .A2(n_88), .B1(n_449), .B2(n_729), .C1(n_732), .C2(n_733), .Y(n_448) );
INVxp67_ASAP7_75t_L g180 ( .A(n_36), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_37), .A2(n_141), .B(n_144), .C(n_152), .Y(n_140) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_38), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_39), .A2(n_137), .B(n_141), .C(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g482 ( .A(n_41), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_42), .A2(n_194), .B(n_195), .C(n_197), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_43), .B(n_149), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_44), .B(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_45), .A2(n_123), .B1(n_124), .B2(n_443), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_45), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_46), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_47), .Y(n_175) );
INVx1_ASAP7_75t_L g205 ( .A(n_48), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_49), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_50), .B(n_173), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_51), .A2(n_141), .B1(n_210), .B2(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_52), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_53), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g192 ( .A(n_54), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_55), .A2(n_194), .B(n_268), .C(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_56), .Y(n_531) );
INVx1_ASAP7_75t_L g490 ( .A(n_57), .Y(n_490) );
INVx1_ASAP7_75t_L g138 ( .A(n_58), .Y(n_138) );
INVx1_ASAP7_75t_L g156 ( .A(n_59), .Y(n_156) );
INVx1_ASAP7_75t_SL g267 ( .A(n_60), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_62), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g256 ( .A(n_63), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_64), .A2(n_268), .B(n_472), .C(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g474 ( .A(n_65), .Y(n_474) );
INVx1_ASAP7_75t_L g103 ( .A(n_66), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_67), .A2(n_173), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_68), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_69), .A2(n_173), .B(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_70), .Y(n_486) );
INVx1_ASAP7_75t_L g525 ( .A(n_71), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_72), .A2(n_172), .B(n_174), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_73), .Y(n_139) );
INVx1_ASAP7_75t_L g219 ( .A(n_74), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_75), .A2(n_137), .B(n_141), .C(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_76), .A2(n_100), .B1(n_111), .B2(n_736), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_77), .A2(n_173), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g222 ( .A(n_78), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_79), .B(n_146), .Y(n_507) );
INVx2_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
INVx1_ASAP7_75t_L g237 ( .A(n_81), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_82), .B(n_472), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_83), .A2(n_137), .B(n_141), .C(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g106 ( .A(n_84), .Y(n_106) );
OR2x2_ASAP7_75t_L g121 ( .A(n_84), .B(n_107), .Y(n_121) );
OR2x2_ASAP7_75t_L g728 ( .A(n_84), .B(n_108), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_85), .A2(n_141), .B(n_255), .C(n_258), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_86), .B(n_153), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_87), .Y(n_465) );
CKINVDCx14_ASAP7_75t_R g732 ( .A(n_88), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_89), .A2(n_137), .B(n_141), .C(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_90), .Y(n_520) );
INVx1_ASAP7_75t_L g470 ( .A(n_91), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_92), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_93), .B(n_146), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_94), .B(n_161), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_95), .B(n_161), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_96), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g209 ( .A(n_97), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_98), .A2(n_173), .B(n_469), .Y(n_468) );
CKINVDCx12_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g737 ( .A(n_101), .Y(n_737) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g733 ( .A(n_104), .Y(n_733) );
INVx3_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
NOR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g725 ( .A(n_106), .B(n_108), .Y(n_725) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_447), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g735 ( .A(n_115), .Y(n_735) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_444), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_121), .Y(n_446) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_125), .A2(n_450), .B1(n_723), .B2(n_726), .Y(n_449) );
INVx1_ASAP7_75t_SL g731 ( .A(n_125), .Y(n_731) );
OR5x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_337), .C(n_401), .D(n_417), .E(n_432), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_271), .C(n_298), .D(n_321), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_214), .B(n_225), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_SL g248 ( .A(n_130), .Y(n_248) );
AND2x4_ASAP7_75t_L g284 ( .A(n_130), .B(n_273), .Y(n_284) );
OR2x2_ASAP7_75t_L g294 ( .A(n_130), .B(n_250), .Y(n_294) );
OR2x2_ASAP7_75t_L g340 ( .A(n_130), .B(n_166), .Y(n_340) );
AND2x2_ASAP7_75t_L g354 ( .A(n_130), .B(n_249), .Y(n_354) );
AND2x2_ASAP7_75t_L g397 ( .A(n_130), .B(n_287), .Y(n_397) );
AND2x2_ASAP7_75t_L g404 ( .A(n_130), .B(n_261), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_130), .B(n_313), .Y(n_423) );
AND2x2_ASAP7_75t_L g441 ( .A(n_130), .B(n_283), .Y(n_441) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_158), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_140), .C(n_153), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_132), .A2(n_234), .B(n_235), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_132), .A2(n_253), .B(n_254), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_132), .A2(n_458), .B(n_459), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_132), .A2(n_183), .B1(n_480), .B2(n_484), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_132), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
AND2x4_ASAP7_75t_L g173 ( .A(n_133), .B(n_137), .Y(n_173) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g151 ( .A(n_134), .Y(n_151) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx1_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx1_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx3_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
INVx1_ASAP7_75t_L g472 ( .A(n_136), .Y(n_472) );
BUFx3_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx4_ASAP7_75t_SL g183 ( .A(n_137), .Y(n_183) );
INVx5_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_142), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_148), .C(n_150), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_146), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_146), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_147), .B(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_147), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_147), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx4_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_151), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_153), .A2(n_190), .B(n_199), .Y(n_189) );
INVx1_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_153), .A2(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_154), .B(n_155), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx3_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_160), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_160), .A2(n_252), .B(n_259), .Y(n_251) );
NOR2xp33_ASAP7_75t_SL g509 ( .A(n_160), .B(n_510), .Y(n_509) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_161), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g169 ( .A(n_162), .Y(n_169) );
INVx1_ASAP7_75t_L g406 ( .A(n_163), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_188), .Y(n_163) );
AND2x2_ASAP7_75t_L g316 ( .A(n_164), .B(n_249), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_164), .B(n_336), .Y(n_335) );
AOI32xp33_ASAP7_75t_L g349 ( .A1(n_164), .A2(n_350), .A3(n_353), .B1(n_355), .B2(n_359), .Y(n_349) );
AND2x2_ASAP7_75t_L g419 ( .A(n_164), .B(n_313), .Y(n_419) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g283 ( .A(n_166), .B(n_250), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_166), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g325 ( .A(n_166), .B(n_272), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_166), .B(n_404), .Y(n_403) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_184), .Y(n_166) );
INVx1_ASAP7_75t_L g288 ( .A(n_167), .Y(n_288) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_167), .A2(n_524), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_SL g503 ( .A1(n_168), .A2(n_504), .B(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_169), .A2(n_457), .B(n_464), .Y(n_456) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_169), .A2(n_479), .B(n_485), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_169), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_171), .A2(n_185), .B(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_176), .A2(n_183), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_SL g204 ( .A1(n_176), .A2(n_183), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_SL g218 ( .A1(n_176), .A2(n_183), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_176), .A2(n_183), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_176), .A2(n_183), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_176), .A2(n_183), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_176), .A2(n_183), .B(n_535), .C(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_181), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_181), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_181), .B(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g239 ( .A(n_182), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_182), .A2(n_239), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_187), .B(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_187), .A2(n_512), .B(n_519), .Y(n_511) );
AND2x2_ASAP7_75t_L g290 ( .A(n_188), .B(n_229), .Y(n_290) );
AND2x2_ASAP7_75t_L g366 ( .A(n_188), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g438 ( .A(n_188), .Y(n_438) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_200), .Y(n_188) );
OR2x2_ASAP7_75t_L g228 ( .A(n_189), .B(n_201), .Y(n_228) );
AND2x2_ASAP7_75t_L g245 ( .A(n_189), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_189), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g297 ( .A(n_189), .Y(n_297) );
AND2x2_ASAP7_75t_L g324 ( .A(n_189), .B(n_201), .Y(n_324) );
BUFx3_ASAP7_75t_L g327 ( .A(n_189), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_189), .B(n_302), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_189), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx2_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
AND2x2_ASAP7_75t_L g296 ( .A(n_200), .B(n_276), .Y(n_296) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g307 ( .A(n_201), .B(n_216), .Y(n_307) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_201), .Y(n_320) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_202), .A2(n_217), .B(n_224), .Y(n_216) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_202), .A2(n_262), .B(n_270), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_207), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g463 ( .A(n_210), .Y(n_463) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_213), .A2(n_488), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_215), .B(n_327), .Y(n_377) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_SL g246 ( .A(n_216), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_216), .B(n_296), .C(n_297), .Y(n_295) );
OR2x2_ASAP7_75t_L g303 ( .A(n_216), .B(n_276), .Y(n_303) );
AND2x2_ASAP7_75t_L g323 ( .A(n_216), .B(n_276), .Y(n_323) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_231), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_244), .B(n_247), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AND2x2_ASAP7_75t_L g442 ( .A(n_227), .B(n_367), .Y(n_442) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_228), .A2(n_340), .B1(n_382), .B2(n_384), .Y(n_381) );
OR2x2_ASAP7_75t_L g388 ( .A(n_228), .B(n_303), .Y(n_388) );
OR2x2_ASAP7_75t_L g412 ( .A(n_228), .B(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_228), .B(n_332), .Y(n_425) );
AND2x2_ASAP7_75t_L g318 ( .A(n_229), .B(n_319), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_229), .A2(n_391), .B(n_406), .Y(n_405) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_229), .A2(n_316), .A3(n_427), .B1(n_429), .B2(n_430), .Y(n_426) );
OR2x2_ASAP7_75t_L g437 ( .A(n_229), .B(n_438), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g305 ( .A(n_230), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_230), .B(n_319), .Y(n_384) );
BUFx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx4_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
AND2x2_ASAP7_75t_L g342 ( .A(n_231), .B(n_307), .Y(n_342) );
AND3x2_ASAP7_75t_L g351 ( .A(n_231), .B(n_245), .C(n_352), .Y(n_351) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_242), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_232), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_232), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_232), .B(n_531), .Y(n_530) );
O2A1O1Ixp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .C(n_241), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_238), .A2(n_241), .B(n_256), .C(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_241), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_241), .A2(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g277 ( .A(n_246), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_246), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_246), .B(n_276), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g272 ( .A(n_248), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g312 ( .A(n_248), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_248), .B(n_261), .Y(n_330) );
AND2x2_ASAP7_75t_L g348 ( .A(n_248), .B(n_250), .Y(n_348) );
OR2x2_ASAP7_75t_L g362 ( .A(n_248), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g408 ( .A(n_248), .B(n_336), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_249), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
AND2x2_ASAP7_75t_L g309 ( .A(n_250), .B(n_287), .Y(n_309) );
OR2x2_ASAP7_75t_L g363 ( .A(n_250), .B(n_287), .Y(n_363) );
AND2x2_ASAP7_75t_L g416 ( .A(n_250), .B(n_273), .Y(n_416) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g314 ( .A(n_251), .Y(n_314) );
AND2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_261), .Y(n_336) );
INVx2_ASAP7_75t_L g273 ( .A(n_261), .Y(n_273) );
INVx1_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_269), .Y(n_517) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_279), .C(n_291), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_272), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g435 ( .A(n_272), .Y(n_435) );
AND2x2_ASAP7_75t_L g313 ( .A(n_273), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_276), .B(n_277), .Y(n_285) );
INVx1_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_276), .B(n_297), .Y(n_394) );
AND2x2_ASAP7_75t_L g410 ( .A(n_276), .B(n_324), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_277), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_285), .B1(n_286), .B2(n_289), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_282), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_283), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_SL g373 ( .A1(n_284), .A2(n_326), .B1(n_374), .B2(n_379), .C(n_381), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_284), .B(n_347), .Y(n_380) );
INVx1_ASAP7_75t_L g440 ( .A(n_286), .Y(n_440) );
BUFx3_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_293), .B(n_347), .Y(n_400) );
INVx1_ASAP7_75t_L g357 ( .A(n_294), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_294), .B(n_347), .Y(n_358) );
INVxp67_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
AND2x2_ASAP7_75t_L g319 ( .A(n_297), .B(n_320), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B(n_308), .C(n_310), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_SL g333 ( .A(n_301), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_302), .B(n_333), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_302), .B(n_324), .Y(n_375) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_305), .A2(n_311), .B1(n_315), .B2(n_317), .Y(n_310) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g371 ( .A(n_307), .B(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_309), .A2(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_313), .A2(n_322), .B1(n_325), .B2(n_326), .C(n_328), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_313), .B(n_347), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_313), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g429 ( .A(n_319), .Y(n_429) );
INVxp67_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx1_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g398 ( .A(n_323), .B(n_327), .Y(n_398) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_327), .B(n_342), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_335), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g341 ( .A(n_336), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_336), .B(n_368), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_336), .B(n_397), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_336), .B(n_347), .Y(n_436) );
NAND5xp2_ASAP7_75t_L g337 ( .A(n_338), .B(n_360), .C(n_373), .D(n_385), .E(n_386), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_343), .B2(n_345), .C(n_349), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g364 ( .A(n_344), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_347), .B(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_348), .A2(n_361), .B1(n_364), .B2(n_368), .Y(n_360) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OAI211xp5_ASAP7_75t_SL g355 ( .A1(n_351), .A2(n_356), .B(n_357), .C(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g383 ( .A(n_363), .Y(n_383) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_372), .B(n_421), .Y(n_431) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_391), .B2(n_395), .C1(n_398), .C2(n_399), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_414), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_437), .C(n_439), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_444), .B(n_448), .C(n_734), .Y(n_447) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g730 ( .A(n_450), .Y(n_730) );
OR4x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_612), .C(n_672), .D(n_699), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_560), .C(n_591), .D(n_608), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_495), .B(n_497), .C(n_540), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_476), .Y(n_453) );
INVx1_ASAP7_75t_L g602 ( .A(n_454), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_454), .A2(n_643), .B1(n_691), .B2(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_455), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g553 ( .A(n_455), .B(n_478), .Y(n_553) );
AND2x2_ASAP7_75t_L g595 ( .A(n_455), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_455), .B(n_496), .Y(n_607) );
INVx1_ASAP7_75t_L g647 ( .A(n_455), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_455), .B(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g575 ( .A(n_456), .B(n_478), .Y(n_575) );
INVx3_ASAP7_75t_L g579 ( .A(n_456), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_456), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g666 ( .A(n_466), .B(n_487), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_466), .B(n_579), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_466), .B(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g496 ( .A(n_467), .B(n_478), .Y(n_496) );
INVx1_ASAP7_75t_L g548 ( .A(n_467), .Y(n_548) );
BUFx2_ASAP7_75t_L g552 ( .A(n_467), .Y(n_552) );
AND2x2_ASAP7_75t_L g596 ( .A(n_467), .B(n_477), .Y(n_596) );
OR2x2_ASAP7_75t_L g635 ( .A(n_467), .B(n_477), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_467), .B(n_487), .Y(n_660) );
AND2x2_ASAP7_75t_L g719 ( .A(n_467), .B(n_549), .Y(n_719) );
INVx1_ASAP7_75t_L g694 ( .A(n_476), .Y(n_694) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_477), .B(n_487), .Y(n_580) );
AND2x2_ASAP7_75t_L g590 ( .A(n_477), .B(n_579), .Y(n_590) );
BUFx2_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_487), .Y(n_623) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_478), .Y(n_678) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_487), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g549 ( .A(n_487), .Y(n_549) );
BUFx2_ASAP7_75t_L g574 ( .A(n_487), .Y(n_574) );
INVx2_ASAP7_75t_L g593 ( .A(n_487), .Y(n_593) );
AND2x2_ASAP7_75t_L g655 ( .A(n_487), .B(n_579), .Y(n_655) );
AOI321xp33_ASAP7_75t_L g674 ( .A1(n_495), .A2(n_675), .A3(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_496), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_496), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g668 ( .A(n_496), .B(n_647), .Y(n_668) );
AND2x2_ASAP7_75t_L g701 ( .A(n_496), .B(n_593), .Y(n_701) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_521), .Y(n_498) );
OR2x2_ASAP7_75t_L g603 ( .A(n_499), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_511), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g555 ( .A(n_502), .Y(n_555) );
AND2x2_ASAP7_75t_L g565 ( .A(n_502), .B(n_523), .Y(n_565) );
AND2x2_ASAP7_75t_L g570 ( .A(n_502), .B(n_545), .Y(n_570) );
INVx1_ASAP7_75t_L g587 ( .A(n_502), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_502), .B(n_568), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_502), .B(n_544), .Y(n_611) );
OR2x2_ASAP7_75t_L g643 ( .A(n_502), .B(n_632), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_502), .B(n_556), .Y(n_682) );
AND2x2_ASAP7_75t_L g716 ( .A(n_502), .B(n_542), .Y(n_716) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
INVx1_ASAP7_75t_L g543 ( .A(n_511), .Y(n_543) );
INVx2_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
AND2x2_ASAP7_75t_L g598 ( .A(n_511), .B(n_569), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_511), .B(n_545), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g704 ( .A(n_522), .B(n_555), .Y(n_704) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
INVx2_ASAP7_75t_L g545 ( .A(n_523), .Y(n_545) );
AND2x2_ASAP7_75t_L g698 ( .A(n_523), .B(n_558), .Y(n_698) );
AND2x2_ASAP7_75t_L g544 ( .A(n_532), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g559 ( .A(n_532), .Y(n_559) );
INVx1_ASAP7_75t_L g569 ( .A(n_532), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B1(n_550), .B2(n_554), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_541), .A2(n_659), .B1(n_696), .B2(n_697), .Y(n_695) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g610 ( .A(n_543), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_544), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_545), .B(n_558), .Y(n_632) );
INVx1_ASAP7_75t_L g648 ( .A(n_545), .Y(n_648) );
AND2x2_ASAP7_75t_L g589 ( .A(n_547), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_SL g628 ( .A(n_547), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_547), .B(n_553), .Y(n_705) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g714 ( .A(n_550), .Y(n_714) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_551), .B(n_647), .Y(n_689) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_SL g594 ( .A(n_553), .Y(n_594) );
NAND2x1_ASAP7_75t_SL g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g615 ( .A(n_555), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_555), .B(n_559), .Y(n_622) );
AND2x2_ASAP7_75t_L g627 ( .A(n_555), .B(n_568), .Y(n_627) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_555), .Y(n_676) );
OAI311xp33_ASAP7_75t_L g699 ( .A1(n_556), .A2(n_700), .A3(n_702), .B1(n_703), .C1(n_713), .Y(n_699) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g712 ( .A(n_557), .B(n_585), .Y(n_712) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g568 ( .A(n_558), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g616 ( .A(n_558), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
INVx1_ASAP7_75t_L g564 ( .A(n_559), .Y(n_564) );
INVx1_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_559), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g617 ( .A(n_559), .Y(n_617) );
AOI221xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B1(n_571), .B2(n_576), .C(n_581), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx4_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
AND2x2_ASAP7_75t_L g679 ( .A(n_565), .B(n_598), .Y(n_679) );
AND2x2_ASAP7_75t_L g686 ( .A(n_565), .B(n_568), .Y(n_686) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_568), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g597 ( .A(n_570), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_573), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g722 ( .A(n_575), .B(n_666), .Y(n_722) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g707 ( .A(n_579), .B(n_635), .Y(n_707) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_580), .A2(n_673), .B(n_674), .C(n_687), .Y(n_672) );
AOI21xp33_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_586), .B(n_588), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g651 ( .A(n_585), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_586), .A2(n_681), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_680) );
AND2x2_ASAP7_75t_L g657 ( .A(n_587), .B(n_598), .Y(n_657) );
AND2x2_ASAP7_75t_L g710 ( .A(n_587), .B(n_605), .Y(n_710) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_590), .B(n_628), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_595), .B(n_597), .C(n_599), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g638 ( .A(n_593), .B(n_596), .Y(n_638) );
OR2x2_ASAP7_75t_L g681 ( .A(n_593), .B(n_635), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_594), .B(n_660), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_594), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g625 ( .A(n_595), .Y(n_625) );
INVx1_ASAP7_75t_L g691 ( .A(n_598), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_606), .B2(n_607), .Y(n_599) );
INVx1_ASAP7_75t_L g614 ( .A(n_600), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_601), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g677 ( .A(n_602), .B(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g663 ( .A(n_604), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_605), .B(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_665), .B1(n_667), .B2(n_669), .Y(n_664) );
INVx1_ASAP7_75t_L g673 ( .A(n_609), .Y(n_673) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g715 ( .A(n_610), .B(n_710), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_611), .A2(n_645), .B1(n_648), .B2(n_649), .C1(n_652), .C2(n_653), .Y(n_644) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_633), .C(n_644), .D(n_656), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_618), .B2(n_623), .C(n_624), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_616), .B(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g642 ( .A(n_617), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_618), .A2(n_688), .B1(n_690), .B2(n_692), .C(n_695), .Y(n_687) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_622), .B(n_631), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_623), .A2(n_685), .B(n_686), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_628), .B2(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_639), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g675 ( .A(n_646), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_647), .B(n_666), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_647), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_651), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g683 ( .A(n_655), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g703 ( .A1(n_666), .A2(n_704), .B1(n_705), .B2(n_706), .C1(n_708), .C2(n_711), .Y(n_703) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_670), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g702 ( .A(n_676), .Y(n_702) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp33_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_716), .B2(n_717), .C(n_720), .Y(n_713) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_723), .A2(n_728), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
endmodule