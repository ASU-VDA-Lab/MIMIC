module fake_jpeg_22117_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_48;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_7),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_SL g17 ( 
.A1(n_8),
.A2(n_15),
.B(n_12),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_12),
.C(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_23),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.C(n_2),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_16),
.C(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_16),
.C(n_10),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_39),
.B1(n_28),
.B2(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_11),
.B1(n_15),
.B2(n_22),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_15),
.B1(n_11),
.B2(n_4),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_24),
.B(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_39),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_38),
.C(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_48),
.A3(n_35),
.B1(n_37),
.B2(n_5),
.C1(n_4),
.C2(n_3),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_4),
.Y(n_52)
);


endmodule