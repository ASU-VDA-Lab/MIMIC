module fake_jpeg_28332_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_52),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_35),
.B(n_40),
.C(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_17),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_42),
.B1(n_43),
.B2(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_30),
.B1(n_33),
.B2(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_58),
.B1(n_34),
.B2(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_24),
.B1(n_20),
.B2(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_21),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_81),
.B1(n_53),
.B2(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_43),
.B1(n_36),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_78),
.B1(n_42),
.B2(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_31),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_36),
.B1(n_32),
.B2(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_82),
.B1(n_84),
.B2(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_63),
.B1(n_79),
.B2(n_73),
.Y(n_111)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_45),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_80),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_45),
.B(n_32),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_105),
.B(n_28),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_69),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_55),
.B1(n_56),
.B2(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_104),
.B1(n_78),
.B2(n_77),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_3),
.C(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_55),
.B1(n_56),
.B2(n_49),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_56),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

AOI22x1_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_97),
.B1(n_105),
.B2(n_99),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_116),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_123),
.B1(n_27),
.B2(n_6),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_65),
.C(n_74),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_131),
.C(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_18),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_66),
.B1(n_69),
.B2(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_91),
.B1(n_69),
.B2(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_4),
.B(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_98),
.C(n_101),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_25),
.B1(n_28),
.B2(n_18),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_133),
.A2(n_22),
.B(n_16),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_69),
.A3(n_18),
.B1(n_19),
.B2(n_110),
.C1(n_31),
.C2(n_27),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_123),
.A3(n_114),
.B1(n_133),
.B2(n_120),
.C1(n_118),
.C2(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_121),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_148),
.B(n_155),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_109),
.B(n_108),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_11),
.B(n_12),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_109),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_130),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_19),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_96),
.C(n_27),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_124),
.C(n_116),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_19),
.B(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_154),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_169),
.C(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_171),
.B1(n_172),
.B2(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_132),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_170),
.B(n_162),
.Y(n_180)
);

XNOR2x2_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_130),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_145),
.C(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_138),
.C(n_136),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_160),
.B1(n_168),
.B2(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_151),
.B1(n_154),
.B2(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_142),
.C(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_188),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_197),
.B1(n_175),
.B2(n_186),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_170),
.B(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_192),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_163),
.B(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_171),
.B(n_148),
.C(n_158),
.Y(n_195)
);

AOI21x1_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_185),
.B(n_184),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_176),
.C(n_174),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_141),
.B1(n_12),
.B2(n_13),
.Y(n_197)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_205),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_11),
.C(n_12),
.Y(n_204)
);

OR2x2_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_191),
.Y(n_205)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_203),
.B(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_11),
.B1(n_14),
.B2(n_199),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_216),
.B(n_209),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_208),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_211),
.B(n_207),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_219),
.B(n_212),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_210),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_220),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_221),
.B(n_14),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_14),
.Y(n_224)
);


endmodule