module fake_jpeg_2061_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx4f_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_2),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_20),
.B(n_22),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_10),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_7),
.B1(n_10),
.B2(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_32),
.B1(n_22),
.B2(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_16),
.B1(n_22),
.B2(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.C(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_16),
.A3(n_18),
.B1(n_21),
.B2(n_22),
.C1(n_31),
.C2(n_27),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_39),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_39),
.B1(n_34),
.B2(n_40),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_30),
.B(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_25),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_36),
.Y(n_45)
);

NOR2xp67_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_42),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_47),
.B(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_43),
.Y(n_55)
);


endmodule