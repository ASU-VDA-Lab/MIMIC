module fake_jpeg_14894_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_21),
.CON(n_43),
.SN(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_26),
.B(n_21),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_43),
.B(n_55),
.C(n_24),
.Y(n_77)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_37),
.B1(n_27),
.B2(n_25),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_21),
.B(n_26),
.C(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_35),
.B1(n_28),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_80),
.B1(n_76),
.B2(n_69),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_18),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_65),
.B(n_78),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_85),
.Y(n_91)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_34),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_75),
.B(n_16),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_31),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_24),
.B1(n_30),
.B2(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_18),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_57),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_97),
.B(n_108),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_24),
.B(n_47),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_113),
.B(n_75),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_44),
.B1(n_41),
.B2(n_33),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_95),
.B1(n_100),
.B2(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_20),
.B1(n_30),
.B2(n_32),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_104),
.Y(n_140)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_18),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_84),
.B1(n_75),
.B2(n_76),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_85),
.B1(n_86),
.B2(n_64),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_74),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_32),
.B(n_16),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_16),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_141),
.B(n_107),
.Y(n_163)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_72),
.B(n_33),
.C(n_81),
.D(n_79),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_103),
.A3(n_19),
.B1(n_22),
.B2(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_89),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_64),
.B1(n_33),
.B2(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_103),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_30),
.B1(n_20),
.B2(n_62),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_9),
.B1(n_15),
.B2(n_13),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_20),
.B1(n_62),
.B2(n_19),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_137),
.B1(n_88),
.B2(n_106),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_22),
.Y(n_136)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_62),
.B1(n_19),
.B2(n_22),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_91),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_0),
.B(n_1),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx4f_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_110),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_151),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_169),
.B(n_172),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_147),
.B(n_150),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_98),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_108),
.C(n_87),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_164),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_163),
.B1(n_165),
.B2(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_166),
.Y(n_185)
);

AO22x2_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_89),
.B1(n_108),
.B2(n_105),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_128),
.B1(n_119),
.B2(n_122),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_100),
.C(n_90),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_95),
.B1(n_89),
.B2(n_105),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_171),
.B1(n_127),
.B2(n_132),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_115),
.B(n_89),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_101),
.B1(n_99),
.B2(n_106),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_8),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_173),
.A2(n_174),
.B(n_141),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_198),
.B1(n_143),
.B2(n_173),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_190),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_197),
.B1(n_171),
.B2(n_167),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_201),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_193),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_134),
.B(n_133),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_143),
.Y(n_215)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_202),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_130),
.B1(n_142),
.B2(n_129),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_129),
.B1(n_137),
.B2(n_103),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_2),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_152),
.C(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_205),
.C(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_SL g242 ( 
.A(n_209),
.B(n_214),
.C(n_215),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_146),
.B(n_164),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_177),
.B(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_158),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_193),
.B1(n_197),
.B2(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_22),
.C(n_3),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_223),
.C(n_202),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_7),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_233),
.B1(n_243),
.B2(n_209),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_238),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_234),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.C(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_195),
.C(n_182),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_2),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_175),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_178),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_198),
.B1(n_184),
.B2(n_183),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_256),
.C(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_214),
.B1(n_203),
.B2(n_206),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_257),
.B1(n_251),
.B2(n_254),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_221),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_203),
.B(n_190),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_179),
.B(n_223),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_240),
.B1(n_234),
.B2(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_266),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_237),
.CI(n_255),
.CON(n_262),
.SN(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_248),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_226),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_227),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_270),
.A2(n_250),
.B1(n_256),
.B2(n_2),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_9),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_268),
.B1(n_264),
.B2(n_261),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_262),
.B1(n_264),
.B2(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_286),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_3),
.C(n_4),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_285),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_3),
.C(n_4),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_288),
.B(n_6),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_6),
.B(n_7),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_281),
.B1(n_272),
.B2(n_274),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_276),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_285),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_287),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_297),
.C(n_290),
.Y(n_298)
);

AOI321xp33_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.A3(n_289),
.B1(n_11),
.B2(n_12),
.C(n_10),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_6),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_10),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_11),
.Y(n_302)
);


endmodule