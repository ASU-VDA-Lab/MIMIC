module fake_ariane_526_n_318 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_318);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_318;

wire n_295;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_183;
wire n_299;
wire n_133;
wire n_205;
wire n_109;
wire n_245;
wire n_283;
wire n_187;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_189;
wire n_286;
wire n_117;
wire n_139;
wire n_130;
wire n_214;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_279;
wire n_207;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_115;
wire n_267;
wire n_291;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_227;
wire n_188;
wire n_129;
wire n_126;
wire n_282;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_276;
wire n_108;
wire n_303;
wire n_168;
wire n_206;
wire n_238;
wire n_136;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_221;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_287;
wire n_302;
wire n_284;
wire n_249;
wire n_123;
wire n_212;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_150;
wire n_113;
wire n_114;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_246;
wire n_159;
wire n_131;
wire n_263;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_185;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_258;
wire n_118;
wire n_121;
wire n_241;
wire n_191;
wire n_211;
wire n_251;
wire n_116;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_50),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_18),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_8),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_60),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_39),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_26),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_43),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_35),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_16),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_3),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_41),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_85),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_64),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_44),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_36),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_49),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_89),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_97),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_17),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_38),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_24),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_37),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_17),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_1),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_1),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_2),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_4),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_5),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_6),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_6),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_129),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_7),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_9),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_9),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_118),
.B(n_10),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_12),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_137),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_13),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_14),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_15),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_19),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_149),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_20),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_22),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_167),
.B1(n_158),
.B2(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_165),
.B1(n_166),
.B2(n_164),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_163),
.B1(n_162),
.B2(n_109),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_185),
.B1(n_191),
.B2(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_110),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_123),
.B1(n_124),
.B2(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

AO22x2_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_157),
.B1(n_156),
.B2(n_155),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_140),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_146),
.B1(n_144),
.B2(n_143),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_175),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_171),
.A2(n_148),
.B1(n_132),
.B2(n_33),
.Y(n_223)
);

AO22x2_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_169),
.B(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_187),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_198),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_222),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_218),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_177),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_208),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_201),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_204),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_243),
.Y(n_256)
);

OR2x6_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_231),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_205),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_176),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_252),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_251),
.B(n_252),
.Y(n_269)
);

BUFx2_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

BUFx2_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_261),
.B1(n_263),
.B2(n_259),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_270),
.B1(n_271),
.B2(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_272),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_245),
.B1(n_275),
.B2(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_181),
.B1(n_174),
.B2(n_190),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_42),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_48),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_53),
.B(n_54),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_62),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_290),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_285),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

OAI22x1_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_309)
);

AO22x2_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_312),
.B1(n_88),
.B2(n_90),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

AOI221xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.C(n_99),
.Y(n_317)
);

AOI211xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_100),
.B(n_101),
.C(n_103),
.Y(n_318)
);


endmodule