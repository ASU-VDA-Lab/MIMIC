module fake_jpeg_14464_n_593 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_593);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_593;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_61),
.B(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_19),
.A2(n_7),
.B(n_15),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_67),
.A2(n_46),
.B(n_21),
.C(n_41),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_7),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_73),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_84),
.B(n_93),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_85),
.Y(n_163)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_88),
.Y(n_126)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_7),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_100),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_85),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_16),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_6),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_13),
.Y(n_184)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_57),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_32),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_19),
.B(n_6),
.C(n_14),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_32),
.C(n_30),
.Y(n_174)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_124),
.B(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_48),
.B1(n_45),
.B2(n_54),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_132),
.A2(n_182),
.B1(n_105),
.B2(n_101),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_148),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_85),
.A2(n_29),
.B1(n_32),
.B2(n_48),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_86),
.B1(n_107),
.B2(n_110),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_18),
.B(n_47),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_158),
.B(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_161),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_88),
.A2(n_41),
.B(n_42),
.C(n_49),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_70),
.B(n_18),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_60),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_59),
.A2(n_47),
.B1(n_53),
.B2(n_46),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_43),
.B(n_92),
.C(n_82),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_112),
.A2(n_31),
.B1(n_53),
.B2(n_49),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_76),
.B(n_21),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_66),
.B(n_30),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_198),
.B(n_43),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_203),
.A2(n_214),
.B(n_224),
.Y(n_286)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_97),
.B1(n_31),
.B2(n_72),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_78),
.B1(n_63),
.B2(n_83),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_206),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_207),
.A2(n_212),
.B1(n_264),
.B2(n_189),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_38),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_208),
.B(n_216),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_140),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_209),
.B(n_226),
.Y(n_293)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_210),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_142),
.A2(n_116),
.B1(n_96),
.B2(n_74),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_148),
.B(n_108),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_38),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_136),
.A2(n_119),
.B1(n_42),
.B2(n_25),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_218),
.A2(n_240),
.B1(n_241),
.B2(n_262),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_219),
.A2(n_232),
.B1(n_211),
.B2(n_222),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_142),
.B(n_0),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_246),
.Y(n_295)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_140),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_250),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_154),
.Y(n_237)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_135),
.A2(n_43),
.B1(n_77),
.B2(n_98),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_127),
.A2(n_43),
.B1(n_57),
.B2(n_6),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_123),
.B(n_0),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_137),
.Y(n_247)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_249),
.B(n_258),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_158),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_253),
.Y(n_322)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_152),
.Y(n_252)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_150),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_143),
.Y(n_255)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_255),
.Y(n_309)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_256),
.Y(n_304)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_15),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_129),
.Y(n_259)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_133),
.Y(n_260)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_261),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_197),
.A2(n_15),
.B1(n_11),
.B2(n_9),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_155),
.B(n_1),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_268),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_169),
.A2(n_15),
.B1(n_11),
.B2(n_6),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_139),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_267),
.B1(n_271),
.B2(n_146),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_1),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_269),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_171),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_194),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_145),
.Y(n_317)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_139),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_178),
.B(n_2),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_164),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_181),
.B(n_5),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_5),
.Y(n_296)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_181),
.A3(n_185),
.B1(n_130),
.B2(n_175),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_276),
.B(n_294),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_278),
.A2(n_268),
.B1(n_234),
.B2(n_220),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_219),
.A2(n_131),
.B1(n_166),
.B2(n_189),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_288),
.A2(n_327),
.B1(n_328),
.B2(n_242),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_253),
.A2(n_131),
.B1(n_166),
.B2(n_176),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_303),
.B1(n_313),
.B2(n_329),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_228),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_296),
.B(n_263),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_299),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_191),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_224),
.A2(n_159),
.B1(n_146),
.B2(n_176),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_310),
.A2(n_221),
.B1(n_225),
.B2(n_238),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_215),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_317),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_239),
.A2(n_232),
.B1(n_252),
.B2(n_165),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_156),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_330),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_203),
.A2(n_145),
.A3(n_159),
.B1(n_165),
.B2(n_151),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_317),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_208),
.B(n_190),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_323),
.B(n_217),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_270),
.A2(n_190),
.B1(n_216),
.B2(n_239),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_237),
.A2(n_223),
.B1(n_227),
.B2(n_272),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_272),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_343),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_358),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_278),
.A2(n_202),
.B1(n_254),
.B2(n_247),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_243),
.B1(n_271),
.B2(n_256),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_342),
.B(n_355),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_293),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_258),
.B(n_214),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_344),
.A2(n_325),
.B(n_314),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_233),
.C(n_231),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_348),
.C(n_374),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_292),
.B(n_226),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_350),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_235),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_351),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_244),
.C(n_248),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_213),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_288),
.A2(n_265),
.B1(n_210),
.B2(n_204),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_368),
.B1(n_372),
.B2(n_376),
.Y(n_381)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_296),
.A2(n_236),
.B1(n_245),
.B2(n_259),
.Y(n_358)
);

OAI22x1_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_304),
.B1(n_311),
.B2(n_283),
.Y(n_382)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_360),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_315),
.A2(n_255),
.B1(n_257),
.B2(n_261),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_373),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_297),
.B1(n_327),
.B2(n_276),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_295),
.B(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_275),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_370),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_286),
.A2(n_297),
.B1(n_282),
.B2(n_285),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_298),
.B(n_299),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_298),
.A2(n_321),
.B1(n_285),
.B2(n_299),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_339),
.B(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_275),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_280),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_374),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_274),
.B1(n_305),
.B2(n_300),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_279),
.A2(n_274),
.B1(n_305),
.B2(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_280),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_277),
.B(n_326),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_362),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_289),
.A2(n_290),
.B1(n_304),
.B2(n_301),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_369),
.A2(n_301),
.B1(n_304),
.B2(n_289),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_377),
.A2(n_384),
.B1(n_397),
.B2(n_400),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_368),
.A2(n_332),
.B(n_363),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_394),
.B(n_402),
.Y(n_433)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_387),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_332),
.A2(n_290),
.B1(n_319),
.B2(n_309),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_366),
.A2(n_311),
.B1(n_320),
.B2(n_324),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_386),
.A2(n_403),
.B(n_409),
.Y(n_441)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_364),
.A3(n_337),
.B1(n_346),
.B2(n_342),
.C1(n_333),
.C2(n_350),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_390),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_336),
.A2(n_325),
.B(n_308),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_SL g396 ( 
.A1(n_341),
.A2(n_316),
.B(n_287),
.C(n_308),
.Y(n_396)
);

AO21x1_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_381),
.B(n_399),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_355),
.A2(n_287),
.B1(n_316),
.B2(n_334),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_334),
.A2(n_351),
.B1(n_347),
.B2(n_343),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_344),
.A2(n_372),
.B(n_335),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_405),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_375),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_354),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_356),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_335),
.A2(n_345),
.B(n_373),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_409),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_361),
.A2(n_358),
.B1(n_349),
.B2(n_340),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_413),
.A2(n_399),
.B1(n_410),
.B2(n_408),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_360),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_414),
.B(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_365),
.C(n_370),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_426),
.C(n_430),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_378),
.A2(n_352),
.B(n_353),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_418),
.A2(n_435),
.B(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_384),
.A2(n_354),
.B1(n_371),
.B2(n_397),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_424),
.A2(n_446),
.B(n_391),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_425),
.B(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_400),
.C(n_403),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_383),
.B(n_405),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_383),
.Y(n_431)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_410),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_436),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_402),
.B(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_437),
.A2(n_449),
.B(n_422),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_390),
.A2(n_395),
.B(n_393),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_380),
.B(n_389),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_440),
.A2(n_396),
.B1(n_390),
.B2(n_382),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_385),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_437),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_444),
.A2(n_448),
.B1(n_391),
.B2(n_396),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_388),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_445),
.A2(n_403),
.B(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_390),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_386),
.B1(n_403),
.B2(n_381),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_394),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_450),
.B(n_464),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_377),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_458),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_426),
.B(n_387),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_454),
.B(n_423),
.Y(n_499)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_415),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_456),
.B(n_462),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_457),
.A2(n_461),
.B1(n_447),
.B2(n_446),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_390),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_418),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_433),
.A2(n_382),
.B(n_392),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_466),
.A2(n_471),
.B1(n_478),
.B2(n_440),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_427),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_472),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_391),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_475),
.C(n_433),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_396),
.B1(n_391),
.B2(n_406),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_474),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_406),
.C(n_411),
.Y(n_475)
);

XOR2x2_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_438),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_441),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_396),
.B1(n_411),
.B2(n_442),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_432),
.Y(n_518)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_473),
.Y(n_484)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

OA22x2_ASAP7_75t_L g527 ( 
.A1(n_485),
.A2(n_495),
.B1(n_498),
.B2(n_423),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_487),
.B(n_499),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_441),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_496),
.Y(n_514)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_489),
.Y(n_521)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_490),
.Y(n_516)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_491),
.Y(n_508)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_492),
.A2(n_493),
.B1(n_445),
.B2(n_468),
.Y(n_522)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_436),
.C(n_443),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_505),
.C(n_475),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_464),
.A2(n_423),
.B(n_447),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_497),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_416),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_460),
.A2(n_423),
.B(n_447),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_422),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_501),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_428),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_488),
.Y(n_515)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_504),
.B(n_482),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_432),
.C(n_428),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g506 ( 
.A(n_505),
.B(n_460),
.CI(n_476),
.CON(n_506),
.SN(n_506)
);

MAJIxp5_ASAP7_75t_SL g538 ( 
.A(n_506),
.B(n_499),
.C(n_487),
.Y(n_538)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_509),
.B(n_515),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_463),
.C(n_450),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_518),
.C(n_520),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_480),
.B(n_479),
.Y(n_519)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_519),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_478),
.Y(n_520)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_522),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_483),
.A2(n_423),
.B1(n_440),
.B2(n_466),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_523),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_468),
.C(n_461),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_525),
.C(n_481),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_486),
.B(n_471),
.C(n_477),
.Y(n_525)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_513),
.A2(n_500),
.B(n_485),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_528),
.A2(n_535),
.B(n_538),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_501),
.Y(n_530)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_492),
.Y(n_533)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_537),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_511),
.A2(n_500),
.B(n_493),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_525),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_459),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_503),
.C(n_491),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_539),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_517),
.A2(n_423),
.B1(n_502),
.B2(n_421),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_540),
.A2(n_544),
.B1(n_500),
.B2(n_511),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_508),
.A2(n_423),
.B1(n_451),
.B2(n_477),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_515),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_547),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_514),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_541),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_551),
.B(n_553),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_552),
.A2(n_532),
.B1(n_531),
.B2(n_533),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_518),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_555),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_520),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_531),
.A2(n_508),
.B1(n_524),
.B2(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_556),
.B(n_558),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_535),
.A2(n_527),
.B(n_506),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_514),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_559),
.B(n_545),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_542),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_564),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_559),
.B(n_530),
.Y(n_565)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_565),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_528),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_546),
.C(n_555),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_567),
.B(n_568),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_547),
.B(n_539),
.C(n_548),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_549),
.B(n_534),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_568),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_572),
.B(n_575),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_558),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_577),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_569),
.A2(n_532),
.B(n_557),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_574),
.A2(n_560),
.B(n_537),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_527),
.C(n_538),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_578),
.B(n_561),
.Y(n_581)
);

AOI21x1_ASAP7_75t_SL g586 ( 
.A1(n_581),
.A2(n_584),
.B(n_573),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_570),
.C(n_566),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_583),
.A2(n_579),
.B(n_577),
.Y(n_585)
);

AO21x1_ASAP7_75t_L g589 ( 
.A1(n_585),
.A2(n_587),
.B(n_526),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_586),
.A2(n_582),
.B(n_527),
.Y(n_588)
);

AO21x1_ASAP7_75t_L g587 ( 
.A1(n_580),
.A2(n_575),
.B(n_506),
.Y(n_587)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_588),
.A2(n_589),
.B(n_526),
.Y(n_590)
);

O2A1O1Ixp33_ASAP7_75t_SL g591 ( 
.A1(n_590),
.A2(n_419),
.B(n_420),
.C(n_429),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_434),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_396),
.Y(n_593)
);


endmodule