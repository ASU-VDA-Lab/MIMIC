module fake_jpeg_29246_n_534 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_60),
.Y(n_107)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx2_ASAP7_75t_SL g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_101),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_91),
.Y(n_147)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_28),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_17),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_89),
.Y(n_145)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_17),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_103),
.B1(n_49),
.B2(n_38),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_40),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_21),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_24),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_38),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_37),
.B(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_48),
.B1(n_21),
.B2(n_27),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_140),
.B1(n_151),
.B2(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_152),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_48),
.B1(n_25),
.B2(n_24),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_138),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_49),
.B1(n_42),
.B2(n_38),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_74),
.B(n_25),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_58),
.A2(n_60),
.B1(n_59),
.B2(n_62),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_66),
.B(n_19),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_20),
.B1(n_37),
.B2(n_46),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_56),
.B(n_38),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_82),
.B(n_50),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_64),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_93),
.B(n_50),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_166),
.A2(n_182),
.B1(n_133),
.B2(n_110),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_132),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_171),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_46),
.B(n_47),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_170),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_22),
.B1(n_29),
.B2(n_39),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_197),
.Y(n_224)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_50),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_180),
.Y(n_228)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_29),
.Y(n_180)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx6p67_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_201),
.B1(n_211),
.B2(n_107),
.Y(n_234)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_103),
.B1(n_97),
.B2(n_96),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_139),
.A2(n_38),
.B1(n_47),
.B2(n_29),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_203),
.B1(n_205),
.B2(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_199),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_126),
.A2(n_22),
.B1(n_47),
.B2(n_39),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_40),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_202),
.B(n_206),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_149),
.A2(n_39),
.B1(n_22),
.B2(n_98),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_208),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_124),
.A2(n_99),
.B1(n_100),
.B2(n_40),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_116),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_107),
.A2(n_40),
.B(n_1),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_213),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_210),
.Y(n_255)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_140),
.A2(n_40),
.B1(n_41),
.B2(n_2),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_124),
.A2(n_40),
.B1(n_41),
.B2(n_2),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_142),
.C(n_130),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_217),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_113),
.B1(n_143),
.B2(n_156),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_221),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_220),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_155),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_122),
.B(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_128),
.A2(n_41),
.B1(n_9),
.B2(n_10),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_167),
.B(n_131),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_253),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_215),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_150),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_245),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_251),
.B1(n_256),
.B2(n_259),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_173),
.A2(n_125),
.B1(n_162),
.B2(n_157),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_244),
.A2(n_252),
.B1(n_218),
.B2(n_220),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_125),
.B(n_164),
.C(n_142),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_133),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_249),
.B(n_262),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_250),
.A2(n_177),
.B1(n_219),
.B2(n_169),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_173),
.A2(n_110),
.B1(n_106),
.B2(n_156),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_106),
.B1(n_155),
.B2(n_41),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_196),
.B(n_7),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_170),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_254),
.A2(n_270),
.B1(n_206),
.B2(n_168),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_16),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_12),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_262),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_215),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_304),
.B1(n_235),
.B2(n_257),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_202),
.B1(n_181),
.B2(n_215),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_277),
.A2(n_293),
.B1(n_303),
.B2(n_305),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_175),
.A3(n_171),
.B1(n_194),
.B2(n_192),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_279),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

NAND2x1_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_207),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_280),
.A2(n_235),
.B(n_258),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_285),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_267),
.C(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_236),
.C(n_229),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_256),
.B1(n_259),
.B2(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

BUFx24_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_172),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_183),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_297),
.B(n_307),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_186),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_299),
.A2(n_302),
.B1(n_257),
.B2(n_246),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_265),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_300),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_301),
.B(n_239),
.Y(n_333)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_179),
.B1(n_213),
.B2(n_210),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_234),
.A2(n_209),
.B1(n_189),
.B2(n_184),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_242),
.B1(n_268),
.B2(n_261),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_214),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_193),
.Y(n_339)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_231),
.B(n_188),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_200),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_309),
.B(n_311),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_242),
.B(n_254),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_273),
.B(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_335),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_273),
.A2(n_242),
.B(n_268),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_344),
.B(n_306),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_345),
.C(n_237),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_281),
.A2(n_227),
.B(n_257),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_319),
.A2(n_339),
.B(n_281),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_229),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_332),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_321),
.A2(n_323),
.B1(n_348),
.B2(n_233),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_301),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_333),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_269),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_291),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_334),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_258),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_341),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_233),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_343),
.B(n_260),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_306),
.A2(n_239),
.B(n_230),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_230),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_276),
.A2(n_260),
.B1(n_185),
.B2(n_233),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_349),
.A2(n_338),
.B(n_346),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_341),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_376),
.Y(n_394)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_272),
.B(n_297),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_352),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_354),
.B(n_370),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_319),
.A2(n_300),
.B(n_276),
.Y(n_354)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx3_ASAP7_75t_SL g395 ( 
.A(n_356),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_316),
.A2(n_304),
.B1(n_288),
.B2(n_271),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_357),
.A2(n_359),
.B1(n_362),
.B2(n_321),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_303),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_358),
.B(n_363),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_275),
.B1(n_279),
.B2(n_272),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_SL g360 ( 
.A1(n_314),
.A2(n_280),
.B(n_275),
.C(n_278),
.Y(n_360)
);

AOI21x1_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_371),
.B(n_373),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_225),
.Y(n_361)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_325),
.A2(n_280),
.B1(n_307),
.B2(n_311),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_342),
.A2(n_274),
.B1(n_294),
.B2(n_292),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_225),
.Y(n_367)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_322),
.B1(n_334),
.B2(n_313),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_325),
.B(n_237),
.Y(n_369)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_289),
.Y(n_370)
);

NAND2x1_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_284),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_339),
.A2(n_283),
.B(n_302),
.Y(n_373)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_344),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_323),
.A2(n_290),
.B1(n_237),
.B2(n_220),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_378),
.Y(n_412)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_290),
.C(n_14),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_320),
.C(n_317),
.Y(n_388)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_380),
.Y(n_409)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_381),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_413),
.B1(n_357),
.B2(n_371),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_345),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_388),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_401),
.B1(n_406),
.B2(n_381),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_333),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_393),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_391),
.B(n_354),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_312),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_332),
.C(n_336),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_397),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_312),
.C(n_339),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_313),
.C(n_337),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_399),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_362),
.C(n_349),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_377),
.A2(n_337),
.B1(n_348),
.B2(n_329),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_404),
.A2(n_382),
.B(n_363),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_346),
.B1(n_329),
.B2(n_324),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_370),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_379),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_355),
.B(n_324),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_366),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_359),
.A2(n_326),
.B1(n_343),
.B2(n_290),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_405),
.B(n_366),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_414),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_412),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_406),
.Y(n_417)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_331),
.Y(n_462)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_395),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_372),
.Y(n_422)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_370),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_426),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_402),
.B(n_382),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_427),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_355),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_428),
.B(n_429),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_383),
.A2(n_353),
.B(n_371),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_430),
.A2(n_440),
.B1(n_401),
.B2(n_397),
.Y(n_456)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_431),
.A2(n_434),
.B1(n_437),
.B2(n_438),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_439),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_409),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_435),
.A2(n_436),
.B1(n_413),
.B2(n_384),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_365),
.B1(n_360),
.B2(n_373),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_380),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_390),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_411),
.A2(n_365),
.B1(n_360),
.B2(n_356),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_393),
.C(n_388),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_444),
.C(n_448),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_442),
.A2(n_445),
.B1(n_449),
.B2(n_458),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_391),
.C(n_399),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_435),
.A2(n_411),
.B1(n_385),
.B2(n_360),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_398),
.C(n_396),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_436),
.A2(n_411),
.B1(n_385),
.B2(n_360),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_456),
.A2(n_459),
.B1(n_437),
.B2(n_432),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_383),
.B1(n_400),
.B2(n_386),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_430),
.A2(n_326),
.B1(n_389),
.B2(n_331),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_331),
.C(n_14),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_461),
.B(n_434),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_429),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_471),
.Y(n_494)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_461),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_466),
.B(n_468),
.Y(n_483)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_414),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_473),
.Y(n_491)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_455),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_479),
.B1(n_455),
.B2(n_449),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_442),
.A2(n_440),
.B1(n_415),
.B2(n_426),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_L g482 ( 
.A1(n_474),
.A2(n_427),
.B1(n_424),
.B2(n_428),
.C(n_418),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_425),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_477),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_431),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_452),
.B(n_437),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_416),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_416),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_460),
.C(n_441),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_476),
.A2(n_463),
.B1(n_453),
.B2(n_445),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_481),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_484),
.B(n_486),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_487),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_469),
.A2(n_452),
.B1(n_451),
.B2(n_458),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_448),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_488),
.A2(n_422),
.B(n_421),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_493),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_465),
.A2(n_457),
.B1(n_419),
.B2(n_425),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_492),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_471),
.A2(n_438),
.B1(n_457),
.B2(n_439),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_460),
.C(n_462),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_495),
.B(n_477),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_465),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_502),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_498),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_472),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_505),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_478),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_473),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_504),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_506),
.A2(n_485),
.B1(n_481),
.B2(n_489),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_447),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_493),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_515),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_483),
.Y(n_514)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_490),
.C(n_487),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_517),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_507),
.A2(n_420),
.B1(n_14),
.B2(n_15),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_519),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_512),
.A2(n_507),
.B(n_500),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_522),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_503),
.C(n_502),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_521),
.A2(n_511),
.B(n_516),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_511),
.B(n_510),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_528),
.C(n_524),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_523),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_518),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_501),
.B(n_519),
.Y(n_532)
);

AOI211xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_504),
.B(n_13),
.C(n_15),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_13),
.B1(n_15),
.B2(n_366),
.Y(n_534)
);


endmodule