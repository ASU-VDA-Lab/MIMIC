module fake_jpeg_13971_n_526 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_526);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_23),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_94),
.Y(n_130)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_18),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_63),
.B(n_89),
.Y(n_141)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx2_ASAP7_75t_SL g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g157 ( 
.A(n_75),
.Y(n_157)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_0),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_36),
.B(n_0),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_39),
.Y(n_132)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_28),
.B(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_44),
.B1(n_42),
.B2(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_105),
.A2(n_121),
.B1(n_136),
.B2(n_133),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_50),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_22),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_44),
.B1(n_42),
.B2(n_47),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_110),
.A2(n_87),
.B(n_83),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_50),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_117),
.B(n_134),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_59),
.A2(n_42),
.B1(n_44),
.B2(n_25),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_37),
.B1(n_33),
.B2(n_40),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_129),
.A2(n_138),
.B1(n_147),
.B2(n_160),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_40),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_48),
.B1(n_25),
.B2(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_137),
.B(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_62),
.A2(n_48),
.B1(n_43),
.B2(n_31),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_47),
.B1(n_39),
.B2(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_47),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_68),
.A2(n_47),
.B1(n_39),
.B2(n_22),
.Y(n_160)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_168),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_160),
.B1(n_93),
.B2(n_75),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_172),
.A2(n_183),
.B(n_200),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_174),
.B(n_192),
.Y(n_247)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_175),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_1),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_122),
.A2(n_67),
.B1(n_52),
.B2(n_72),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_197),
.Y(n_235)
);

AO22x2_ASAP7_75t_SL g183 ( 
.A1(n_105),
.A2(n_90),
.B1(n_99),
.B2(n_91),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_143),
.B1(n_139),
.B2(n_106),
.Y(n_248)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_190),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_122),
.A2(n_78),
.B1(n_74),
.B2(n_69),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_47),
.B1(n_39),
.B2(n_22),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_189),
.Y(n_251)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_194),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_199),
.Y(n_227)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_195),
.A2(n_202),
.B(n_14),
.Y(n_268)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_121),
.A2(n_80),
.B1(n_71),
.B2(n_39),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_183),
.B1(n_195),
.B2(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_203),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_22),
.B(n_3),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_136),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_204),
.A2(n_209),
.B1(n_211),
.B2(n_6),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_205),
.A2(n_206),
.B1(n_218),
.B2(n_219),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_207),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_212),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_17),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_115),
.C(n_151),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_145),
.A2(n_125),
.B1(n_112),
.B2(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_2),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_217),
.Y(n_256)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_108),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_171),
.B(n_118),
.CI(n_157),
.CON(n_223),
.SN(n_223)
);

MAJIxp5_ASAP7_75t_SL g285 ( 
.A(n_223),
.B(n_207),
.C(n_208),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_232),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_250),
.B1(n_255),
.B2(n_262),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_198),
.B(n_113),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_151),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_240),
.C(n_252),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_236),
.B(n_248),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_193),
.B(n_139),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_237),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_152),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_108),
.B(n_103),
.C(n_7),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_249),
.A2(n_223),
.B(n_266),
.C(n_261),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_106),
.B1(n_6),
.B2(n_7),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_2),
.C(n_6),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_172),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_258),
.A2(n_270),
.B1(n_238),
.B2(n_254),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_8),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_202),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_11),
.C(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_271),
.C(n_189),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_168),
.B1(n_197),
.B2(n_170),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_11),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_266),
.B(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_188),
.B(n_13),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_162),
.B(n_176),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_16),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_274),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_169),
.B1(n_219),
.B2(n_196),
.Y(n_275)
);

OAI22x1_ASAP7_75t_L g319 ( 
.A1(n_275),
.A2(n_295),
.B1(n_269),
.B2(n_238),
.Y(n_319)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_277),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_283),
.B1(n_288),
.B2(n_290),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_194),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_289),
.C(n_292),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_175),
.B(n_176),
.C(n_220),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_310),
.B(n_313),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_201),
.B1(n_203),
.B2(n_217),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_285),
.A2(n_293),
.B(n_300),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_286),
.B(n_253),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_190),
.B1(n_191),
.B2(n_206),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_226),
.B(n_205),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_271),
.B1(n_262),
.B2(n_236),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_165),
.B1(n_177),
.B2(n_16),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_309),
.B1(n_317),
.B2(n_260),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_234),
.B(n_16),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_247),
.A2(n_16),
.B(n_17),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_221),
.B(n_17),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_297),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_264),
.A2(n_17),
.B1(n_235),
.B2(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_240),
.B(n_227),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_227),
.B(n_225),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_302),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_223),
.A2(n_249),
.B1(n_224),
.B2(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_245),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_237),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_318),
.C(n_269),
.Y(n_347)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g333 ( 
.A1(n_306),
.A2(n_287),
.B(n_300),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_222),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_307),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_258),
.A2(n_248),
.B1(n_267),
.B2(n_241),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_256),
.A2(n_229),
.B(n_241),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_244),
.A2(n_254),
.B(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_248),
.B(n_257),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_316),
.A2(n_308),
.B(n_304),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_252),
.B(n_246),
.C(n_259),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_289),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_335),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_323),
.A2(n_340),
.B1(n_349),
.B2(n_352),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_287),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_338),
.C(n_341),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_257),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_259),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_273),
.A2(n_248),
.B1(n_264),
.B2(n_269),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_231),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_231),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_273),
.A2(n_290),
.B1(n_309),
.B2(n_283),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_274),
.A2(n_281),
.B(n_316),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_351),
.A2(n_357),
.B(n_272),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_296),
.B1(n_279),
.B2(n_288),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_318),
.C(n_286),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_328),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_356),
.A2(n_285),
.B(n_308),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_310),
.B(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_361),
.A2(n_371),
.B(n_375),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_313),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_362),
.B(n_384),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_351),
.A2(n_291),
.B1(n_298),
.B2(n_301),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_363),
.A2(n_365),
.B1(n_385),
.B2(n_388),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_359),
.A2(n_306),
.B1(n_276),
.B2(n_305),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_278),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_366),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_370),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_377),
.C(n_376),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_336),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_353),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_374),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_346),
.Y(n_374)
);

FAx1_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_357),
.CI(n_337),
.CON(n_375),
.SN(n_375)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_334),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_382),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_325),
.B(n_330),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_359),
.A2(n_337),
.B(n_354),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_389),
.B(n_326),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_327),
.B(n_332),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_349),
.A2(n_329),
.B1(n_325),
.B2(n_330),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_334),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_340),
.B1(n_344),
.B2(n_322),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_354),
.A2(n_347),
.B(n_319),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_390),
.Y(n_398)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_320),
.B(n_358),
.Y(n_392)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_345),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_342),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_343),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_394),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_373),
.A2(n_355),
.B1(n_338),
.B2(n_326),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_395),
.A2(n_409),
.B1(n_360),
.B2(n_364),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_341),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_414),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_405),
.C(n_382),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_403),
.A2(n_412),
.B(n_375),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_331),
.C(n_342),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_373),
.A2(n_331),
.B1(n_350),
.B2(n_321),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_321),
.B(n_361),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_392),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_381),
.B1(n_374),
.B2(n_370),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_420),
.B1(n_410),
.B2(n_423),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_417),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_390),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_378),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_388),
.A2(n_385),
.B1(n_363),
.B2(n_368),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_420),
.A2(n_423),
.B1(n_389),
.B2(n_383),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_379),
.B(n_387),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_422),
.B(n_375),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_387),
.B1(n_379),
.B2(n_375),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_425),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_428),
.B(n_439),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_431),
.A2(n_432),
.B(n_448),
.Y(n_456)
);

FAx1_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_386),
.CI(n_394),
.CON(n_432),
.SN(n_432)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_427),
.Y(n_451)
);

XOR2x2_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_440),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_367),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_444),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_409),
.A2(n_391),
.B1(n_364),
.B2(n_360),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_437),
.B(n_442),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_414),
.B(n_380),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_395),
.B(n_372),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_404),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_403),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_404),
.Y(n_445)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

OAI31xp33_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_406),
.A3(n_424),
.B(n_417),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_410),
.A2(n_402),
.B1(n_399),
.B2(n_398),
.Y(n_449)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_449),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_460),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_405),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_458),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_424),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_413),
.C(n_421),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_413),
.C(n_421),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_470),
.Y(n_483)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_466),
.Y(n_471)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_422),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_428),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_435),
.C(n_431),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_461),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_474),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_425),
.C(n_434),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_479),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_434),
.C(n_441),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_486),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_443),
.Y(n_481)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_453),
.B(n_447),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_464),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_415),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_485),
.A2(n_398),
.B1(n_443),
.B2(n_399),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_426),
.C(n_437),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_489),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_463),
.B1(n_467),
.B2(n_454),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_450),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_486),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_465),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_498),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_485),
.A2(n_397),
.B1(n_470),
.B2(n_402),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_456),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_493),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_496),
.B(n_472),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_502),
.B(n_507),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_474),
.C(n_484),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_506),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_487),
.A2(n_456),
.B(n_432),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_504),
.A2(n_448),
.B(n_494),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_471),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_418),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_491),
.B(n_499),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_500),
.B(n_505),
.Y(n_516)
);

AOI21x1_ASAP7_75t_SL g518 ( 
.A1(n_511),
.A2(n_512),
.B(n_514),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_490),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_516),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_515),
.A2(n_505),
.B(n_501),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_517),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_432),
.B(n_493),
.Y(n_519)
);

O2A1O1Ixp33_ASAP7_75t_SL g522 ( 
.A1(n_521),
.A2(n_518),
.B(n_519),
.C(n_513),
.Y(n_522)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_520),
.B(n_401),
.C(n_407),
.D(n_479),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_407),
.B(n_401),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_464),
.B1(n_482),
.B2(n_469),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_475),
.B(n_453),
.Y(n_526)
);


endmodule