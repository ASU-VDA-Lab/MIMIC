module fake_jpeg_31920_n_364 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_364);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_364;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_0),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_63),
.B(n_31),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_57),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_30),
.B1(n_23),
.B2(n_34),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_75),
.B1(n_80),
.B2(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_30),
.B1(n_23),
.B2(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_81),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_79),
.B1(n_42),
.B2(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_33),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_35),
.B(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_91),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_99),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_131),
.B(n_37),
.C(n_91),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_128),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_105),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_112),
.Y(n_157)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_117),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_125),
.B1(n_20),
.B2(n_25),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_71),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_123),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_37),
.B(n_22),
.C(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_130),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_37),
.B(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_63),
.B(n_67),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_35),
.B1(n_20),
.B2(n_22),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_57),
.C(n_56),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_37),
.C(n_59),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_27),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_75),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_25),
.B1(n_20),
.B2(n_37),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_60),
.B1(n_88),
.B2(n_68),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_137),
.B1(n_147),
.B2(n_149),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_110),
.B(n_116),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_128),
.B1(n_101),
.B2(n_126),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_100),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_155),
.B1(n_134),
.B2(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_59),
.C(n_68),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_153),
.C(n_110),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_53),
.B1(n_66),
.B2(n_56),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_46),
.B1(n_62),
.B2(n_90),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_46),
.C(n_62),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_125),
.B1(n_103),
.B2(n_106),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_83),
.B(n_92),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_114),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_104),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_166),
.B(n_174),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_142),
.B1(n_94),
.B2(n_159),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_135),
.B1(n_152),
.B2(n_144),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_178),
.Y(n_204)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_113),
.B1(n_112),
.B2(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_93),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_185),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_182),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_184),
.B(n_191),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_93),
.B(n_129),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_124),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_147),
.B1(n_149),
.B2(n_160),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_14),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_133),
.A3(n_119),
.B1(n_15),
.B2(n_14),
.C1(n_7),
.C2(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_107),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_115),
.B(n_116),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_119),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_140),
.B(n_90),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_162),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_139),
.C(n_153),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_180),
.C(n_197),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_212),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_191),
.B(n_185),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_135),
.B1(n_160),
.B2(n_146),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_216),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_152),
.B1(n_158),
.B2(n_138),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_230),
.B1(n_225),
.B2(n_216),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_226),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_162),
.B(n_154),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_172),
.B(n_164),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_177),
.Y(n_247)
);

OR2x6_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_159),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_174),
.B(n_169),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_154),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_176),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_158),
.B1(n_108),
.B2(n_102),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_246),
.B(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_236),
.B1(n_252),
.B2(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_230),
.B1(n_218),
.B2(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_249),
.C(n_208),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_173),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_245),
.B(n_215),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_170),
.B(n_169),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_189),
.C(n_181),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_255),
.Y(n_263)
);

OA21x2_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_169),
.B(n_138),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_258),
.B(n_229),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_82),
.B(n_83),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_8),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_12),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_214),
.B(n_17),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_267),
.C(n_279),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_208),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_249),
.C(n_238),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_213),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_213),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_240),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_209),
.B1(n_203),
.B2(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_247),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_232),
.A2(n_219),
.B1(n_209),
.B2(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_277),
.B1(n_258),
.B2(n_256),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_207),
.B1(n_221),
.B2(n_228),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_220),
.B1(n_206),
.B2(n_217),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_233),
.C(n_243),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_236),
.A2(n_217),
.B1(n_211),
.B2(n_212),
.Y(n_281)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_245),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_251),
.B1(n_234),
.B2(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_291),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_250),
.C(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_293),
.C(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_265),
.B(n_241),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_215),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_294),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_270),
.A2(n_254),
.B1(n_242),
.B2(n_248),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_298),
.B(n_300),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_255),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_301),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_260),
.A2(n_231),
.B(n_239),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_237),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_235),
.B(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_228),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_224),
.B(n_210),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_280),
.B(n_272),
.C(n_264),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_270),
.B1(n_279),
.B2(n_269),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_311),
.B1(n_283),
.B2(n_302),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_287),
.C(n_267),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_313),
.C(n_316),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_261),
.B(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_259),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_2),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_269),
.B1(n_272),
.B2(n_264),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_263),
.C(n_280),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_314),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_210),
.C(n_83),
.Y(n_316)
);

AO22x1_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_17),
.B1(n_82),
.B2(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_17),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_330),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_292),
.B1(n_295),
.B2(n_288),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_323),
.A2(n_325),
.B1(n_311),
.B2(n_304),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_285),
.B1(n_293),
.B2(n_299),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_294),
.B1(n_298),
.B2(n_12),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_326),
.A2(n_328),
.B1(n_2),
.B2(n_4),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_7),
.B(n_13),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_320),
.B(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_82),
.B1(n_4),
.B2(n_5),
.Y(n_328)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_306),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_316),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_17),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_317),
.B(n_314),
.Y(n_338)
);

OAI221xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_334),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_335),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

A2O1A1O1Ixp25_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_304),
.B(n_308),
.C(n_313),
.D(n_305),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_341),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_332),
.A2(n_2),
.B(n_4),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_344),
.B(n_345),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_2),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_337),
.A2(n_332),
.B(n_327),
.Y(n_348)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

NAND2x1_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_331),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_328),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_345),
.A2(n_322),
.B(n_323),
.C(n_329),
.Y(n_353)
);

O2A1O1Ixp33_ASAP7_75t_SL g357 ( 
.A1(n_353),
.A2(n_5),
.B(n_6),
.C(n_17),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_355),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_351),
.A2(n_339),
.B1(n_325),
.B2(n_6),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_17),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_359),
.C(n_349),
.Y(n_361)
);

OAI321xp33_ASAP7_75t_L g362 ( 
.A1(n_357),
.A2(n_350),
.A3(n_352),
.B1(n_353),
.B2(n_359),
.C(n_358),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_347),
.C(n_350),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_362),
.C(n_357),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_360),
.Y(n_364)
);


endmodule