module fake_ariane_1015_n_183 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_183);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_183;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_29),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

OR2x6_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_41),
.C(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_41),
.C(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_46),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_38),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_55),
.B(n_56),
.C(n_66),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_56),
.Y(n_93)
);

AO31x2_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_66),
.A3(n_53),
.B(n_52),
.Y(n_94)
);

AO31x2_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_70),
.A3(n_59),
.B(n_62),
.Y(n_95)
);

NOR2x1_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_68),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_65),
.B(n_85),
.C(n_88),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_63),
.B(n_70),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AOI21x1_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_68),
.B(n_32),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_86),
.B(n_74),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_99),
.B(n_100),
.C(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_86),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_81),
.B(n_68),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_96),
.B1(n_71),
.B2(n_60),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_99),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_111),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_113),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_113),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_111),
.B(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_123),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_111),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_84),
.B1(n_108),
.B2(n_128),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_79),
.C(n_97),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_129),
.B1(n_69),
.B2(n_124),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_124),
.Y(n_144)
);

OAI221xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_69),
.B1(n_72),
.B2(n_78),
.C(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_114),
.Y(n_146)
);

NAND4xp25_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_1),
.C(n_3),
.D(n_4),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_60),
.B1(n_78),
.B2(n_75),
.C(n_82),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_1),
.C(n_3),
.D(n_4),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_114),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_6),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_6),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_95),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2x1p5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_115),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_115),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_148),
.C(n_8),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_7),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_7),
.B(n_9),
.C(n_13),
.Y(n_163)
);

NAND3x1_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_9),
.C(n_13),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_103),
.B1(n_107),
.B2(n_102),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_161),
.C(n_162),
.Y(n_168)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_153),
.A3(n_158),
.B1(n_154),
.B2(n_82),
.C(n_102),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_154),
.B1(n_103),
.B2(n_75),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_159),
.B1(n_167),
.B2(n_103),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_101),
.B1(n_98),
.B2(n_95),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_95),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_75),
.B1(n_95),
.B2(n_94),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_95),
.B1(n_94),
.B2(n_23),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_177),
.B1(n_174),
.B2(n_94),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_19),
.B(n_22),
.C(n_24),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_94),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_178),
.B1(n_181),
.B2(n_179),
.Y(n_183)
);


endmodule