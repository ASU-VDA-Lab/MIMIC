module fake_jpeg_23836_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_56),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_26),
.CON(n_45),
.SN(n_45)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_36),
.B1(n_15),
.B2(n_17),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_0),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_22),
.B(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_64),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_37),
.B1(n_38),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_77),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_17),
.B1(n_29),
.B2(n_15),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_73),
.B1(n_35),
.B2(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_69),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_17),
.B(n_29),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_83),
.B(n_22),
.Y(n_99)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_29),
.B1(n_15),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_34),
.B1(n_16),
.B2(n_30),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_39),
.B1(n_35),
.B2(n_16),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_44),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_79),
.Y(n_113)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_39),
.B1(n_35),
.B2(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_103),
.B1(n_110),
.B2(n_82),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_58),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_28),
.B(n_18),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_39),
.B1(n_35),
.B2(n_42),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_36),
.C(n_51),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_58),
.C(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_60),
.B1(n_75),
.B2(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_125),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_127),
.B1(n_20),
.B2(n_27),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_126),
.C(n_125),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_131),
.Y(n_154)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_120),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_133),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_81),
.B(n_79),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_107),
.B(n_98),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_32),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_33),
.C(n_32),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_24),
.B(n_19),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_33),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_92),
.A2(n_24),
.B1(n_21),
.B2(n_71),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_33),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_111),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_97),
.B(n_110),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_144),
.B(n_151),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_136),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_145),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_140),
.A2(n_108),
.B1(n_86),
.B2(n_21),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_33),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_113),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_150),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_91),
.B1(n_101),
.B2(n_94),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_168),
.B1(n_116),
.B2(n_139),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_155),
.C(n_156),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_91),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_115),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_90),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_90),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_137),
.B1(n_134),
.B2(n_128),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_168),
.B(n_173),
.Y(n_175)
);

AO22x2_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_13),
.CI(n_12),
.CON(n_201),
.SN(n_201)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_30),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_13),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_181),
.B1(n_197),
.B2(n_201),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_170),
.B1(n_160),
.B2(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_186),
.Y(n_219)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_129),
.B(n_27),
.C(n_23),
.D(n_20),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_205),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_0),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_8),
.B(n_14),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_169),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_148),
.A2(n_19),
.B(n_27),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_23),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_0),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_153),
.C(n_143),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_218),
.C(n_203),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_170),
.B1(n_166),
.B2(n_145),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_223),
.B1(n_175),
.B2(n_197),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_190),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_221),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_181),
.B1(n_198),
.B2(n_191),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_0),
.C(n_1),
.Y(n_218)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_12),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_12),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_205),
.Y(n_233)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_196),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_242),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_229),
.B1(n_217),
.B2(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_246),
.B1(n_248),
.B2(n_226),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_211),
.C(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_179),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_212),
.B(n_230),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_251),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_177),
.B1(n_188),
.B2(n_189),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_191),
.B(n_185),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_192),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_240),
.C(n_201),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_4),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_216),
.B1(n_223),
.B2(n_214),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_251),
.B(n_239),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_183),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_268),
.B1(n_233),
.B2(n_236),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_9),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_208),
.B1(n_201),
.B2(n_176),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_252),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_272),
.A2(n_273),
.B1(n_282),
.B2(n_254),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_275),
.C(n_278),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_240),
.C(n_2),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_10),
.B(n_9),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_4),
.B(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_10),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_1),
.C(n_2),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_264),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_1),
.B(n_3),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_259),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_268),
.Y(n_285)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_256),
.B(n_257),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_286),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_288),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_263),
.C(n_261),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_266),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_261),
.B(n_254),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_5),
.C(n_6),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_4),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_283),
.B(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_302),
.C(n_286),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_300),
.B(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_6),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_312),
.B(n_309),
.C(n_304),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.B(n_309),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_314),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_6),
.B(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_7),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_7),
.Y(n_318)
);


endmodule