module fake_jpeg_11606_n_622 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_622);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_622;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_76),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_73),
.Y(n_216)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_0),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_88),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_93),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_105),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_17),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_42),
.A2(n_2),
.B(n_3),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_106),
.B(n_2),
.Y(n_191)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_50),
.Y(n_118)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_124),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_55),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

BUFx2_ASAP7_75t_SL g212 ( 
.A(n_127),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_19),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_30),
.B1(n_56),
.B2(n_48),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_130),
.A2(n_201),
.B1(n_37),
.B2(n_33),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_49),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_153),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_69),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_132),
.B(n_142),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_63),
.A2(n_30),
.B1(n_56),
.B2(n_48),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_147),
.A2(n_177),
.B1(n_37),
.B2(n_36),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_92),
.A2(n_58),
.B1(n_57),
.B2(n_52),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_149),
.A2(n_196),
.B1(n_79),
.B2(n_82),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_41),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_166),
.C(n_24),
.Y(n_238)
);

FAx1_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_57),
.CI(n_52),
.CON(n_166),
.SN(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_186),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_61),
.A2(n_39),
.B1(n_24),
.B2(n_46),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_49),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_181),
.B(n_215),
.Y(n_260)
);

BUFx4f_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_62),
.A2(n_51),
.B1(n_33),
.B2(n_41),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_65),
.A2(n_20),
.B1(n_46),
.B2(n_40),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_77),
.A2(n_20),
.B1(n_40),
.B2(n_39),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_102),
.Y(n_243)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_102),
.B(n_51),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_77),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_36),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_220),
.A2(n_230),
.B1(n_218),
.B2(n_208),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_145),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_221),
.Y(n_325)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_158),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_233),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_226),
.B(n_231),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_227),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_228),
.Y(n_344)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_152),
.A2(n_72),
.B1(n_78),
.B2(n_66),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_235),
.B(n_238),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_236),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_239),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_240),
.B(n_268),
.Y(n_305)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_243),
.B(n_256),
.Y(n_341)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_244),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_169),
.B(n_152),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_245),
.B(n_253),
.Y(n_335)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_247),
.Y(n_319)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_166),
.A2(n_95),
.B1(n_88),
.B2(n_90),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_121),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_156),
.B(n_104),
.C(n_101),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_205),
.C(n_195),
.Y(n_324)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_135),
.A2(n_99),
.B1(n_91),
.B2(n_87),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_257),
.A2(n_258),
.B1(n_265),
.B2(n_277),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_134),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_191),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_199),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_179),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_154),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_267),
.B(n_269),
.Y(n_351)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_179),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_184),
.B(n_12),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_270),
.B(n_271),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_184),
.B(n_12),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_272),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_138),
.B(n_13),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_273),
.B(n_274),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_275),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_176),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_276),
.Y(n_333)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_144),
.Y(n_277)
);

AO22x1_ASAP7_75t_SL g278 ( 
.A1(n_129),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_278),
.B(n_290),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_14),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_14),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_329)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_183),
.Y(n_281)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_163),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_216),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_163),
.B1(n_160),
.B2(n_141),
.Y(n_297)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVx6_ASAP7_75t_SL g285 ( 
.A(n_212),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_174),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_192),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_150),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_136),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_292),
.Y(n_302)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_137),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_159),
.A2(n_14),
.B1(n_16),
.B2(n_170),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_242),
.B(n_222),
.Y(n_349)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_203),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_294),
.Y(n_307)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_167),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_147),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_343),
.C(n_246),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_297),
.A2(n_349),
.B(n_256),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_298),
.A2(n_310),
.B1(n_316),
.B2(n_321),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_301),
.B(n_250),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_218),
.B1(n_208),
.B2(n_177),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_235),
.A2(n_148),
.B1(n_193),
.B2(n_164),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_315),
.A2(n_317),
.B1(n_336),
.B2(n_342),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_226),
.A2(n_193),
.B1(n_164),
.B2(n_148),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_232),
.A2(n_259),
.B1(n_254),
.B2(n_233),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_219),
.A2(n_212),
.B(n_140),
.C(n_143),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_334),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_205),
.B1(n_195),
.B2(n_206),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_342),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_237),
.A2(n_161),
.B1(n_288),
.B2(n_264),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_332),
.B1(n_337),
.B2(n_275),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_182),
.B1(n_187),
.B2(n_168),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_241),
.B(n_194),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_257),
.A2(n_165),
.B1(n_188),
.B2(n_171),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_249),
.A2(n_151),
.B1(n_16),
.B2(n_162),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_227),
.A2(n_162),
.A3(n_291),
.B1(n_252),
.B2(n_234),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_223),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_265),
.A2(n_258),
.B1(n_281),
.B2(n_248),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_SL g343 ( 
.A(n_282),
.B(n_236),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_354),
.B(n_373),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_244),
.B1(n_272),
.B2(n_268),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_355),
.A2(n_359),
.B1(n_375),
.B2(n_340),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_357),
.A2(n_364),
.B(n_365),
.Y(n_412)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_294),
.B1(n_266),
.B2(n_221),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_361),
.A2(n_362),
.B1(n_374),
.B2(n_382),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_300),
.A2(n_229),
.B1(n_247),
.B2(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_343),
.B(n_222),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_366),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_335),
.B(n_225),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_370),
.Y(n_409)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_302),
.Y(n_369)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_228),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_303),
.Y(n_372)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_300),
.A2(n_263),
.B1(n_336),
.B2(n_315),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_305),
.A2(n_317),
.B1(n_321),
.B2(n_298),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_357),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_350),
.A2(n_296),
.B(n_338),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_381),
.B(n_393),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_295),
.B(n_324),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_380),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_309),
.A2(n_308),
.B1(n_339),
.B2(n_349),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_379),
.A2(n_304),
.B(n_325),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_328),
.B(n_351),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_313),
.B(n_332),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_349),
.A2(n_334),
.B1(n_348),
.B2(n_331),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_333),
.C(n_318),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_389),
.C(n_345),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_323),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g408 ( 
.A1(n_384),
.A2(n_386),
.B(n_396),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_301),
.B(n_333),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_388),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_323),
.Y(n_386)
);

AO21x2_ASAP7_75t_SL g387 ( 
.A1(n_309),
.A2(n_319),
.B(n_303),
.Y(n_387)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_319),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_330),
.C(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_328),
.B(n_308),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_391),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_306),
.B(n_330),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_297),
.A2(n_337),
.B(n_329),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_316),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_353),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_311),
.A2(n_327),
.B1(n_314),
.B2(n_344),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_395),
.A2(n_314),
.B1(n_327),
.B2(n_325),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_322),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_399),
.B(n_389),
.Y(n_456)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_340),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_403),
.B(n_376),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_348),
.B1(n_312),
.B2(n_346),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_369),
.B(n_299),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_415),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_299),
.C(n_346),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_424),
.C(n_389),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_388),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_419),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_371),
.B(n_322),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_418),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_383),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_375),
.A2(n_344),
.B1(n_312),
.B2(n_325),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_429),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_381),
.B(n_382),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_358),
.B(n_363),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_433),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_364),
.A2(n_360),
.B(n_365),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_428),
.A2(n_400),
.B(n_411),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_353),
.B1(n_370),
.B2(n_360),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_431),
.A2(n_387),
.B1(n_356),
.B2(n_374),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_377),
.B(n_390),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_434),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_380),
.B(n_385),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_437),
.B(n_449),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_438),
.B(n_465),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_366),
.Y(n_441)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_434),
.Y(n_442)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_442),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_443),
.A2(n_459),
.B(n_425),
.C(n_412),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_449),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_446),
.A2(n_428),
.B(n_412),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_411),
.A2(n_379),
.B(n_393),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_384),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_448),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_386),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_458),
.B1(n_467),
.B2(n_420),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_456),
.C(n_419),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_457),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_367),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_387),
.B1(n_356),
.B2(n_394),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_426),
.A2(n_387),
.B1(n_372),
.B2(n_355),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_460),
.Y(n_491)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_463),
.B(n_464),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_391),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_421),
.B(n_373),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_387),
.B1(n_359),
.B2(n_362),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_414),
.B(n_396),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_448),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_445),
.B(n_421),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_470),
.B(n_401),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_441),
.A2(n_422),
.B(n_416),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_472),
.B(n_466),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_473),
.A2(n_450),
.B(n_460),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_424),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_475),
.B(n_476),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_410),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_410),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_492),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_451),
.A2(n_402),
.B1(n_406),
.B2(n_429),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_479),
.A2(n_488),
.B1(n_454),
.B2(n_453),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_481),
.A2(n_483),
.B1(n_458),
.B2(n_467),
.Y(n_505)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_439),
.A2(n_430),
.B1(n_398),
.B2(n_405),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_490),
.C(n_493),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_399),
.C(n_403),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_444),
.B(n_414),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_398),
.C(n_405),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_447),
.B(n_408),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_494),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_496),
.A2(n_439),
.B1(n_443),
.B2(n_436),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_455),
.B(n_409),
.C(n_432),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_499),
.C(n_500),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_468),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_409),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_432),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_503),
.A2(n_506),
.B1(n_522),
.B2(n_495),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_505),
.A2(n_510),
.B(n_498),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_479),
.A2(n_436),
.B1(n_453),
.B2(n_466),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_471),
.Y(n_507)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_507),
.Y(n_552)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_508),
.Y(n_530)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_459),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_511),
.B(n_523),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_457),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_525),
.Y(n_537)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_514),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g515 ( 
.A(n_473),
.B(n_461),
.CI(n_469),
.CON(n_515),
.SN(n_515)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_515),
.B(n_520),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_516),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_483),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_489),
.B(n_463),
.C(n_462),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_524),
.C(n_487),
.Y(n_531)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_440),
.C(n_442),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_490),
.B(n_440),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_527),
.B1(n_488),
.B2(n_480),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_484),
.A2(n_430),
.B1(n_459),
.B2(n_435),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_491),
.Y(n_539)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_474),
.Y(n_529)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_529),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_531),
.B(n_541),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_532),
.B(n_535),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_493),
.C(n_492),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_533),
.B(n_545),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_519),
.B(n_487),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_536),
.A2(n_505),
.B1(n_510),
.B2(n_503),
.Y(n_557)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_539),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_502),
.A2(n_495),
.B(n_481),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_540),
.A2(n_511),
.B(n_506),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_477),
.Y(n_541)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_497),
.Y(n_543)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_543),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_500),
.C(n_481),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_518),
.B(n_499),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_548),
.B(n_513),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_459),
.Y(n_549)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_549),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_481),
.C(n_435),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_551),
.B(n_519),
.C(n_524),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_544),
.B(n_504),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_553),
.A2(n_552),
.B1(n_543),
.B2(n_561),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_517),
.Y(n_556)
);

CKINVDCx14_ASAP7_75t_R g581 ( 
.A(n_556),
.Y(n_581)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_540),
.A2(n_511),
.B(n_515),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_558),
.A2(n_566),
.B(n_532),
.Y(n_572)
);

FAx1_ASAP7_75t_SL g562 ( 
.A(n_545),
.B(n_515),
.CI(n_517),
.CON(n_562),
.SN(n_562)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_541),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_548),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_525),
.C(n_531),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_567),
.B(n_569),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_537),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_546),
.B(n_528),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_570),
.Y(n_574)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_571),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_572),
.A2(n_573),
.B(n_566),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_558),
.A2(n_534),
.B(n_536),
.Y(n_573)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_575),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_576),
.B(n_580),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_560),
.A2(n_538),
.B1(n_534),
.B2(n_530),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_577),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_584),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_553),
.B(n_546),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_537),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_585),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_557),
.B(n_559),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_560),
.A2(n_530),
.B1(n_539),
.B2(n_551),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_581),
.B(n_567),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_588),
.B(n_589),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_576),
.B(n_555),
.C(n_564),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_577),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_572),
.A2(n_570),
.B(n_565),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_594),
.B(n_596),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_583),
.A2(n_565),
.B1(n_554),
.B2(n_562),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_564),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_597),
.B(n_568),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_592),
.B(n_579),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_598),
.B(n_595),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_599),
.A2(n_601),
.B(n_603),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_592),
.B(n_584),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_563),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_605),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_586),
.A2(n_583),
.B(n_562),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_606),
.B(n_600),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_609),
.Y(n_615)
);

AO221x1_ASAP7_75t_L g611 ( 
.A1(n_606),
.A2(n_594),
.B1(n_593),
.B2(n_587),
.C(n_554),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_608),
.C(n_574),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_604),
.A2(n_590),
.B(n_593),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_612),
.B(n_601),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_610),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_613),
.A2(n_614),
.B(n_616),
.Y(n_618)
);

AOI321xp33_ASAP7_75t_L g617 ( 
.A1(n_615),
.A2(n_596),
.A3(n_573),
.B1(n_559),
.B2(n_509),
.C(n_535),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_617),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_618),
.B(n_547),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_620),
.A2(n_547),
.B1(n_459),
.B2(n_395),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_621),
.B(n_459),
.Y(n_622)
);


endmodule