module real_jpeg_16213_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_584, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_584;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_123),
.B1(n_128),
.B2(n_130),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_0),
.A2(n_130),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_0),
.A2(n_130),
.B1(n_364),
.B2(n_367),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_80),
.B1(n_159),
.B2(n_162),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_2),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_162),
.B1(n_267),
.B2(n_271),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_2),
.A2(n_162),
.B1(n_443),
.B2(n_448),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_2),
.A2(n_162),
.B1(n_503),
.B2(n_508),
.Y(n_502)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_3),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_3),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g490 ( 
.A(n_3),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_4),
.A2(n_71),
.B1(n_283),
.B2(n_286),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_4),
.A2(n_71),
.B1(n_140),
.B2(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_4),
.A2(n_71),
.B1(n_423),
.B2(n_425),
.Y(n_422)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_5),
.B(n_163),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_5),
.A2(n_51),
.A3(n_87),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_5),
.B(n_75),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_5),
.A2(n_79),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_5),
.A2(n_102),
.B1(n_524),
.B2(n_531),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_6),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_112),
.B1(n_117),
.B2(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_7),
.A2(n_117),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_7),
.A2(n_117),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_7),
.A2(n_117),
.B1(n_567),
.B2(n_569),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_8),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_8),
.A2(n_185),
.B1(n_220),
.B2(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_9),
.Y(n_224)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_9),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_9),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_113),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_10),
.A2(n_173),
.B1(n_328),
.B2(n_333),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_10),
.A2(n_173),
.B1(n_574),
.B2(n_577),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_11),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_12),
.A2(n_35),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_12),
.A2(n_35),
.B1(n_375),
.B2(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_12),
.A2(n_35),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_13),
.A2(n_136),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_13),
.A2(n_136),
.B1(n_437),
.B2(n_441),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_13),
.A2(n_136),
.B1(n_521),
.B2(n_525),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_15),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_15),
.A2(n_231),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_15),
.A2(n_231),
.B1(n_307),
.B2(n_313),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_15),
.A2(n_231),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_16),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g184 ( 
.A(n_16),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_16),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g570 ( 
.A(n_17),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_554),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_393),
.B(n_549),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_320),
.C(n_355),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_258),
.B(n_290),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_24),
.B(n_258),
.C(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_164),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_25),
.B(n_165),
.C(n_225),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_76),
.C(n_134),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_27),
.B(n_134),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_42),
.B1(n_65),
.B2(n_74),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_29),
.A2(n_75),
.B1(n_266),
.B2(n_278),
.Y(n_265)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_33),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_34),
.Y(n_270)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_38),
.Y(n_577)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_40),
.Y(n_301)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_41),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_42),
.A2(n_65),
.B1(n_74),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_42),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_42),
.A2(n_74),
.B1(n_252),
.B2(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_42),
.A2(n_74),
.B1(n_298),
.B2(n_469),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_42),
.A2(n_74),
.B1(n_363),
.B2(n_573),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_57),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22x1_ASAP7_75t_SL g150 ( 
.A1(n_49),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_150)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_54),
.Y(n_366)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_55),
.Y(n_348)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_58),
.Y(n_230)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_58),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_59),
.Y(n_332)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_59),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_61),
.Y(n_414)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_70),
.Y(n_576)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_75),
.A2(n_266),
.B1(n_278),
.B2(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_75),
.A2(n_278),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_76),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_101),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_77),
.B(n_101),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_90),
.B2(n_94),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_SL g280 ( 
.A1(n_78),
.A2(n_79),
.B(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_79),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_79),
.B(n_484),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_79),
.A2(n_483),
.B(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_79),
.B(n_131),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g537 ( 
.A(n_79),
.B(n_189),
.Y(n_537)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_89),
.Y(n_255)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_89),
.Y(n_371)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_89),
.Y(n_473)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_145),
.B(n_150),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_97),
.Y(n_248)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_97),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_110),
.B1(n_122),
.B2(n_131),
.Y(n_101)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_102),
.A2(n_122),
.B1(n_169),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_102),
.A2(n_180),
.B(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_102),
.A2(n_453),
.B1(n_456),
.B2(n_460),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_102),
.A2(n_502),
.B1(n_524),
.B2(n_534),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_103),
.A2(n_167),
.B1(n_306),
.B2(n_422),
.Y(n_421)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_106),
.Y(n_241)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_109),
.Y(n_521)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_111),
.A2(n_167),
.B1(n_306),
.B2(n_314),
.Y(n_305)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_112),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_115),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_116),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_132),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_133),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_144),
.B1(n_157),
.B2(n_163),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_135),
.A2(n_144),
.B1(n_163),
.B2(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_143),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_143),
.Y(n_388)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_143),
.Y(n_568)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_144),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_155),
.Y(n_257)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_158),
.A2(n_244),
.B1(n_245),
.B2(n_250),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_225),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_186),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_166),
.A2(n_187),
.B(n_209),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_179),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_167),
.A2(n_501),
.B1(n_510),
.B2(n_512),
.Y(n_500)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_183),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_209),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_200),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_188),
.A2(n_210),
.B1(n_282),
.B2(n_289),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_188),
.A2(n_210),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_188),
.A2(n_210),
.B1(n_436),
.B2(n_442),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_188),
.A2(n_210),
.B1(n_403),
.B2(n_442),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_188),
.A2(n_210),
.B1(n_436),
.B2(n_494),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_188),
.A2(n_210),
.B(n_374),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_189),
.A2(n_201),
.B1(n_228),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_189),
.A2(n_228),
.B1(n_402),
.B2(n_408),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_196),
.Y(n_424)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_213),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_216),
.Y(n_482)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_242),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_237),
.Y(n_226)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_236),
.Y(n_486)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_243),
.B(n_251),
.C(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_244),
.A2(n_250),
.B1(n_342),
.B2(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_244),
.A2(n_250),
.B1(n_384),
.B2(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_259),
.A2(n_260),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_264),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_279),
.C(n_281),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_281),
.Y(n_293)
);

INVx8_ASAP7_75t_L g470 ( 
.A(n_267),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_282),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_285),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_317),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_291),
.B(n_317),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_292),
.B(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_294),
.B(n_295),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_305),
.C(n_316),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_296),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_305),
.B(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_311),
.Y(n_454)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_314),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_315),
.Y(n_511)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

A2O1A1O1Ixp25_ASAP7_75t_L g549 ( 
.A1(n_320),
.A2(n_355),
.B(n_550),
.C(n_552),
.D(n_553),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_354),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_321),
.B(n_354),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_339),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_391),
.C(n_392),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_335),
.B1(n_336),
.B2(n_338),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_326),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_336),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_331),
.Y(n_481)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_332),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_336),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_335),
.A2(n_389),
.B1(n_561),
.B2(n_584),
.Y(n_560)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_353),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_345),
.C(n_353),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_390),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_356),
.B(n_390),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_357),
.B(n_557),
.C(n_558),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_378),
.Y(n_358)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_359),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_372),
.B(n_377),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_372),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_377),
.A2(n_563),
.B1(n_580),
.B2(n_581),
.Y(n_562)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_377),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_378),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_381),
.B2(n_389),
.Y(n_378)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_382),
.Y(n_561)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_430),
.B(n_548),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_395),
.B(n_397),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.C(n_409),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_399),
.B(n_544),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_401),
.A2(n_409),
.B1(n_410),
.B2(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_420),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_411),
.A2(n_420),
.B1(n_421),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_542),
.B(n_547),
.Y(n_430)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_476),
.B(n_541),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_463),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_433),
.B(n_463),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_452),
.C(n_461),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_435),
.B1(n_461),
.B2(n_462),
.Y(n_497)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_450),
.Y(n_495)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_452),
.B(n_497),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

OAI32xp33_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_480),
.A3(n_482),
.B1(n_483),
.B2(n_487),
.Y(n_479)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

BUFx5_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_464),
.B(n_467),
.C(n_475),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_467),
.A2(n_468),
.B1(n_474),
.B2(n_475),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_498),
.B(n_540),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_496),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_478),
.B(n_496),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_492),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_479),
.A2(n_492),
.B1(n_493),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_479),
.Y(n_514)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_491),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_515),
.B(n_539),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_513),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_500),
.B(n_513),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_532),
.B(n_538),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_523),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_522),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_537),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_537),
.Y(n_538)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx12f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_SL g542 ( 
.A(n_543),
.B(n_546),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_543),
.B(n_546),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_582),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_559),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_556),
.B(n_559),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_562),
.Y(n_559)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_563),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_564),
.A2(n_565),
.B1(n_571),
.B2(n_579),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_571),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_578),
.Y(n_571)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);


endmodule