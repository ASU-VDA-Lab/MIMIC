module real_jpeg_5527_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_1),
.B(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_1),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_3),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_4),
.Y(n_164)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_10),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_12),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_12),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_13),
.B(n_110),
.Y(n_109)
);

XNOR2x2_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_120),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_119),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_72),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_18),
.B(n_72),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.C(n_54),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_20),
.B(n_28),
.C(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_21),
.Y(n_139)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_22),
.Y(n_170)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_33),
.B(n_37),
.Y(n_105)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_39),
.B(n_54),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_52),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_40),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_41),
.B(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_45),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_62),
.C(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_101),
.B2(n_102),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_89),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_118),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_140),
.B(n_184),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_124),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_138),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_128),
.B1(n_138),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_178),
.B(n_183),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_161),
.B(n_177),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_150),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_147),
.C(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_171),
.B(n_176),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_175),
.Y(n_176)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);


endmodule