module real_jpeg_17450_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_70;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_41;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_0),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_0),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_0),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_0),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_0),
.B(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_2),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_4),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_4),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_5),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_102),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_8),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_10),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_10),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_10),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_13),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_14),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_14),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_14),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_15),
.Y(n_50)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_160),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_159),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_132),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_20),
.B(n_132),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_91),
.B2(n_92),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_69),
.B2(n_70),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_29),
.Y(n_195)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_29),
.Y(n_210)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.C(n_48),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_48),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_46),
.Y(n_184)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_102),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_49),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_50),
.B(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_51),
.Y(n_227)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_68),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.C(n_77),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_77),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.C(n_89),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_78),
.A2(n_79),
.B1(n_89),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_83),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_89),
.Y(n_187)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_120),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_100),
.B(n_106),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_127),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_122),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.C(n_155),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.C(n_148),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21x1_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_188),
.B(n_243),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_164),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_185),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.C(n_181),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_204),
.B(n_242),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_202),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_200),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_193),
.A2(n_200),
.B1(n_201),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_196),
.Y(n_214)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_236),
.B(n_241),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_224),
.B(n_235),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_207),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_217),
.C(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_229),
.B(n_234),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);


endmodule