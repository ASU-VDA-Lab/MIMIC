module fake_jpeg_2270_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_2),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_39),
.B1(n_51),
.B2(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_36),
.C(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_49),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_56),
.B(n_54),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_77),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_52),
.B1(n_51),
.B2(n_56),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_64),
.B1(n_48),
.B2(n_34),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_56),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_64),
.B1(n_60),
.B2(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_89),
.B1(n_93),
.B2(n_32),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_64),
.B1(n_65),
.B2(n_48),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_92),
.B1(n_75),
.B2(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_6),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_7),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_8),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_20),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_108),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_18),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_21),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_111),
.B1(n_88),
.B2(n_10),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_31),
.C(n_30),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_112),
.CI(n_24),
.CON(n_115),
.SN(n_115)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_28),
.C(n_26),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_82),
.B(n_83),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_117),
.B(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_124),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_100),
.B(n_107),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_89),
.B1(n_93),
.B2(n_88),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_125),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_23),
.B(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_121),
.C(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_126),
.B(n_119),
.Y(n_136)
);

NAND4xp25_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.C(n_133),
.D(n_132),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_129),
.A3(n_134),
.B1(n_118),
.B2(n_116),
.C1(n_115),
.C2(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_11),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_14),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_115),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_15),
.B(n_16),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_15),
.Y(n_144)
);


endmodule