module fake_jpeg_12375_n_96 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_31),
.B(n_33),
.Y(n_36)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_32),
.B1(n_22),
.B2(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_17),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_5),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_11),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_11),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_19),
.B(n_16),
.C(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_30),
.C(n_27),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_26),
.B(n_14),
.Y(n_65)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_27),
.C(n_28),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_18),
.C(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_16),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_45),
.C(n_8),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_68),
.B(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_8),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_52),
.B1(n_26),
.B2(n_49),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_74),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_76),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_56),
.B(n_54),
.C(n_47),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_59),
.C(n_66),
.Y(n_79)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_9),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_56),
.B1(n_46),
.B2(n_51),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_69),
.A3(n_73),
.B1(n_46),
.B2(n_78),
.C(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_59),
.C(n_67),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_59),
.C(n_66),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_72),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_65),
.Y(n_88)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_73),
.B1(n_74),
.B2(n_72),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_92),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_86),
.C(n_10),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

AOI31xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_93),
.A3(n_5),
.B(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);


endmodule