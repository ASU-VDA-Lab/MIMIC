module real_jpeg_8258_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_327, n_326, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_327;
input n_326;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_68),
.B1(n_69),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_2),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_142),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_142),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_142),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_4),
.A2(n_52),
.B1(n_68),
.B2(n_69),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_9),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_9),
.A2(n_68),
.B1(n_69),
.B2(n_113),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_113),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_113),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_62),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_62),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_11),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_101),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_101),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_101),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_12),
.A2(n_44),
.B1(n_68),
.B2(n_69),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_31),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_13),
.B(n_31),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_13),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_27),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_13),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_13),
.B(n_53),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_28),
.B(n_48),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_126),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_15),
.A2(n_37),
.B1(n_68),
.B2(n_69),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_16),
.A2(n_68),
.B1(n_69),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_16),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_106),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_106),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_17),
.A2(n_68),
.B1(n_69),
.B2(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_81),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_73),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_54),
.B1(n_55),
.B2(n_72),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_25),
.A2(n_34),
.B1(n_86),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_26),
.A2(n_30),
.B1(n_58),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_26),
.A2(n_30),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_30),
.B1(n_152),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_26),
.A2(n_30),
.B1(n_168),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_26),
.A2(n_30),
.B1(n_208),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_26),
.A2(n_30),
.B1(n_219),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_26),
.A2(n_30),
.B1(n_245),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_50)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_29),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_30),
.B(n_126),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_31),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_31),
.B(n_33),
.Y(n_156)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_32),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_46),
.B1(n_50),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_47),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_43),
.A2(n_47),
.B(n_126),
.C(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_45),
.A2(n_53),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_50),
.B1(n_61),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_46),
.A2(n_50),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_46),
.A2(n_50),
.B1(n_223),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_46),
.A2(n_50),
.B1(n_248),
.B2(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_46),
.A2(n_50),
.B1(n_80),
.B2(n_266),
.Y(n_290)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.C(n_63),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_63),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_67),
.B(n_71),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_67),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_64),
.A2(n_67),
.B1(n_112),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_64),
.A2(n_67),
.B1(n_139),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_64),
.A2(n_67),
.B1(n_148),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_64),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_64),
.A2(n_67),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_64),
.A2(n_67),
.B1(n_231),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_64),
.A2(n_67),
.B1(n_240),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_67),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_67),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_71),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.C(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_311),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.C(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_79),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_79),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_82),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI321xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_308),
.A3(n_318),
.B1(n_323),
.B2(n_324),
.C(n_326),
.Y(n_89)
);

AOI321xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_256),
.A3(n_296),
.B1(n_302),
.B2(n_307),
.C(n_327),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_213),
.C(n_252),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_183),
.B(n_212),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_162),
.B(n_182),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_144),
.B(n_161),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_133),
.B(n_143),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_119),
.B(n_132),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_107),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_102),
.A2(n_103),
.B1(n_160),
.B2(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_123),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_118),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_127),
.B(n_131),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_125),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_141),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_123),
.A2(n_124),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_123),
.A2(n_124),
.B1(n_194),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_123),
.A2(n_124),
.B1(n_228),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_123),
.A2(n_124),
.B(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.C(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_146),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.CI(n_153),
.CON(n_146),
.SN(n_146)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_176),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_178),
.C(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_174),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.C(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_185),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_198),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_197),
.C(n_198),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_192),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_206),
.B2(n_207),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_206),
.C(n_209),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_203),
.A2(n_205),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_214),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_233),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_215),
.B(n_233),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.C(n_232),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_224),
.C(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_232),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_250),
.B2(n_251),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_241),
.C(n_251),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_239),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_246),
.C(n_249),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_250),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_254),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_275),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_257),
.B(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_268),
.C(n_274),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_259),
.B1(n_268),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_264),
.C(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_262),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_268),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_270),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_269),
.A2(n_290),
.B(n_292),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_271),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_271),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_294),
.B2(n_295),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_287),
.C(n_295),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_283),
.B(n_285),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_283),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_285),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_285),
.A2(n_310),
.B1(n_314),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_316),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.C(n_315),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);


endmodule