module fake_netlist_1_6403_n_723 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_723);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_723;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_67), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_7), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_19), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_15), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_81), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_72), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_3), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_57), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_18), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_41), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_73), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_37), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_53), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_38), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_5), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_9), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_23), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_25), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_27), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_18), .B(n_33), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_36), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_48), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_29), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_70), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_35), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_6), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_22), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_8), .Y(n_131) );
OR2x6_ASAP7_75t_L g132 ( .A(n_85), .B(n_1), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_119), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_116), .B(n_1), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_117), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_131), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_97), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_100), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_105), .Y(n_140) );
NOR2xp33_ASAP7_75t_R g141 ( .A(n_84), .B(n_45), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_116), .B(n_2), .Y(n_142) );
NOR2xp67_ASAP7_75t_L g143 ( .A(n_82), .B(n_4), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_108), .Y(n_145) );
INVx1_ASAP7_75t_SL g146 ( .A(n_115), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_83), .Y(n_148) );
NOR2xp67_ASAP7_75t_L g149 ( .A(n_83), .B(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
XOR2xp5_ASAP7_75t_L g151 ( .A(n_90), .B(n_7), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_116), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_110), .B(n_8), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_89), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_104), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_109), .B(n_10), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_104), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_130), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_93), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_93), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_86), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_91), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_91), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_88), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_96), .Y(n_172) );
NOR2xp33_ASAP7_75t_R g173 ( .A(n_88), .B(n_49), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_96), .B(n_10), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_98), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_92), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_174), .B(n_98), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_144), .B(n_111), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_174), .A2(n_92), .B1(n_128), .B2(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_133), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
BUFx4_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_136), .B(n_94), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_160), .B(n_94), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_174), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_160), .B(n_95), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_153), .B(n_111), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_133), .B(n_95), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_135), .B(n_99), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_168), .B(n_99), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_163), .B(n_118), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_150), .A2(n_118), .B(n_128), .C(n_126), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_163), .B(n_120), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_137), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_171), .B(n_120), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_168), .B(n_176), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_176), .B(n_102), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_145), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
BUFx4_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_169), .B(n_101), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_147), .Y(n_218) );
INVxp67_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_170), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_148), .A2(n_101), .B1(n_106), .B2(n_122), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_164), .B(n_102), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_132), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_145), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_152), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_172), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_175), .B(n_103), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_162), .B(n_103), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_155), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_138), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_173), .B(n_112), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_132), .B(n_106), .Y(n_238) );
INVx5_ASAP7_75t_L g239 ( .A(n_155), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_209), .B(n_158), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_209), .B(n_143), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_197), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_212), .B(n_149), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_223), .B(n_129), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_212), .B(n_141), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_206), .B(n_112), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_182), .A2(n_122), .B1(n_123), .B2(n_114), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_229), .B(n_125), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_238), .B(n_123), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_206), .B(n_121), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_107), .B1(n_113), .B2(n_124), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_205), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_193), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_218), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_182), .A2(n_159), .B1(n_148), .B2(n_151), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
NOR2xp33_ASAP7_75t_R g265 ( .A(n_184), .B(n_159), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_193), .B(n_166), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_238), .B(n_12), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_177), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_229), .B(n_167), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_178), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_182), .A2(n_167), .B1(n_166), .B2(n_138), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_192), .B(n_167), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_180), .B(n_13), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_236), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_184), .B(n_14), .C(n_15), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_179), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_204), .B(n_167), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_183), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_179), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g285 ( .A(n_224), .B(n_16), .C(n_17), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_179), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_215), .B(n_167), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_217), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_215), .B(n_166), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_180), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_190), .Y(n_293) );
OR2x4_ASAP7_75t_L g294 ( .A(n_198), .B(n_166), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_210), .B(n_166), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_220), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_220), .B(n_20), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_189), .B(n_21), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_200), .B(n_26), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_181), .B(n_28), .Y(n_301) );
NOR3xp33_ASAP7_75t_SL g302 ( .A(n_211), .B(n_30), .C(n_32), .Y(n_302) );
AND2x6_ASAP7_75t_L g303 ( .A(n_187), .B(n_34), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_236), .Y(n_304) );
NOR2xp33_ASAP7_75t_R g305 ( .A(n_211), .B(n_39), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_196), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_194), .B(n_40), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_187), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_268), .A2(n_200), .B1(n_208), .B2(n_195), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_240), .B(n_200), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_247), .B(n_208), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_288), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_240), .B(n_195), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_249), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_306), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_249), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_249), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_255), .B(n_195), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_249), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
NOR2xp67_ASAP7_75t_R g323 ( .A(n_273), .B(n_213), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_255), .A2(n_221), .B(n_203), .C(n_222), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_241), .Y(n_329) );
O2A1O1Ixp5_ASAP7_75t_L g330 ( .A1(n_299), .A2(n_202), .B(n_237), .C(n_232), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_268), .A2(n_208), .B1(n_181), .B2(n_216), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_281), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_260), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_281), .B(n_196), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_260), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_277), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g339 ( .A1(n_255), .A2(n_199), .B1(n_216), .B2(n_219), .C1(n_230), .C2(n_213), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_260), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_301), .A2(n_199), .B(n_231), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_269), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_241), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_265), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_265), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_273), .B(n_239), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_268), .B(n_42), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_263), .B(n_43), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_269), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_286), .B(n_46), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_242), .A2(n_231), .B(n_235), .C(n_233), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_286), .B(n_47), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_300), .B(n_50), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_271), .B(n_51), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_271), .B(n_54), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_266), .A2(n_233), .B(n_235), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_272), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_281), .Y(n_360) );
INVx3_ASAP7_75t_SL g361 ( .A(n_303), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_260), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_256), .A2(n_234), .B(n_225), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_339), .A2(n_257), .B1(n_252), .B2(n_247), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_309), .A2(n_252), .B1(n_300), .B2(n_257), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_315), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_339), .A2(n_274), .B1(n_308), .B2(n_281), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_313), .B(n_245), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_310), .B(n_304), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_314), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_326), .B(n_284), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_350), .A2(n_274), .B1(n_284), .B2(n_303), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_312), .Y(n_374) );
CKINVDCx14_ASAP7_75t_R g375 ( .A(n_315), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_355), .A2(n_296), .B1(n_297), .B2(n_246), .Y(n_376) );
CKINVDCx9p33_ASAP7_75t_R g377 ( .A(n_345), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_316), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_314), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_316), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_329), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_331), .A2(n_264), .B1(n_272), .B2(n_284), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_314), .Y(n_384) );
AND2x6_ASAP7_75t_L g385 ( .A(n_355), .B(n_264), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
OR2x2_ASAP7_75t_SL g387 ( .A(n_350), .B(n_285), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_284), .B1(n_298), .B2(n_283), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_318), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_318), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_311), .A2(n_303), .B1(n_261), .B2(n_279), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_332), .B(n_289), .Y(n_392) );
INVx11_ASAP7_75t_L g393 ( .A(n_338), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_355), .A2(n_250), .B(n_358), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_326), .B(n_261), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_314), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_320), .A2(n_279), .B1(n_245), .B2(n_262), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_346), .B1(n_338), .B2(n_344), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_378), .B(n_332), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_382), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_373), .B(n_302), .C(n_278), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_370), .B(n_346), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_378), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_385), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_361), .B1(n_348), .B2(n_349), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_392), .B(n_337), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
OR2x6_ASAP7_75t_L g412 ( .A(n_388), .B(n_349), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_370), .A2(n_341), .B1(n_348), .B2(n_361), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_368), .A2(n_341), .B1(n_361), .B2(n_305), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_394), .A2(n_324), .B(n_330), .C(n_307), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_365), .A2(n_305), .B1(n_326), .B2(n_256), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_385), .A2(n_326), .B1(n_323), .B2(n_342), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_376), .A2(n_337), .B1(n_342), .B2(n_326), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_381), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_366), .A2(n_326), .B1(n_294), .B2(n_343), .Y(n_421) );
BUFx4f_ASAP7_75t_SL g422 ( .A(n_393), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_369), .A2(n_296), .B1(n_253), .B2(n_254), .C(n_248), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_343), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_376), .A2(n_357), .B(n_356), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_389), .B(n_351), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_389), .B(n_390), .Y(n_428) );
NOR2xp33_ASAP7_75t_R g429 ( .A(n_422), .B(n_375), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_402), .A2(n_385), .B1(n_374), .B2(n_367), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_419), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_406), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_410), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_410), .B(n_390), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_398), .B1(n_383), .B2(n_396), .C(n_380), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_401), .B(n_386), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_408), .A2(n_294), .B1(n_385), .B2(n_387), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_419), .A2(n_379), .B(n_356), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_404), .B(n_386), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_404), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_402), .A2(n_385), .B1(n_391), .B2(n_307), .Y(n_446) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_399), .A2(n_387), .B1(n_243), .B2(n_244), .C1(n_290), .C2(n_293), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_404), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_400), .B(n_386), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_425), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_426), .A2(n_357), .B(n_251), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_351), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_423), .B(n_347), .C(n_333), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_409), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_409), .B(n_359), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_408), .A2(n_360), .B1(n_333), .B2(n_359), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_395), .B1(n_372), .B2(n_295), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_414), .A2(n_395), .B1(n_372), .B2(n_295), .Y(n_458) );
OAI33xp33_ASAP7_75t_L g459 ( .A1(n_420), .A2(n_275), .A3(n_282), .B1(n_251), .B2(n_287), .B3(n_291), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_409), .B(n_397), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_428), .B(n_384), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_428), .B(n_424), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_426), .A2(n_384), .B(n_371), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_424), .B(n_371), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_435), .B(n_427), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_435), .B(n_425), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_450), .B(n_427), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_450), .B(n_407), .Y(n_468) );
AOI31xp33_ASAP7_75t_L g469 ( .A1(n_447), .A2(n_418), .A3(n_417), .B(n_416), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_434), .B(n_406), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_449), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_449), .B(n_407), .Y(n_477) );
OAI221xp5_ASAP7_75t_L g478 ( .A1(n_430), .A2(n_415), .B1(n_412), .B2(n_411), .C(n_335), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_448), .B(n_406), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_434), .B(n_406), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_436), .B(n_462), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_444), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_434), .B(n_411), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_447), .B(n_421), .C(n_353), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_436), .B(n_411), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_454), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_454), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_438), .B(n_352), .C(n_354), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_439), .B(n_406), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_462), .B(n_412), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_461), .B(n_412), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_440), .A2(n_335), .A3(n_377), .B(n_258), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_439), .B(n_406), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_438), .B(n_372), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_442), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_445), .B(n_412), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_439), .B(n_412), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_443), .B(n_397), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g506 ( .A(n_445), .B(n_397), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_461), .B(n_452), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_443), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_452), .B(n_397), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_455), .Y(n_511) );
NAND2x1_ASAP7_75t_SL g512 ( .A(n_455), .B(n_372), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_464), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_455), .B(n_314), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_470), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_466), .B(n_464), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_470), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_502), .B(n_433), .Y(n_518) );
NOR2xp33_ASAP7_75t_SL g519 ( .A(n_498), .B(n_429), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_497), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_487), .Y(n_521) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_487), .B(n_463), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_466), .B(n_460), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_469), .B(n_459), .C(n_453), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_503), .B(n_433), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_475), .B(n_460), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_465), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_507), .B(n_460), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_481), .B(n_456), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_502), .B(n_441), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_472), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_474), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_503), .B(n_463), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_465), .B(n_458), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_507), .B(n_463), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_478), .A2(n_446), .A3(n_457), .B(n_453), .Y(n_539) );
AND3x2_ASAP7_75t_L g540 ( .A(n_488), .B(n_393), .C(n_441), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_513), .B(n_451), .Y(n_541) );
AND4x1_ASAP7_75t_L g542 ( .A(n_485), .B(n_459), .C(n_363), .D(n_270), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_463), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_500), .B(n_451), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_491), .B(n_463), .C(n_186), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_488), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_468), .B(n_441), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_513), .B(n_451), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_467), .B(n_451), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_468), .B(n_441), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_476), .Y(n_551) );
NAND4xp25_ASAP7_75t_L g552 ( .A(n_486), .B(n_267), .C(n_358), .D(n_395), .Y(n_552) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_505), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_482), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_477), .B(n_335), .Y(n_556) );
NAND2xp33_ASAP7_75t_SL g557 ( .A(n_512), .B(n_317), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_482), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_489), .B(n_317), .Y(n_560) );
NOR3xp33_ASAP7_75t_SL g561 ( .A(n_510), .B(n_267), .C(n_58), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_484), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_509), .B(n_317), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_497), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_497), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_493), .B(n_321), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_504), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_508), .B(n_317), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_505), .B(n_317), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_509), .B(n_395), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
NAND2xp33_ASAP7_75t_SL g573 ( .A(n_512), .B(n_319), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_521), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_521), .Y(n_576) );
OAI222xp33_ASAP7_75t_L g577 ( .A1(n_553), .A2(n_493), .B1(n_495), .B2(n_508), .C1(n_511), .C2(n_479), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_519), .A2(n_495), .B1(n_499), .B2(n_492), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_527), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_529), .B(n_483), .Y(n_580) );
OAI221xp5_ASAP7_75t_SL g581 ( .A1(n_539), .A2(n_492), .B1(n_499), .B2(n_511), .C(n_479), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_517), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_524), .A2(n_483), .B1(n_514), .B2(n_480), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_552), .A2(n_504), .B1(n_490), .B2(n_501), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_556), .A2(n_504), .B1(n_490), .B2(n_501), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_514), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_522), .B(n_483), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_544), .A2(n_494), .B(n_471), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_534), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_546), .B(n_494), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_525), .B(n_471), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_516), .B(n_480), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_561), .A2(n_480), .B(n_473), .C(n_319), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_480), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_544), .A2(n_473), .B(n_191), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_536), .B(n_473), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_560), .A2(n_473), .B(n_321), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_551), .B(n_334), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_546), .B(n_340), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_522), .A2(n_340), .B1(n_334), .B2(n_336), .Y(n_604) );
OAI321xp33_ASAP7_75t_L g605 ( .A1(n_549), .A2(n_362), .A3(n_336), .B1(n_186), .B2(n_322), .C(n_325), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_528), .B(n_334), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_531), .A2(n_227), .B(n_191), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g608 ( .A1(n_531), .A2(n_340), .A3(n_325), .B(n_322), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_537), .A2(n_362), .B1(n_336), .B2(n_328), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_540), .A2(n_362), .B(n_336), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_558), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_559), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_569), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_562), .B(n_56), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_555), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_545), .A2(n_362), .B1(n_336), .B2(n_328), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_531), .A2(n_227), .B(n_188), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_571), .A2(n_228), .B1(n_188), .B2(n_214), .C(n_225), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_518), .A2(n_362), .B1(n_328), .B2(n_327), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_518), .A2(n_328), .B1(n_327), .B2(n_228), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_555), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_542), .A2(n_226), .B(n_214), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_566), .Y(n_625) );
AOI21xp33_ASAP7_75t_SL g626 ( .A1(n_518), .A2(n_59), .B(n_60), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_570), .A2(n_328), .B1(n_327), .B2(n_226), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_575), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_616), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_622), .B(n_550), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_582), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_600), .B(n_540), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_593), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_579), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_583), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_624), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_625), .B(n_526), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_589), .B(n_547), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_576), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_585), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_611), .A2(n_560), .B(n_557), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_594), .B(n_565), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_574), .B(n_538), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_595), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_610), .B(n_548), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_614), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_612), .B(n_541), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_598), .B(n_564), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_613), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_603), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_626), .A2(n_557), .B(n_573), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_603), .Y(n_657) );
INVxp33_ASAP7_75t_L g658 ( .A(n_580), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_596), .B(n_543), .Y(n_659) );
NOR4xp25_ASAP7_75t_SL g660 ( .A(n_581), .B(n_573), .C(n_565), .D(n_564), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_591), .B(n_568), .Y(n_661) );
NOR3xp33_ASAP7_75t_SL g662 ( .A(n_577), .B(n_563), .C(n_63), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_608), .B(n_568), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_591), .B(n_567), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_586), .B(n_599), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_663), .B(n_578), .C(n_590), .D(n_604), .Y(n_668) );
NAND3x2_ASAP7_75t_L g669 ( .A(n_651), .B(n_606), .C(n_623), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_651), .A2(n_642), .B1(n_666), .B2(n_662), .C(n_640), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_643), .A2(n_617), .B(n_623), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_635), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_635), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_633), .B(n_520), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_639), .B(n_520), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_647), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_650), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_632), .A2(n_615), .B1(n_621), .B2(n_620), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_658), .A2(n_567), .B1(n_607), .B2(n_618), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_633), .B(n_601), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_656), .B(n_619), .C(n_605), .Y(n_681) );
AOI32xp33_ASAP7_75t_L g682 ( .A1(n_632), .A2(n_617), .A3(n_609), .B1(n_597), .B2(n_627), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_638), .A2(n_234), .B(n_239), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_644), .Y(n_684) );
AOI322xp5_ASAP7_75t_L g685 ( .A1(n_639), .A2(n_186), .A3(n_64), .B1(n_65), .B2(n_66), .C1(n_69), .C2(n_71), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_644), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_648), .Y(n_687) );
AOI221x1_ASAP7_75t_L g688 ( .A1(n_629), .A2(n_186), .B1(n_327), .B2(n_76), .C(n_77), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_632), .A2(n_655), .B1(n_665), .B2(n_657), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_670), .A2(n_634), .B1(n_655), .B2(n_630), .C(n_659), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_672), .B(n_634), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_677), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_669), .A2(n_660), .B1(n_653), .B2(n_647), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_680), .Y(n_694) );
AO22x2_ASAP7_75t_L g695 ( .A1(n_673), .A2(n_628), .B1(n_631), .B2(n_646), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_676), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_689), .B(n_665), .Y(n_697) );
NAND2x1p5_ASAP7_75t_L g698 ( .A(n_684), .B(n_653), .Y(n_698) );
NOR2xp33_ASAP7_75t_R g699 ( .A(n_679), .B(n_645), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_686), .A2(n_661), .B1(n_648), .B2(n_654), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_667), .B(n_652), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_671), .A2(n_664), .B(n_649), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_668), .A2(n_654), .B1(n_641), .B2(n_636), .C(n_637), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_683), .A2(n_641), .B1(n_636), .B2(n_637), .Y(n_704) );
AOI321xp33_ASAP7_75t_L g705 ( .A1(n_681), .A2(n_61), .A3(n_74), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_679), .A2(n_327), .B1(n_186), .B2(n_239), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_681), .A2(n_239), .B1(n_687), .B2(n_675), .C(n_674), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_682), .A2(n_239), .B(n_678), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_685), .B(n_239), .C(n_688), .D(n_675), .Y(n_709) );
AO22x2_ASAP7_75t_L g710 ( .A1(n_677), .A2(n_640), .B1(n_672), .B2(n_684), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_710), .A2(n_690), .B1(n_692), .B2(n_695), .Y(n_711) );
OR3x2_ASAP7_75t_L g712 ( .A(n_709), .B(n_708), .C(n_694), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_696), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_691), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_698), .B(n_693), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_703), .B1(n_701), .B2(n_696), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_712), .A2(n_695), .B1(n_707), .B2(n_697), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_711), .A2(n_704), .B1(n_702), .B2(n_705), .C(n_700), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_717), .A2(n_711), .B1(n_714), .B2(n_713), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
BUFx3_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_719), .B1(n_716), .B2(n_699), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_721), .B(n_706), .Y(n_723) );
endmodule