module fake_jpeg_12005_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_18),
.Y(n_38)
);

A2O1A1O1Ixp25_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_17),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_67)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_19),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_27),
.B1(n_13),
.B2(n_14),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_13),
.B1(n_21),
.B2(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_34),
.B1(n_37),
.B2(n_21),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_63),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_31),
.B(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_16),
.B1(n_22),
.B2(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_67),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_16),
.B(n_22),
.C(n_20),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_47),
.C(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_0),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_40),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_40),
.Y(n_72)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_78),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_85),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_45),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_82),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_39),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_67),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_70),
.B(n_65),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_86),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_83),
.C(n_72),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_109),
.C(n_39),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_108),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_57),
.Y(n_118)
);

OAI322xp33_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_70),
.A3(n_62),
.B1(n_58),
.B2(n_63),
.C1(n_86),
.C2(n_59),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_90),
.C(n_93),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_62),
.C(n_86),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_89),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_95),
.B1(n_109),
.B2(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_96),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_92),
.C(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.C(n_119),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_104),
.B(n_102),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_116),
.B(n_91),
.Y(n_127)
);

AOI21x1_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_3),
.B(n_4),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_52),
.C(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

NAND4xp25_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_52),
.C(n_118),
.D(n_4),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

OA21x2_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_8),
.B(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_133),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_123),
.B(n_10),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_8),
.B(n_11),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_134),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.Y(n_140)
);


endmodule