module real_aes_78_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_0), .B(n_203), .Y(n_244) );
INVx1_ASAP7_75t_L g541 ( .A(n_0), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_1), .A2(n_215), .B(n_294), .Y(n_293) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_2), .A2(n_51), .B1(n_94), .B2(n_98), .Y(n_97) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_3), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_3), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_3), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g190 ( .A(n_4), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_5), .B(n_224), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_6), .A2(n_23), .B1(n_122), .B2(n_126), .Y(n_121) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_7), .A2(n_21), .B1(n_94), .B2(n_95), .Y(n_93) );
NAND2xp33_ASAP7_75t_L g287 ( .A(n_8), .B(n_222), .Y(n_287) );
INVx2_ASAP7_75t_L g213 ( .A(n_9), .Y(n_213) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_18), .B1(n_203), .B2(n_215), .C(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_11), .B(n_203), .Y(n_283) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_12), .A2(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_13), .B(n_229), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_14), .A2(n_49), .B1(n_155), .B2(n_158), .Y(n_154) );
INVx1_ASAP7_75t_L g169 ( .A(n_15), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_15), .B(n_224), .Y(n_275) );
AO21x1_ASAP7_75t_L g202 ( .A1(n_16), .A2(n_203), .B(n_210), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_17), .A2(n_165), .B1(n_172), .B2(n_173), .Y(n_164) );
INVx1_ASAP7_75t_SL g172 ( .A(n_17), .Y(n_172) );
NAND2x1_ASAP7_75t_L g242 ( .A(n_19), .B(n_224), .Y(n_242) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_19), .A2(n_83), .B1(n_84), .B2(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_19), .Y(n_521) );
NAND2x1_ASAP7_75t_L g301 ( .A(n_20), .B(n_222), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g182 ( .A1(n_21), .A2(n_51), .B1(n_57), .B2(n_183), .C(n_185), .Y(n_182) );
OR2x2_ASAP7_75t_L g212 ( .A(n_22), .B(n_66), .Y(n_212) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_22), .A2(n_66), .B(n_213), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_24), .A2(n_40), .B1(n_130), .B2(n_132), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_25), .B(n_222), .Y(n_296) );
INVx3_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_27), .A2(n_56), .B1(n_142), .B2(n_144), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_28), .B(n_224), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_29), .A2(n_48), .B1(n_149), .B2(n_151), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_30), .B(n_222), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_31), .A2(n_215), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_SL g103 ( .A(n_32), .Y(n_103) );
INVx1_ASAP7_75t_L g192 ( .A(n_33), .Y(n_192) );
AND2x2_ASAP7_75t_L g209 ( .A(n_33), .B(n_190), .Y(n_209) );
AND2x2_ASAP7_75t_L g216 ( .A(n_33), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_34), .B(n_203), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_35), .A2(n_65), .B1(n_113), .B2(n_116), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_36), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_37), .B(n_222), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_38), .A2(n_215), .B(n_300), .Y(n_299) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_39), .A2(n_57), .B1(n_94), .B2(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_41), .B(n_222), .Y(n_243) );
INVx1_ASAP7_75t_L g206 ( .A(n_42), .Y(n_206) );
INVx1_ASAP7_75t_L g219 ( .A(n_42), .Y(n_219) );
INVx1_ASAP7_75t_L g104 ( .A(n_43), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_224), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_45), .A2(n_215), .B(n_241), .Y(n_240) );
AO21x1_ASAP7_75t_L g214 ( .A1(n_46), .A2(n_215), .B(n_220), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_47), .B(n_203), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_50), .B(n_203), .Y(n_303) );
INVxp33_ASAP7_75t_L g187 ( .A(n_51), .Y(n_187) );
AND2x2_ASAP7_75t_L g259 ( .A(n_52), .B(n_230), .Y(n_259) );
INVx1_ASAP7_75t_L g208 ( .A(n_53), .Y(n_208) );
INVx1_ASAP7_75t_L g217 ( .A(n_53), .Y(n_217) );
AND2x2_ASAP7_75t_L g305 ( .A(n_54), .B(n_246), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_55), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_55), .Y(n_176) );
INVxp67_ASAP7_75t_L g186 ( .A(n_57), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_58), .B(n_203), .Y(n_277) );
AND2x2_ASAP7_75t_L g290 ( .A(n_59), .B(n_246), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_60), .A2(n_166), .B1(n_167), .B2(n_171), .Y(n_165) );
INVx1_ASAP7_75t_L g171 ( .A(n_60), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_61), .A2(n_63), .B1(n_88), .B2(n_108), .Y(n_87) );
AND2x2_ASAP7_75t_L g210 ( .A(n_62), .B(n_211), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_64), .A2(n_83), .B1(n_84), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_64), .Y(n_530) );
AND2x2_ASAP7_75t_L g249 ( .A(n_67), .B(n_246), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_68), .B(n_222), .Y(n_276) );
INVx1_ASAP7_75t_L g82 ( .A(n_69), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_70), .B(n_224), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_71), .B(n_222), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_72), .A2(n_215), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_73), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_74), .B(n_224), .Y(n_295) );
BUFx2_ASAP7_75t_L g178 ( .A(n_75), .Y(n_178) );
BUFx2_ASAP7_75t_SL g184 ( .A(n_76), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_77), .A2(n_215), .B(n_285), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_179), .B1(n_193), .B2(n_518), .C(n_519), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_162), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NOR2xp67_ASAP7_75t_L g85 ( .A(n_86), .B(n_135), .Y(n_85) );
NAND4xp25_ASAP7_75t_L g86 ( .A(n_87), .B(n_112), .C(n_121), .D(n_129), .Y(n_86) );
INVx2_ASAP7_75t_SL g88 ( .A(n_89), .Y(n_88) );
INVx8_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x4_ASAP7_75t_L g90 ( .A(n_91), .B(n_99), .Y(n_90) );
AND2x2_ASAP7_75t_L g114 ( .A(n_91), .B(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g124 ( .A(n_91), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g139 ( .A(n_91), .B(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g91 ( .A(n_92), .B(n_96), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x4_ASAP7_75t_L g111 ( .A(n_93), .B(n_96), .Y(n_111) );
INVx1_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
AND2x2_ASAP7_75t_L g128 ( .A(n_93), .B(n_97), .Y(n_128) );
INVx2_ASAP7_75t_L g95 ( .A(n_94), .Y(n_95) );
INVx1_ASAP7_75t_L g98 ( .A(n_94), .Y(n_98) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_94), .A2(n_102), .B1(n_103), .B2(n_104), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_94), .Y(n_102) );
INVx1_ASAP7_75t_L g107 ( .A(n_94), .Y(n_107) );
INVxp67_ASAP7_75t_L g147 ( .A(n_96), .Y(n_147) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g119 ( .A(n_97), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g118 ( .A(n_99), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g127 ( .A(n_99), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_105), .Y(n_99) );
AND2x2_ASAP7_75t_L g115 ( .A(n_100), .B(n_106), .Y(n_115) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g125 ( .A(n_101), .B(n_105), .Y(n_125) );
AND2x2_ASAP7_75t_L g140 ( .A(n_101), .B(n_106), .Y(n_140) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_101), .Y(n_153) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g143 ( .A(n_111), .B(n_115), .Y(n_143) );
AND2x2_ASAP7_75t_L g150 ( .A(n_111), .B(n_125), .Y(n_150) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g131 ( .A(n_115), .B(n_119), .Y(n_131) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx8_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g157 ( .A(n_119), .B(n_125), .Y(n_157) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx6_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g133 ( .A(n_128), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g152 ( .A(n_128), .B(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND4xp25_ASAP7_75t_SL g135 ( .A(n_136), .B(n_141), .C(n_148), .D(n_154), .Y(n_135) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx6_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g146 ( .A(n_140), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g159 ( .A(n_140), .B(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx12f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B1(n_174), .B2(n_175), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
AND3x1_ASAP7_75t_SL g181 ( .A(n_182), .B(n_188), .C(n_191), .Y(n_181) );
INVxp67_ASAP7_75t_L g527 ( .A(n_182), .Y(n_527) );
CKINVDCx8_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_188), .Y(n_525) );
AO21x1_ASAP7_75t_SL g534 ( .A1(n_188), .A2(n_535), .B(n_539), .Y(n_534) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_SL g533 ( .A(n_189), .B(n_191), .Y(n_533) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g218 ( .A(n_190), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_191), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2x1p5_ASAP7_75t_L g536 ( .A(n_192), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_417), .Y(n_194) );
NOR3xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_354), .C(n_377), .Y(n_195) );
NAND3xp33_ASAP7_75t_SL g196 ( .A(n_197), .B(n_306), .C(n_323), .Y(n_196) );
OAI31xp33_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_236), .A3(n_260), .B(n_267), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_198), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_228), .Y(n_199) );
AND2x4_ASAP7_75t_L g309 ( .A(n_200), .B(n_228), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_200), .B(n_251), .Y(n_338) );
AND2x4_ASAP7_75t_L g340 ( .A(n_200), .B(n_334), .Y(n_340) );
AND2x2_ASAP7_75t_L g471 ( .A(n_200), .B(n_264), .Y(n_471) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g316 ( .A(n_201), .Y(n_316) );
OAI21x1_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_214), .B(n_226), .Y(n_201) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_203), .Y(n_518) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_209), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
AND2x6_ASAP7_75t_L g222 ( .A(n_205), .B(n_217), .Y(n_222) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_L g224 ( .A(n_207), .B(n_219), .Y(n_224) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx5_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
INVx1_ASAP7_75t_L g227 ( .A(n_210), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_211), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_SL g271 ( .A(n_211), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_211), .A2(n_283), .B(n_284), .Y(n_282) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_212), .B(n_213), .Y(n_230) );
AND2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g538 ( .A(n_217), .Y(n_538) );
INVx2_ASAP7_75t_L g540 ( .A(n_219), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_223), .B(n_225), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_225), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_225), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_256), .B(n_257), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_225), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_225), .A2(n_286), .B(n_287), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_225), .A2(n_295), .B(n_296), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_225), .A2(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g250 ( .A(n_228), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_228), .B(n_315), .Y(n_407) );
AND2x2_ASAP7_75t_L g413 ( .A(n_228), .B(n_252), .Y(n_413) );
AND2x2_ASAP7_75t_L g502 ( .A(n_228), .B(n_503), .Y(n_502) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_231), .B(n_235), .Y(n_228) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_231), .B(n_235), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_229), .A2(n_292), .B(n_293), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_229), .Y(n_304) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_SL g484 ( .A(n_236), .Y(n_484) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
BUFx2_ASAP7_75t_L g313 ( .A(n_237), .Y(n_313) );
AND2x2_ASAP7_75t_L g347 ( .A(n_237), .B(n_251), .Y(n_347) );
AND2x2_ASAP7_75t_L g396 ( .A(n_237), .B(n_252), .Y(n_396) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g353 ( .A(n_238), .B(n_252), .Y(n_353) );
INVxp67_ASAP7_75t_L g365 ( .A(n_238), .Y(n_365) );
BUFx3_ASAP7_75t_L g410 ( .A(n_238), .Y(n_410) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_245), .B(n_249), .Y(n_238) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_245), .B(n_249), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_244), .Y(n_239) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_245), .A2(n_253), .B(n_259), .Y(n_252) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_253), .B(n_259), .Y(n_266) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx4f_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
OAI31xp33_ASAP7_75t_L g306 ( .A1(n_250), .A2(n_307), .A3(n_312), .B(n_317), .Y(n_306) );
AND2x2_ASAP7_75t_L g314 ( .A(n_251), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g333 ( .A(n_252), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_254), .B(n_258), .Y(n_253) );
AOI322xp5_ASAP7_75t_L g507 ( .A1(n_260), .A2(n_382), .A3(n_411), .B1(n_416), .B2(n_508), .C1(n_511), .C2(n_512), .Y(n_507) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_261), .B(n_353), .Y(n_358) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_261), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g439 ( .A(n_261), .B(n_343), .Y(n_439) );
INVx1_ASAP7_75t_SL g453 ( .A(n_261), .Y(n_453) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_262), .Y(n_477) );
AND2x2_ASAP7_75t_L g406 ( .A(n_263), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_263), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_SL g263 ( .A(n_264), .B(n_265), .Y(n_263) );
BUFx2_ASAP7_75t_L g311 ( .A(n_264), .Y(n_311) );
INVx1_ASAP7_75t_L g503 ( .A(n_264), .Y(n_503) );
OR2x2_ASAP7_75t_L g370 ( .A(n_265), .B(n_315), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_265), .B(n_340), .Y(n_404) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g343 ( .A(n_266), .B(n_315), .Y(n_343) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_288), .Y(n_267) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g399 ( .A(n_269), .Y(n_399) );
OR2x2_ASAP7_75t_L g426 ( .A(n_269), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_280), .Y(n_269) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_270), .B(n_289), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_270), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g499 ( .A(n_270), .B(n_361), .Y(n_499) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_278), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_271), .B(n_279), .Y(n_278) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_271), .A2(n_272), .B(n_278), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
OR2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
INVx2_ASAP7_75t_L g361 ( .A(n_280), .Y(n_361) );
INVx1_ASAP7_75t_L g402 ( .A(n_280), .Y(n_402) );
AND2x2_ASAP7_75t_L g433 ( .A(n_280), .B(n_289), .Y(n_433) );
AND2x2_ASAP7_75t_L g464 ( .A(n_280), .B(n_391), .Y(n_464) );
AND2x2_ASAP7_75t_L g360 ( .A(n_288), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_288), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_288), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g468 ( .A(n_288), .B(n_330), .Y(n_468) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_297), .Y(n_288) );
INVx5_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_289), .B(n_322), .Y(n_400) );
BUFx2_ASAP7_75t_L g460 ( .A(n_289), .Y(n_460) );
OR2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx4_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
AND2x2_ASAP7_75t_L g445 ( .A(n_297), .B(n_328), .Y(n_445) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B(n_305), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_308), .A2(n_435), .B1(n_438), .B2(n_440), .C(n_441), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g456 ( .A(n_309), .B(n_347), .Y(n_456) );
INVx1_ASAP7_75t_SL g482 ( .A(n_309), .Y(n_482) );
AND2x2_ASAP7_75t_L g467 ( .A(n_310), .B(n_439), .Y(n_467) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_311), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g336 ( .A(n_313), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g342 ( .A(n_313), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
AND2x2_ASAP7_75t_L g424 ( .A(n_314), .B(n_352), .Y(n_424) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g345 ( .A(n_321), .Y(n_345) );
OR2x2_ASAP7_75t_L g513 ( .A(n_321), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g329 ( .A(n_322), .Y(n_329) );
AND2x4_ASAP7_75t_L g385 ( .A(n_322), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_322), .B(n_390), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_322), .B(n_328), .Y(n_427) );
AND2x2_ASAP7_75t_L g487 ( .A(n_322), .B(n_390), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_331), .B1(n_344), .B2(n_346), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_324), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND3x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .C(n_330), .Y(n_326) );
AND2x4_ASAP7_75t_L g344 ( .A(n_327), .B(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_328), .B(n_385), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_329), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g429 ( .A(n_330), .Y(n_429) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_330), .A2(n_459), .A3(n_495), .B1(n_497), .B2(n_500), .C1(n_504), .C2(n_505), .Y(n_494) );
NAND4xp25_ASAP7_75t_SL g331 ( .A(n_332), .B(n_335), .C(n_339), .D(n_341), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_333), .B(n_349), .Y(n_461) );
BUFx2_ASAP7_75t_L g352 ( .A(n_334), .Y(n_352) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g476 ( .A(n_337), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g490 ( .A(n_338), .B(n_365), .Y(n_490) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g356 ( .A(n_340), .B(n_357), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_340), .A2(n_409), .B(n_411), .C(n_414), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_340), .B(n_347), .Y(n_466) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_342), .A2(n_424), .B1(n_425), .B2(n_428), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_379), .B1(n_383), .B2(n_387), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_343), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_343), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_343), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g510 ( .A(n_343), .Y(n_510) );
INVx1_ASAP7_75t_L g449 ( .A(n_344), .Y(n_449) );
OAI21xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_348), .B(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g357 ( .A(n_347), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_347), .B(n_352), .Y(n_506) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g442 ( .A(n_349), .B(n_353), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_351), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g509 ( .A(n_352), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g483 ( .A(n_353), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_359), .C(n_362), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp33_ASAP7_75t_SL g469 ( .A1(n_357), .A2(n_388), .B1(n_435), .B2(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_361), .B(n_384), .Y(n_392) );
OR2x2_ASAP7_75t_L g421 ( .A(n_361), .B(n_422), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_367), .B(n_371), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI211xp5_ASAP7_75t_SL g420 ( .A1(n_368), .A2(n_421), .B(n_423), .C(n_431), .Y(n_420) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp67_ASAP7_75t_SL g454 ( .A(n_373), .B(n_400), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_373), .Y(n_457) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_375), .B(n_384), .Y(n_514) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g386 ( .A(n_376), .Y(n_386) );
INVx2_ASAP7_75t_L g391 ( .A(n_376), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_393), .C(n_405), .D(n_408), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_381), .A2(n_513), .B1(n_515), .B2(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x4_ASAP7_75t_L g480 ( .A(n_384), .B(n_410), .Y(n_480) );
AND2x2_ASAP7_75t_L g401 ( .A(n_385), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_385), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
INVx1_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .A3(n_400), .B1(n_401), .B2(n_403), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_394), .A2(n_442), .B(n_443), .Y(n_441) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_397), .A2(n_474), .B1(n_476), .B2(n_478), .C(n_481), .Y(n_473) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g458 ( .A(n_399), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g416 ( .A(n_400), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_401), .A2(n_439), .B1(n_489), .B2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g415 ( .A(n_402), .Y(n_415) );
AND2x2_ASAP7_75t_L g493 ( .A(n_402), .B(n_446), .Y(n_493) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_409), .B(n_461), .Y(n_496) );
INVx1_ASAP7_75t_L g515 ( .A(n_409), .Y(n_515) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_418), .B(n_472), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_462), .Y(n_418) );
NOR3xp33_ASAP7_75t_SL g419 ( .A(n_420), .B(n_434), .C(n_447), .Y(n_419) );
INVx1_ASAP7_75t_L g437 ( .A(n_422), .Y(n_437) );
INVx1_ASAP7_75t_SL g448 ( .A(n_424), .Y(n_448) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g430 ( .A(n_427), .Y(n_430) );
INVx2_ASAP7_75t_L g440 ( .A(n_428), .Y(n_440) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AND2x4_ASAP7_75t_L g486 ( .A(n_429), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g504 ( .A(n_433), .B(n_487), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
AOI32xp33_ASAP7_75t_L g455 ( .A1(n_444), .A2(n_456), .A3(n_457), .B1(n_458), .B2(n_461), .Y(n_455) );
NOR2xp33_ASAP7_75t_SL g474 ( .A(n_444), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g475 ( .A(n_446), .Y(n_475) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B(n_450), .C(n_455), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g511 ( .A(n_459), .B(n_499), .Y(n_511) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_460), .B(n_499), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_467), .B2(n_468), .C(n_469), .Y(n_462) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_473), .B(n_488), .C(n_494), .D(n_507), .Y(n_472) );
INVxp33_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .C(n_485), .Y(n_481) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OAI222xp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_528), .B2(n_531), .C1(n_534), .C2(n_541), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
endmodule