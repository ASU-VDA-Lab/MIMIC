module real_aes_7791_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_1170;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_792;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_1200;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_1113;
wire n_766;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_1034;
wire n_491;
wire n_694;
wire n_923;
wire n_894;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_1140;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_994;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_1199;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_1053;
wire n_559;
wire n_1182;
wire n_636;
wire n_976;
wire n_906;
wire n_477;
wire n_872;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_656;
wire n_1025;
wire n_532;
wire n_746;
wire n_1168;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1135;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_1174;
wire n_1167;
wire n_1193;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_449;
wire n_1006;
wire n_417;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_1198;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_1103;
wire n_880;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_1145;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_1179;
wire n_1201;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1105;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_1187;
wire n_727;
wire n_1014;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_899;
wire n_526;
wire n_928;
wire n_637;
wire n_653;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_1162;
wire n_861;
wire n_705;
wire n_1191;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_1172;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_1190;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_1114;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_474;
wire n_1159;
wire n_1156;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_652;
wire n_703;
wire n_500;
wire n_1101;
wire n_1102;
wire n_601;
wire n_463;
wire n_661;
wire n_1076;
wire n_804;
wire n_447;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_0), .Y(n_1189) );
INVx1_ASAP7_75t_L g780 ( .A(n_1), .Y(n_780) );
AOI222xp33_ASAP7_75t_L g519 ( .A1(n_2), .A2(n_195), .B1(n_351), .B2(n_492), .C1(n_520), .C2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_3), .A2(n_108), .B1(n_930), .B2(n_1019), .Y(n_1056) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_4), .A2(n_344), .B1(n_930), .B2(n_990), .C(n_991), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g1144 ( .A(n_5), .Y(n_1144) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_6), .A2(n_177), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_7), .A2(n_98), .B1(n_618), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_8), .A2(n_248), .B1(n_550), .B2(n_553), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_9), .B(n_672), .Y(n_671) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_10), .A2(n_236), .B1(n_423), .B2(n_428), .Y(n_431) );
INVx1_ASAP7_75t_L g1136 ( .A(n_10), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_11), .A2(n_188), .B1(n_419), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_12), .A2(n_375), .B1(n_486), .B2(n_517), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_13), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_14), .A2(n_172), .B1(n_533), .B2(n_735), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1105 ( .A(n_15), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g1116 ( .A(n_16), .Y(n_1116) );
INVx1_ASAP7_75t_L g855 ( .A(n_17), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_18), .A2(n_263), .B1(n_474), .B2(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_19), .A2(n_111), .B1(n_654), .B2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_20), .A2(n_143), .B1(n_434), .B2(n_439), .Y(n_1193) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_21), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_22), .A2(n_336), .B1(n_654), .B2(n_1024), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_23), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_24), .A2(n_337), .B1(n_609), .B2(n_1146), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_25), .A2(n_325), .B1(n_717), .B2(n_990), .Y(n_1084) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_26), .A2(n_69), .B1(n_297), .B2(n_483), .C1(n_486), .C2(n_490), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_27), .A2(n_324), .B1(n_509), .B2(n_1027), .Y(n_1026) );
AOI22xp5_ASAP7_75t_SL g728 ( .A1(n_28), .A2(n_260), .B1(n_533), .B2(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_29), .Y(n_1034) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_30), .A2(n_38), .B1(n_457), .B2(n_797), .C(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_31), .A2(n_322), .B1(n_717), .B2(n_1019), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_32), .A2(n_382), .B1(n_477), .B2(n_678), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_33), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_34), .Y(n_1100) );
AO22x2_ASAP7_75t_L g433 ( .A1(n_35), .A2(n_127), .B1(n_423), .B2(n_424), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_36), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_37), .A2(n_58), .B1(n_538), .B2(n_618), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_39), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_40), .Y(n_1190) );
INVx1_ASAP7_75t_L g758 ( .A(n_41), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_42), .A2(n_66), .B1(n_449), .B2(n_500), .Y(n_884) );
INVx1_ASAP7_75t_L g832 ( .A(n_43), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_44), .A2(n_182), .B1(n_419), .B2(n_614), .Y(n_968) );
INVx1_ASAP7_75t_L g994 ( .A(n_45), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_46), .A2(n_194), .B1(n_656), .B2(n_874), .Y(n_1198) );
INVx1_ASAP7_75t_L g964 ( .A(n_47), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_48), .B(n_792), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_49), .A2(n_225), .B1(n_466), .B2(n_493), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g1000 ( .A1(n_50), .A2(n_148), .B1(n_157), .B2(n_520), .C1(n_600), .C2(n_701), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_51), .A2(n_89), .B1(n_608), .B2(n_1195), .Y(n_1194) );
AOI22xp5_ASAP7_75t_SL g726 ( .A1(n_52), .A2(n_332), .B1(n_439), .B2(n_727), .Y(n_726) );
AOI222xp33_ASAP7_75t_L g1068 ( .A1(n_53), .A2(n_313), .B1(n_335), .B2(n_570), .C1(n_704), .C2(n_917), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_54), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_55), .A2(n_128), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI22xp5_ASAP7_75t_SL g883 ( .A1(n_56), .A2(n_235), .B1(n_727), .B2(n_735), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_57), .A2(n_78), .B1(n_701), .B2(n_792), .Y(n_1010) );
INVx1_ASAP7_75t_L g862 ( .A(n_59), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_60), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_61), .A2(n_193), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_62), .A2(n_345), .B1(n_460), .B2(n_465), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_63), .A2(n_316), .B1(n_564), .B2(n_566), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g1096 ( .A(n_64), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_65), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_67), .B(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_68), .A2(n_259), .B1(n_550), .B2(n_553), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_70), .A2(n_287), .B1(n_518), .B2(n_792), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_71), .A2(n_380), .B1(n_870), .B2(n_871), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_72), .A2(n_97), .B1(n_465), .B2(n_492), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_73), .A2(n_138), .B1(n_471), .B2(n_544), .Y(n_675) );
INVx1_ASAP7_75t_L g777 ( .A(n_74), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_75), .A2(n_160), .B1(n_509), .B2(n_612), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_76), .A2(n_215), .B1(n_509), .B2(n_536), .Y(n_1197) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_77), .B(n_733), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_79), .A2(n_232), .B1(n_458), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_80), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_81), .A2(n_245), .B1(n_536), .B2(n_605), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_82), .A2(n_1140), .B1(n_1163), .B2(n_1164), .Y(n_1139) );
CKINVDCx20_ASAP7_75t_R g1163 ( .A(n_82), .Y(n_1163) );
INVx1_ASAP7_75t_L g859 ( .A(n_83), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_84), .A2(n_102), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_85), .A2(n_243), .B1(n_447), .B2(n_806), .Y(n_805) );
AOI22xp5_ASAP7_75t_SL g886 ( .A1(n_86), .A2(n_103), .B1(n_618), .B2(n_806), .Y(n_886) );
INVx1_ASAP7_75t_L g841 ( .A(n_87), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_88), .A2(n_164), .B1(n_612), .B2(n_615), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_90), .A2(n_171), .B1(n_553), .B2(n_826), .Y(n_825) );
AO22x2_ASAP7_75t_L g427 ( .A1(n_91), .A2(n_272), .B1(n_423), .B2(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g1133 ( .A(n_91), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_92), .A2(n_286), .B1(n_477), .B2(n_480), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_93), .A2(n_371), .B1(n_490), .B2(n_836), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_94), .A2(n_369), .B1(n_434), .B2(n_614), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_95), .A2(n_387), .B1(n_608), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g1009 ( .A(n_96), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_99), .A2(n_305), .B1(n_609), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_100), .A2(n_327), .B1(n_500), .B2(n_544), .Y(n_1045) );
OA22x2_ASAP7_75t_L g1052 ( .A1(n_101), .A2(n_1053), .B1(n_1054), .B2(n_1069), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_101), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_104), .A2(n_221), .B1(n_733), .B2(n_819), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_105), .A2(n_121), .B1(n_471), .B2(n_618), .Y(n_969) );
INVx1_ASAP7_75t_L g830 ( .A(n_106), .Y(n_830) );
INVx1_ASAP7_75t_L g880 ( .A(n_107), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_109), .A2(n_251), .B1(n_826), .B2(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g815 ( .A(n_110), .Y(n_815) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_112), .A2(n_174), .B1(n_566), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_113), .A2(n_227), .B1(n_797), .B2(n_1013), .Y(n_1082) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_114), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_115), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_116), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_117), .B(n_960), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_118), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_119), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_120), .A2(n_256), .B1(n_477), .B2(n_874), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g949 ( .A1(n_122), .A2(n_296), .B1(n_447), .B2(n_727), .Y(n_949) );
INVx1_ASAP7_75t_L g821 ( .A(n_123), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_124), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_125), .Y(n_1091) );
INVx1_ASAP7_75t_L g945 ( .A(n_126), .Y(n_945) );
INVx1_ASAP7_75t_L g1137 ( .A(n_127), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_129), .A2(n_156), .B1(n_609), .B2(n_1022), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_130), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g1181 ( .A(n_131), .Y(n_1181) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_132), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g1158 ( .A(n_133), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_134), .A2(n_216), .B1(n_461), .B2(n_864), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_135), .A2(n_142), .B1(n_819), .B2(n_928), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_136), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_137), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_139), .A2(n_220), .B1(n_536), .B2(n_605), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_140), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_141), .A2(n_273), .B1(n_564), .B2(n_566), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g1154 ( .A(n_144), .Y(n_1154) );
AOI211xp5_ASAP7_75t_L g1098 ( .A1(n_145), .A2(n_917), .B(n_1099), .C(n_1103), .Y(n_1098) );
INVx1_ASAP7_75t_L g954 ( .A(n_146), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_147), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_149), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_150), .Y(n_534) );
INVx1_ASAP7_75t_L g973 ( .A(n_151), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_152), .A2(n_355), .B1(n_953), .B2(n_1062), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_153), .A2(n_270), .B1(n_518), .B2(n_792), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g1085 ( .A1(n_154), .A2(n_234), .B1(n_434), .B2(n_1086), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_155), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_158), .A2(n_378), .B1(n_486), .B2(n_517), .Y(n_962) );
AOI211xp5_ASAP7_75t_L g1087 ( .A1(n_159), .A2(n_870), .B(n_1088), .C(n_1092), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_161), .A2(n_811), .B1(n_845), .B2(n_846), .Y(n_810) );
CKINVDCx16_ASAP7_75t_R g845 ( .A(n_161), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g1155 ( .A(n_162), .Y(n_1155) );
CKINVDCx20_ASAP7_75t_R g1173 ( .A(n_163), .Y(n_1173) );
OAI22xp5_ASAP7_75t_SL g1176 ( .A1(n_163), .A2(n_1173), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_165), .A2(n_279), .B1(n_615), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_166), .A2(n_203), .B1(n_480), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_167), .A2(n_377), .B1(n_566), .B2(n_795), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_168), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_169), .A2(n_290), .B1(n_466), .B2(n_795), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_170), .Y(n_1148) );
AND2x6_ASAP7_75t_L g401 ( .A(n_173), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_173), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_175), .A2(n_320), .B1(n_732), .B2(n_819), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g1077 ( .A(n_176), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_178), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_179), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_180), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_181), .A2(n_271), .B1(n_600), .B2(n_919), .Y(n_918) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_183), .A2(n_373), .B1(n_504), .B2(n_717), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_184), .A2(n_254), .B1(n_466), .B2(n_492), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_185), .A2(n_389), .B1(n_419), .B2(n_618), .Y(n_680) );
AO22x1_ASAP7_75t_L g986 ( .A1(n_186), .A2(n_198), .B1(n_987), .B2(n_988), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_187), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_189), .A2(n_354), .B1(n_439), .B2(n_714), .C(n_986), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_190), .A2(n_284), .B1(n_1022), .B2(n_1058), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_191), .A2(n_396), .B1(n_575), .B2(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g912 ( .A(n_192), .Y(n_912) );
INVx1_ASAP7_75t_L g837 ( .A(n_196), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_197), .Y(n_1150) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_199), .A2(n_204), .B1(n_509), .B2(n_928), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_200), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_201), .A2(n_282), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
AO22x2_ASAP7_75t_L g422 ( .A1(n_202), .A2(n_261), .B1(n_423), .B2(n_424), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g1134 ( .A(n_202), .B(n_1135), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_205), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_206), .A2(n_281), .B1(n_439), .B2(n_533), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_207), .A2(n_264), .B1(n_500), .B2(n_501), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_208), .A2(n_323), .B1(n_791), .B2(n_792), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_209), .A2(n_364), .B1(n_501), .B2(n_735), .Y(n_951) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_210), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_211), .A2(n_353), .B1(n_501), .B2(n_808), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g1182 ( .A(n_212), .Y(n_1182) );
CKINVDCx20_ASAP7_75t_R g1079 ( .A(n_213), .Y(n_1079) );
AOI22xp5_ASAP7_75t_SL g731 ( .A1(n_214), .A2(n_292), .B1(n_732), .B2(n_733), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_217), .A2(n_252), .B1(n_419), .B2(n_434), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_218), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_219), .A2(n_399), .B(n_407), .C(n_1138), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_222), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_223), .B(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g1081 ( .A1(n_224), .A2(n_370), .B1(n_465), .B2(n_795), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_226), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_228), .A2(n_262), .B1(n_566), .B2(n_795), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_229), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_230), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_231), .A2(n_982), .B1(n_983), .B2(n_1001), .Y(n_981) );
INVx1_ASAP7_75t_L g1001 ( .A(n_231), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_233), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_237), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_238), .A2(n_625), .B1(n_659), .B2(n_660), .Y(n_624) );
INVx1_ASAP7_75t_L g659 ( .A(n_238), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g1157 ( .A(n_239), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_240), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_241), .A2(n_253), .B1(n_507), .B2(n_990), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_242), .A2(n_374), .B1(n_953), .B2(n_1062), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_244), .B(n_457), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_246), .A2(n_384), .B1(n_434), .B2(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_247), .Y(n_745) );
XNOR2xp5_ASAP7_75t_L g1005 ( .A(n_249), .B(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_250), .A2(n_288), .B1(n_732), .B2(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g406 ( .A(n_255), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_257), .A2(n_343), .B1(n_486), .B2(n_493), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_258), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_265), .A2(n_278), .B1(n_439), .B2(n_447), .Y(n_438) );
OA22x2_ASAP7_75t_L g849 ( .A1(n_266), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_266), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_267), .A2(n_303), .B1(n_544), .B2(n_721), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_268), .A2(n_526), .B1(n_577), .B2(n_578), .Y(n_525) );
INVx1_ASAP7_75t_L g577 ( .A(n_268), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_269), .A2(n_330), .B1(n_471), .B2(n_474), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_274), .A2(n_329), .B1(n_553), .B2(n_677), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_275), .A2(n_379), .B1(n_808), .B2(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g755 ( .A(n_276), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_277), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g1185 ( .A(n_280), .Y(n_1185) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_283), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_285), .A2(n_368), .B1(n_802), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_289), .A2(n_334), .B1(n_797), .B2(n_1066), .Y(n_1065) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_291), .B(n_457), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_293), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_294), .A2(n_348), .B1(n_538), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_295), .A2(n_383), .B1(n_453), .B2(n_457), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_298), .A2(n_397), .B1(n_714), .B2(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_299), .Y(n_894) );
INVx1_ASAP7_75t_L g423 ( .A(n_300), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_301), .A2(n_307), .B1(n_797), .B2(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g834 ( .A(n_302), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_304), .A2(n_585), .B1(n_619), .B2(n_620), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_304), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_306), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_308), .Y(n_1089) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_309), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_310), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_311), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_312), .A2(n_358), .B1(n_471), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g824 ( .A(n_314), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_315), .Y(n_901) );
INVx1_ASAP7_75t_L g913 ( .A(n_317), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_318), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_319), .A2(n_367), .B1(n_461), .B2(n_465), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_321), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_326), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_328), .A2(n_359), .B1(n_517), .B2(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g1015 ( .A(n_331), .B(n_744), .Y(n_1015) );
AO22x2_ASAP7_75t_L g1030 ( .A1(n_333), .A2(n_1031), .B1(n_1047), .B2(n_1048), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_333), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_338), .Y(n_784) );
INVx1_ASAP7_75t_L g405 ( .A(n_339), .Y(n_405) );
AOI22xp5_ASAP7_75t_SL g908 ( .A1(n_340), .A2(n_909), .B1(n_934), .B2(n_935), .Y(n_908) );
INVx1_ASAP7_75t_L g935 ( .A(n_340), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_341), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g1162 ( .A(n_346), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_347), .B(n_515), .Y(n_961) );
INVx1_ASAP7_75t_L g844 ( .A(n_349), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_350), .B(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g781 ( .A(n_352), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_356), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_357), .B(n_453), .Y(n_1101) );
INVx1_ASAP7_75t_L g865 ( .A(n_360), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_361), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_362), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_363), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_365), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_366), .Y(n_628) );
INVx1_ASAP7_75t_L g1117 ( .A(n_372), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_376), .B(n_515), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_381), .Y(n_1114) );
INVx1_ASAP7_75t_L g857 ( .A(n_385), .Y(n_857) );
INVx1_ASAP7_75t_L g992 ( .A(n_386), .Y(n_992) );
XNOR2xp5_ASAP7_75t_L g1071 ( .A(n_388), .B(n_1072), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_390), .Y(n_601) );
INVx1_ASAP7_75t_L g817 ( .A(n_391), .Y(n_817) );
OA22x2_ASAP7_75t_L g690 ( .A1(n_392), .A2(n_691), .B1(n_692), .B2(n_722), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_392), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_393), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_394), .Y(n_1161) );
CKINVDCx20_ASAP7_75t_R g1159 ( .A(n_395), .Y(n_1159) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_402), .Y(n_1129) );
OA21x2_ASAP7_75t_L g1171 ( .A1(n_403), .A2(n_1128), .B(n_1172), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_684), .B2(n_1124), .C(n_1125), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_580), .B2(n_581), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_525), .B2(n_579), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AO22x1_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_496), .B1(n_523), .B2(n_524), .Y(n_414) );
INVx2_ASAP7_75t_SL g523 ( .A(n_415), .Y(n_523) );
AO22x2_ASAP7_75t_L g662 ( .A1(n_415), .A2(n_523), .B1(n_663), .B2(n_683), .Y(n_662) );
XOR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_495), .Y(n_415) );
NAND4xp75_ASAP7_75t_L g416 ( .A(n_417), .B(n_451), .C(n_469), .D(n_482), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_438), .Y(n_417) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g540 ( .A(n_420), .Y(n_540) );
BUFx3_ASAP7_75t_L g658 ( .A(n_420), .Y(n_658) );
BUFx3_ASAP7_75t_L g735 ( .A(n_420), .Y(n_735) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_429), .Y(n_420) );
AND2x2_ASAP7_75t_L g479 ( .A(n_421), .B(n_450), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_421), .B(n_450), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_421), .B(n_429), .Y(n_778) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_426), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_422), .B(n_427), .Y(n_437) );
INVx2_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
AND2x2_ASAP7_75t_L g464 ( .A(n_422), .B(n_431), .Y(n_464) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_425), .Y(n_428) );
INVx1_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g446 ( .A(n_427), .Y(n_446) );
AND2x2_ASAP7_75t_L g456 ( .A(n_427), .B(n_445), .Y(n_456) );
INVx1_ASAP7_75t_L g489 ( .A(n_427), .Y(n_489) );
AND2x4_ASAP7_75t_L g435 ( .A(n_429), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g473 ( .A(n_429), .B(n_444), .Y(n_473) );
AND2x4_ASAP7_75t_L g475 ( .A(n_429), .B(n_456), .Y(n_475) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
OR2x2_ASAP7_75t_L g443 ( .A(n_430), .B(n_433), .Y(n_443) );
AND2x2_ASAP7_75t_L g450 ( .A(n_430), .B(n_433), .Y(n_450) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g468 ( .A(n_431), .B(n_433), .Y(n_468) );
AND2x2_ASAP7_75t_L g488 ( .A(n_432), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g640 ( .A(n_432), .Y(n_640) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g463 ( .A(n_433), .Y(n_463) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_SL g547 ( .A(n_435), .Y(n_547) );
BUFx3_ASAP7_75t_L g618 ( .A(n_435), .Y(n_618) );
BUFx3_ASAP7_75t_L g732 ( .A(n_435), .Y(n_732) );
INVx1_ASAP7_75t_L g773 ( .A(n_435), .Y(n_773) );
BUFx3_ASAP7_75t_L g871 ( .A(n_435), .Y(n_871) );
BUFx2_ASAP7_75t_SL g926 ( .A(n_435), .Y(n_926) );
BUFx2_ASAP7_75t_L g953 ( .A(n_435), .Y(n_953) );
AND2x2_ASAP7_75t_L g733 ( .A(n_436), .B(n_640), .Y(n_733) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_L g481 ( .A(n_437), .B(n_463), .Y(n_481) );
INVx1_ASAP7_75t_L g1113 ( .A(n_439), .Y(n_1113) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g654 ( .A(n_440), .Y(n_654) );
INVx4_ASAP7_75t_L g806 ( .A(n_440), .Y(n_806) );
OAI221xp5_ASAP7_75t_SL g1142 ( .A1(n_440), .A2(n_1028), .B1(n_1143), .B2(n_1144), .C(n_1145), .Y(n_1142) );
INVx11_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx11_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
AND2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
AND2x4_ASAP7_75t_L g455 ( .A(n_442), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g558 ( .A(n_443), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g449 ( .A(n_444), .B(n_450), .Y(n_449) );
AND2x6_ASAP7_75t_L g485 ( .A(n_444), .B(n_468), .Y(n_485) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
INVx2_ASAP7_75t_L g615 ( .A(n_448), .Y(n_615) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_448), .A2(n_472), .B1(n_768), .B2(n_769), .Y(n_767) );
OAI221xp5_ASAP7_75t_SL g820 ( .A1(n_448), .A2(n_821), .B1(n_822), .B2(n_824), .C(n_825), .Y(n_820) );
INVx2_ASAP7_75t_L g930 ( .A(n_448), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_448), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
INVx6_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g533 ( .A(n_449), .Y(n_533) );
BUFx3_ASAP7_75t_L g717 ( .A(n_449), .Y(n_717) );
BUFx3_ASAP7_75t_L g876 ( .A(n_449), .Y(n_876) );
AND2x6_ASAP7_75t_L g458 ( .A(n_450), .B(n_456), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_450), .B(n_456), .Y(n_513) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_459), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
INVx2_ASAP7_75t_L g672 ( .A(n_454), .Y(n_672) );
INVx5_ASAP7_75t_L g744 ( .A(n_454), .Y(n_744) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g559 ( .A(n_456), .Y(n_559) );
INVx1_ASAP7_75t_L g1014 ( .A(n_457), .Y(n_1014) );
BUFx4f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g799 ( .A(n_458), .Y(n_799) );
BUFx2_ASAP7_75t_L g960 ( .A(n_458), .Y(n_960) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_458), .Y(n_1066) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
INVx1_ASAP7_75t_L g565 ( .A(n_461), .Y(n_565) );
BUFx2_ASAP7_75t_L g795 ( .A(n_461), .Y(n_795) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g487 ( .A(n_464), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g493 ( .A(n_464), .B(n_494), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_464), .B(n_640), .Y(n_639) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
BUFx2_ASAP7_75t_SL g947 ( .A(n_466), .Y(n_947) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g646 ( .A(n_467), .Y(n_646) );
INVx1_ASAP7_75t_L g645 ( .A(n_468), .Y(n_645) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
BUFx2_ASAP7_75t_SL g729 ( .A(n_473), .Y(n_729) );
BUFx2_ASAP7_75t_SL g870 ( .A(n_473), .Y(n_870) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_474), .Y(n_1086) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
BUFx3_ASAP7_75t_L g544 ( .A(n_475), .Y(n_544) );
INVx2_ASAP7_75t_L g606 ( .A(n_475), .Y(n_606) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_475), .Y(n_819) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_477), .Y(n_1146) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx5_ASAP7_75t_L g504 ( .A(n_478), .Y(n_504) );
INVx4_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
INVx1_ASAP7_75t_L g677 ( .A(n_478), .Y(n_677) );
INVx3_ASAP7_75t_L g727 ( .A(n_478), .Y(n_727) );
BUFx3_ASAP7_75t_L g827 ( .A(n_478), .Y(n_827) );
INVx8_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx4f_ASAP7_75t_SL g609 ( .A(n_480), .Y(n_609) );
BUFx2_ASAP7_75t_L g678 ( .A(n_480), .Y(n_678) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_480), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1195 ( .A(n_480), .Y(n_1195) );
INVx6_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_SL g553 ( .A(n_481), .Y(n_553) );
INVx1_ASAP7_75t_L g721 ( .A(n_481), .Y(n_721) );
INVx1_ASAP7_75t_SL g928 ( .A(n_481), .Y(n_928) );
INVx2_ASAP7_75t_L g1184 ( .A(n_483), .Y(n_1184) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g698 ( .A(n_484), .Y(n_698) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_484), .A2(n_899), .B1(n_900), .B2(n_901), .Y(n_898) );
INVx4_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx2_ASAP7_75t_SL g572 ( .A(n_485), .Y(n_572) );
INVx2_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
INVx2_ASAP7_75t_L g739 ( .A(n_485), .Y(n_739) );
BUFx3_ASAP7_75t_L g917 ( .A(n_485), .Y(n_917) );
INVx4_ASAP7_75t_L g631 ( .A(n_486), .Y(n_631) );
BUFx2_ASAP7_75t_L g791 ( .A(n_486), .Y(n_791) );
INVx2_ASAP7_75t_L g900 ( .A(n_486), .Y(n_900) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_487), .Y(n_521) );
BUFx4f_ASAP7_75t_SL g570 ( .A(n_487), .Y(n_570) );
BUFx2_ASAP7_75t_L g836 ( .A(n_487), .Y(n_836) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_487), .Y(n_864) );
INVx1_ASAP7_75t_L g494 ( .A(n_489), .Y(n_494) );
INVx1_ASAP7_75t_L g1106 ( .A(n_490), .Y(n_1106) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx4f_ASAP7_75t_SL g704 ( .A(n_492), .Y(n_704) );
BUFx12f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_493), .Y(n_575) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_493), .Y(n_792) );
INVx2_ASAP7_75t_SL g524 ( .A(n_496), .Y(n_524) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_522), .Y(n_496) );
NAND4xp75_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .C(n_510), .D(n_519), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
INVx5_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g530 ( .A(n_502), .Y(n_530) );
INVx2_ASAP7_75t_SL g614 ( .A(n_502), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_502), .B(n_780), .Y(n_779) );
INVx4_ASAP7_75t_L g1025 ( .A(n_502), .Y(n_1025) );
BUFx2_ASAP7_75t_L g608 ( .A(n_504), .Y(n_608) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_504), .Y(n_651) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
BUFx2_ASAP7_75t_L g987 ( .A(n_509), .Y(n_987) );
OA211x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_514), .C(n_516), .Y(n_510) );
BUFx3_ASAP7_75t_L g561 ( .A(n_512), .Y(n_561) );
INVx2_ASAP7_75t_L g591 ( .A(n_512), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_512), .A2(n_588), .B1(n_628), .B2(n_629), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_512), .A2(n_639), .B1(n_758), .B2(n_759), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_512), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_512), .A2(n_556), .B1(n_912), .B2(n_913), .Y(n_911) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g891 ( .A(n_513), .Y(n_891) );
INVx1_ASAP7_75t_SL g567 ( .A(n_518), .Y(n_567) );
INVx2_ASAP7_75t_SL g633 ( .A(n_520), .Y(n_633) );
INVx2_ASAP7_75t_L g788 ( .A(n_520), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_521), .Y(n_595) );
INVx1_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
INVx1_ASAP7_75t_L g578 ( .A(n_526), .Y(n_578) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_554), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_541), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_531), .B1(n_532), .B2(n_534), .C(n_535), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_537), .Y(n_714) );
INVx3_ASAP7_75t_L g933 ( .A(n_537), .Y(n_933) );
BUFx3_ASAP7_75t_L g1024 ( .A(n_537), .Y(n_1024) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_540), .Y(n_808) );
OAI221xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_545), .B1(n_546), .B2(n_548), .C(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_552), .Y(n_1022) );
NOR2xp33_ASAP7_75t_SL g554 ( .A(n_555), .B(n_568), .Y(n_554) );
OAI221xp5_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_560), .B1(n_561), .B2(n_562), .C(n_563), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_556), .A2(n_590), .B1(n_695), .B2(n_696), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_556), .A2(n_890), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g588 ( .A(n_557), .Y(n_588) );
INVx1_ASAP7_75t_SL g831 ( .A(n_557), .Y(n_831) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_558), .A2(n_755), .B(n_756), .Y(n_754) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_558), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_561), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_854) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B1(n_572), .B2(n_573), .C1(n_574), .C2(n_576), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_572), .A2(n_631), .B1(n_761), .B2(n_762), .Y(n_760) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_574), .A2(n_631), .B1(n_632), .B2(n_633), .C1(n_634), .C2(n_635), .Y(n_630) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx3_ASAP7_75t_L g600 ( .A(n_575), .Y(n_600) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_621), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g620 ( .A(n_585), .Y(n_620) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_602), .Y(n_585) );
NOR2xp33_ASAP7_75t_SL g586 ( .A(n_587), .B(n_594), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_592), .C(n_593), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_588), .A2(n_890), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
OAI211xp5_ASAP7_75t_L g1099 ( .A1(n_590), .A2(n_1100), .B(n_1101), .C(n_1102), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_590), .A2(n_831), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI222xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_598), .C1(n_599), .C2(n_601), .Y(n_594) );
OAI222xp33_ASAP7_75t_L g1156 ( .A1(n_595), .A2(n_599), .B1(n_788), .B2(n_1157), .C1(n_1158), .C2(n_1159), .Y(n_1156) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_597), .A2(n_667), .B(n_668), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g944 ( .A1(n_597), .A2(n_945), .B(n_946), .Y(n_944) );
OAI21xp5_ASAP7_75t_SL g963 ( .A1(n_597), .A2(n_964), .B(n_965), .Y(n_963) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_610), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g764 ( .A1(n_606), .A2(n_765), .B(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g802 ( .A(n_606), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_609), .Y(n_995) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_661), .B2(n_662), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g660 ( .A(n_625), .Y(n_660) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_647), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .C(n_636), .Y(n_626) );
INVx3_ASAP7_75t_L g701 ( .A(n_631), .Y(n_701) );
OAI221xp5_ASAP7_75t_SL g833 ( .A1(n_633), .A2(n_834), .B1(n_835), .B2(n_837), .C(n_838), .Y(n_833) );
OAI21xp33_ASAP7_75t_L g858 ( .A1(n_633), .A2(n_859), .B(n_860), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_641), .B2(n_642), .Y(n_636) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx3_ASAP7_75t_L g707 ( .A(n_639), .Y(n_707) );
INVx4_ASAP7_75t_L g843 ( .A(n_639), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_639), .A2(n_862), .B1(n_863), .B2(n_865), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_639), .A2(n_642), .B1(n_998), .B2(n_999), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_642), .A2(n_841), .B1(n_842), .B2(n_844), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_642), .A2(n_707), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_642), .A2(n_707), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g923 ( .A(n_643), .Y(n_923) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g709 ( .A(n_644), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_644), .A2(n_842), .B1(n_1040), .B2(n_1041), .Y(n_1039) );
OR2x6_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g816 ( .A(n_654), .Y(n_816) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx4_ASAP7_75t_SL g683 ( .A(n_663), .Y(n_683) );
XOR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_682), .Y(n_663) );
NAND3x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_674), .C(n_679), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .C(n_673), .Y(n_669) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g1124 ( .A(n_684), .Y(n_1124) );
XNOR2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_978), .Y(n_684) );
AOI22xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_906), .B1(n_976), .B2(n_977), .Y(n_685) );
INVx1_ASAP7_75t_L g976 ( .A(n_686), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_747), .B1(n_904), .B2(n_905), .Y(n_686) );
INVx1_ASAP7_75t_L g904 ( .A(n_687), .Y(n_904) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_723), .B1(n_724), .B2(n_746), .Y(n_689) );
INVx1_ASAP7_75t_L g746 ( .A(n_690), .Y(n_746) );
INVx1_ASAP7_75t_L g722 ( .A(n_692), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .C(n_705), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_707), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_711), .B(n_718), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_SL g814 ( .A(n_714), .Y(n_814) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
XOR2x2_ASAP7_75t_L g782 ( .A(n_724), .B(n_783), .Y(n_782) );
XOR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_745), .Y(n_724) );
NAND4xp75_ASAP7_75t_SL g725 ( .A(n_726), .B(n_728), .C(n_730), .D(n_736), .Y(n_725) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_734), .Y(n_730) );
BUFx2_ASAP7_75t_L g990 ( .A(n_735), .Y(n_990) );
INVx1_ASAP7_75t_L g1020 ( .A(n_735), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B(n_740), .Y(n_737) );
OAI222xp33_ASAP7_75t_L g1074 ( .A1(n_739), .A2(n_1075), .B1(n_1076), .B2(n_1077), .C1(n_1078), .C2(n_1079), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_744), .Y(n_797) );
INVx1_ASAP7_75t_L g905 ( .A(n_747), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_809), .B2(n_903), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_782), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
XOR2x2_ASAP7_75t_L g878 ( .A(n_751), .B(n_879), .Y(n_878) );
XNOR2x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_781), .Y(n_751) );
AND3x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_763), .C(n_770), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .C(n_760), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_776), .C(n_779), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_774), .B2(n_775), .Y(n_771) );
BUFx2_ASAP7_75t_R g993 ( .A(n_775), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g823 ( .A(n_778), .Y(n_823) );
XNOR2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_800), .C(n_804), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_793), .Y(n_786) );
OAI21xp5_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_789), .B(n_790), .Y(n_787) );
OAI21xp5_ASAP7_75t_SL g1008 ( .A1(n_788), .A2(n_1009), .B(n_1010), .Y(n_1008) );
BUFx4f_ASAP7_75t_L g839 ( .A(n_792), .Y(n_839) );
INVx1_ASAP7_75t_L g1078 ( .A(n_792), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .Y(n_800) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g1094 ( .A(n_806), .Y(n_1094) );
INVx2_ASAP7_75t_L g903 ( .A(n_809), .Y(n_903) );
XNOR2x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_847), .Y(n_809) );
INVx1_ASAP7_75t_L g846 ( .A(n_811), .Y(n_846) );
AND2x2_ASAP7_75t_SL g811 ( .A(n_812), .B(n_828), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_820), .Y(n_812) );
OAI221xp5_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .C(n_818), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_814), .A2(n_822), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
INVx4_ASAP7_75t_L g1063 ( .A(n_819), .Y(n_1063) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .C(n_840), .Y(n_828) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx3_ASAP7_75t_SL g893 ( .A(n_843), .Y(n_893) );
AO22x2_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_878), .B2(n_902), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_866), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .C(n_861), .Y(n_853) );
OAI21xp5_ASAP7_75t_SL g895 ( .A1(n_856), .A2(n_896), .B(n_897), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_863), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
BUFx6f_ASAP7_75t_L g919 ( .A(n_864), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_867), .B(n_872), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_871), .Y(n_988) );
INVx2_ASAP7_75t_L g1028 ( .A(n_871), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_877), .Y(n_872) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g902 ( .A(n_878), .Y(n_902) );
XNOR2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
NAND3x1_ASAP7_75t_SL g881 ( .A(n_882), .B(n_885), .C(n_888), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_895), .C(n_898), .Y(n_888) );
OAI22xp5_ASAP7_75t_SL g889 ( .A1(n_890), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g977 ( .A(n_906), .Y(n_977) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OA22x2_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_936), .B1(n_974), .B2(n_975), .Y(n_907) );
INVx1_ASAP7_75t_L g974 ( .A(n_908), .Y(n_974) );
INVx2_ASAP7_75t_SL g934 ( .A(n_909), .Y(n_934) );
AND2x2_ASAP7_75t_SL g909 ( .A(n_910), .B(n_924), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_914), .C(n_920), .Y(n_910) );
OAI21xp33_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B(n_918), .Y(n_914) );
OAI21xp33_ASAP7_75t_L g1036 ( .A1(n_916), .A2(n_1037), .B(n_1038), .Y(n_1036) );
INVx3_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_919), .Y(n_1076) );
AND4x1_ASAP7_75t_L g924 ( .A(n_925), .B(n_927), .C(n_929), .D(n_931), .Y(n_924) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
OAI221xp5_ASAP7_75t_SL g1147 ( .A1(n_933), .A2(n_1148), .B1(n_1149), .B2(n_1150), .C(n_1151), .Y(n_1147) );
INVx1_ASAP7_75t_L g975 ( .A(n_936), .Y(n_975) );
XOR2x2_ASAP7_75t_L g936 ( .A(n_937), .B(n_955), .Y(n_936) );
XOR2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_954), .Y(n_937) );
NAND4xp75_ASAP7_75t_SL g938 ( .A(n_939), .B(n_948), .C(n_951), .D(n_952), .Y(n_938) );
NOR2xp67_ASAP7_75t_SL g939 ( .A(n_940), .B(n_944), .Y(n_939) );
NAND3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .C(n_943), .Y(n_940) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
XOR2x2_ASAP7_75t_SL g955 ( .A(n_956), .B(n_973), .Y(n_955) );
NAND2x1p5_ASAP7_75t_L g956 ( .A(n_957), .B(n_966), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_963), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_961), .C(n_962), .Y(n_958) );
NOR2x1_ASAP7_75t_L g966 ( .A(n_967), .B(n_970), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_1050), .B1(n_1122), .B2(n_1123), .Y(n_978) );
INVx1_ASAP7_75t_L g1123 ( .A(n_979), .Y(n_1123) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1002), .B1(n_1003), .B2(n_1049), .Y(n_980) );
INVx1_ASAP7_75t_L g1049 ( .A(n_981), .Y(n_1049) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
AND4x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_989), .C(n_996), .D(n_1000), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_991) );
OAI22xp5_ASAP7_75t_SL g1088 ( .A1(n_993), .A2(n_1089), .B1(n_1090), .B2(n_1091), .Y(n_1088) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AO22x1_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1029), .B2(n_1030), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
NAND4xp75_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1017), .C(n_1023), .D(n_1026), .Y(n_1006) );
NOR2xp67_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1011), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .C(n_1016), .Y(n_1011) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1021), .Y(n_1017) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_SL g1047 ( .A(n_1031), .Y(n_1047) );
AND2x2_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1042), .Y(n_1031) );
NOR3xp33_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1036), .C(n_1039), .Y(n_1032) );
AND4x1_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1044), .C(n_1045), .D(n_1046), .Y(n_1042) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1050), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1070), .B1(n_1120), .B2(n_1121), .Y(n_1051) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1052), .Y(n_1121) );
INVx1_ASAP7_75t_SL g1069 ( .A(n_1054), .Y(n_1069) );
NAND4xp75_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1059), .C(n_1064), .D(n_1068), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1058), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
INVx3_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
AND2x2_ASAP7_75t_SL g1064 ( .A(n_1065), .B(n_1067), .Y(n_1064) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1070), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1095), .B1(n_1118), .B2(n_1119), .Y(n_1070) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1071), .Y(n_1119) );
NAND3x1_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1083), .C(n_1087), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1080), .Y(n_1073) );
OAI221xp5_ASAP7_75t_SL g1183 ( .A1(n_1076), .A2(n_1184), .B1(n_1185), .B2(n_1186), .C(n_1187), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1086), .Y(n_1149) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1095), .Y(n_1118) );
XNOR2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1107), .Y(n_1097) );
NOR3xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1111), .C(n_1115), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_SL g1125 ( .A(n_1126), .Y(n_1125) );
NOR2x1_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1131), .Y(n_1126) );
OR2x2_ASAP7_75t_SL g1201 ( .A(n_1127), .B(n_1132), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1130), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1129), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1129), .B(n_1168), .Y(n_1172) );
CKINVDCx16_ASAP7_75t_R g1168 ( .A(n_1130), .Y(n_1168) );
CKINVDCx20_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1134), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
OAI322xp33_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1165), .A3(n_1166), .B1(n_1169), .B2(n_1173), .C1(n_1174), .C2(n_1199), .Y(n_1138) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1140), .Y(n_1164) );
AND2x2_ASAP7_75t_SL g1140 ( .A(n_1141), .B(n_1152), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1147), .Y(n_1141) );
NOR3xp33_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1156), .C(n_1160), .Y(n_1152) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
CKINVDCx20_ASAP7_75t_R g1169 ( .A(n_1170), .Y(n_1169) );
CKINVDCx20_ASAP7_75t_R g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_1178), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1191), .Y(n_1178) );
NOR3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1183), .C(n_1188), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1196), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1198), .Y(n_1196) );
CKINVDCx20_ASAP7_75t_R g1199 ( .A(n_1200), .Y(n_1199) );
CKINVDCx20_ASAP7_75t_R g1200 ( .A(n_1201), .Y(n_1200) );
endmodule