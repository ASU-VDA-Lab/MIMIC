module fake_aes_4655_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_SL g3 ( .A(n_1), .Y(n_3) );
BUFx4f_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
AO31x2_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .A3(n_1), .B(n_2), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x4_ASAP7_75t_L g8 ( .A(n_7), .B(n_5), .Y(n_8) );
AOI222xp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_4), .B1(n_6), .B2(n_5), .C1(n_0), .C2(n_2), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
NAND3xp33_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .C(n_5), .Y(n_11) );
OAI21xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_6), .B(n_4), .Y(n_12) );
endmodule