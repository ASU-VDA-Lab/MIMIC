module real_jpeg_30734_n_13 (n_123, n_8, n_116, n_0, n_2, n_114, n_10, n_9, n_12, n_124, n_6, n_121, n_11, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_120, n_13);

input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_124;
input n_6;
input n_121;
input n_11;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_120;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_1),
.B(n_48),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_5),
.A2(n_34),
.A3(n_36),
.B1(n_46),
.B2(n_108),
.C1(n_110),
.C2(n_124),
.Y(n_107)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_11),
.B1(n_71),
.B2(n_75),
.C(n_79),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_71),
.C(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_9),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_22),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI31xp67_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_59),
.A3(n_97),
.B(n_103),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_45),
.C(n_53),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_26),
.A2(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_28),
.B(n_53),
.C(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_115),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OA21x2_ASAP7_75t_SL g104 ( 
.A1(n_45),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_92),
.C(n_93),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_83),
.B(n_91),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_70),
.B1(n_81),
.B2(n_82),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_120),
.Y(n_75)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_114),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_116),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_117),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_118),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_119),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_121),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_122),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_123),
.Y(n_100)
);


endmodule