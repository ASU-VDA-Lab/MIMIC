module fake_jpeg_2276_n_640 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_640);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_640;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_10),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g199 ( 
.A(n_62),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_64),
.Y(n_152)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_60),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_75),
.Y(n_202)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_32),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_89),
.Y(n_181)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_19),
.B(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_95),
.B(n_38),
.Y(n_173)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_31),
.B(n_6),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g165 ( 
.A(n_122),
.Y(n_165)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

AND2x4_ASAP7_75t_SL g124 ( 
.A(n_30),
.B(n_18),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_54),
.Y(n_167)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_55),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_128),
.B(n_16),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_138),
.B(n_153),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_55),
.B1(n_59),
.B2(n_38),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_140),
.A2(n_169),
.B1(n_170),
.B2(n_177),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_173),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_80),
.A2(n_32),
.B1(n_56),
.B2(n_55),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_161),
.A2(n_172),
.B1(n_191),
.B2(n_177),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_30),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_163),
.B(n_164),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_68),
.A2(n_56),
.B1(n_70),
.B2(n_127),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_69),
.A2(n_114),
.B1(n_124),
.B2(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_89),
.A2(n_32),
.B1(n_60),
.B2(n_22),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_63),
.B(n_45),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_174),
.B(n_180),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_73),
.A2(n_56),
.B1(n_55),
.B2(n_49),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_59),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_75),
.A2(n_47),
.B1(n_43),
.B2(n_58),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_184),
.A2(n_186),
.B1(n_57),
.B2(n_5),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_77),
.A2(n_47),
.B1(n_43),
.B2(n_58),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_82),
.B(n_45),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_197),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_80),
.A2(n_41),
.B1(n_54),
.B2(n_36),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_101),
.B(n_48),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_14),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_92),
.A2(n_94),
.B1(n_100),
.B2(n_41),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_54),
.B1(n_57),
.B2(n_37),
.Y(n_261)
);

INVx6_ASAP7_75t_SL g212 ( 
.A(n_122),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g224 ( 
.A(n_212),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_213),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_214),
.B(n_231),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_48),
.B1(n_44),
.B2(n_36),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_217),
.A2(n_261),
.B1(n_264),
.B2(n_278),
.Y(n_337)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_222),
.Y(n_288)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_225),
.Y(n_310)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_227),
.Y(n_317)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_228),
.Y(n_339)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_199),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_143),
.B(n_39),
.C(n_49),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_230),
.B(n_263),
.C(n_1),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_148),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_181),
.A2(n_44),
.B1(n_39),
.B2(n_41),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_232),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_290)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_145),
.Y(n_236)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_132),
.B(n_149),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_241),
.Y(n_298)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_155),
.Y(n_240)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_103),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_243),
.B(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_245),
.Y(n_327)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_246),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_129),
.Y(n_247)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_168),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_163),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_284),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_142),
.A2(n_99),
.B1(n_110),
.B2(n_105),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_254),
.A2(n_206),
.B1(n_146),
.B2(n_200),
.Y(n_332)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_168),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_260),
.Y(n_320)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_134),
.Y(n_257)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_154),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_259),
.Y(n_294)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_41),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_267),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_167),
.B(n_112),
.C(n_106),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_166),
.B1(n_204),
.B2(n_202),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_146),
.Y(n_266)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_131),
.A2(n_54),
.B1(n_106),
.B2(n_112),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_12),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_271),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_195),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_272),
.Y(n_335)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_275),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_274),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_210),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_130),
.B(n_0),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_277),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_201),
.A2(n_57),
.B1(n_5),
.B2(n_13),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_162),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_279),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_5),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_156),
.B1(n_159),
.B2(n_189),
.Y(n_291)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_162),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_141),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_152),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_285),
.B1(n_146),
.B2(n_144),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_179),
.B(n_0),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_199),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_287),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_179),
.B(n_1),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

AOI22x1_ASAP7_75t_L g301 ( 
.A1(n_221),
.A2(n_161),
.B1(n_191),
.B2(n_147),
.Y(n_301)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_301),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_216),
.A2(n_209),
.B1(n_200),
.B2(n_204),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_329),
.B1(n_346),
.B2(n_285),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_251),
.A2(n_137),
.B1(n_150),
.B2(n_157),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g394 ( 
.A1(n_314),
.A2(n_332),
.B1(n_286),
.B2(n_266),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_221),
.B(n_171),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_315),
.B(n_254),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_252),
.A2(n_171),
.B1(n_144),
.B2(n_192),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_322),
.Y(n_358)
);

AO22x1_ASAP7_75t_SL g322 ( 
.A1(n_221),
.A2(n_192),
.B1(n_157),
.B2(n_206),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_261),
.A2(n_277),
.B1(n_234),
.B2(n_284),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_209),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_336),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_215),
.B(n_57),
.C(n_13),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_213),
.C(n_251),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_1),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_250),
.B(n_1),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_338),
.B(n_347),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_219),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_251),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_267),
.B1(n_229),
.B2(n_227),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_263),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_265),
.A2(n_15),
.B(n_18),
.C(n_4),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_298),
.B(n_239),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_352),
.A2(n_365),
.B1(n_372),
.B2(n_375),
.Y(n_417)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_294),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_359),
.Y(n_411)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_230),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_360),
.B(n_361),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_344),
.A2(n_246),
.B1(n_273),
.B2(n_228),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_362),
.A2(n_366),
.B(n_316),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_257),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_363),
.B(n_377),
.C(n_386),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_224),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_367),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_315),
.B(n_244),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_294),
.Y(n_368)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_294),
.Y(n_369)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_224),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_370),
.B(n_376),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_262),
.B1(n_281),
.B2(n_279),
.Y(n_372)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_308),
.A2(n_272),
.B1(n_249),
.B2(n_255),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_312),
.B(n_224),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_292),
.B(n_259),
.C(n_226),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_245),
.B1(n_218),
.B2(n_220),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_379),
.A2(n_381),
.B1(n_389),
.B2(n_332),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_337),
.A2(n_258),
.B1(n_244),
.B2(n_233),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_335),
.Y(n_382)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_382),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_289),
.Y(n_384)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_299),
.A2(n_306),
.B1(n_335),
.B2(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_385),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_320),
.B(n_222),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_387),
.B(n_392),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_223),
.B1(n_274),
.B2(n_235),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_237),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_390),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_391),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_292),
.B(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_289),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_393),
.B(n_395),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_394),
.A2(n_317),
.B1(n_306),
.B2(n_339),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_338),
.B(n_268),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_308),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_401),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_336),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_301),
.B(n_299),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_402),
.A2(n_403),
.B(n_412),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_301),
.B(n_299),
.Y(n_403)
);

AO22x1_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_322),
.B1(n_324),
.B2(n_346),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_425),
.Y(n_472)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_388),
.A2(n_345),
.B1(n_331),
.B2(n_290),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_358),
.B1(n_390),
.B2(n_365),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_305),
.B(n_347),
.Y(n_412)
);

OA22x2_ASAP7_75t_L g470 ( 
.A1(n_424),
.A2(n_328),
.B1(n_317),
.B2(n_321),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_309),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_380),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_351),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_358),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_435),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_431),
.A2(n_432),
.B(n_402),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_366),
.A2(n_349),
.B(n_358),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_352),
.A2(n_330),
.B1(n_303),
.B2(n_304),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_433),
.A2(n_417),
.B1(n_409),
.B2(n_407),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_386),
.B(n_363),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_436),
.A2(n_438),
.B1(n_444),
.B2(n_445),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_439),
.B1(n_453),
.B2(n_456),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_360),
.B1(n_349),
.B2(n_389),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_417),
.A2(n_362),
.B1(n_395),
.B2(n_356),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_397),
.Y(n_440)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_374),
.B1(n_375),
.B2(n_378),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_406),
.A2(n_361),
.B1(n_392),
.B2(n_372),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_368),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_455),
.C(n_458),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_447),
.B(n_463),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_406),
.A2(n_382),
.B1(n_391),
.B2(n_369),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_449),
.A2(n_451),
.B(n_459),
.Y(n_491)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_452),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_379),
.B1(n_353),
.B2(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_303),
.C(n_304),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_393),
.B1(n_384),
.B2(n_291),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_414),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_457),
.B(n_416),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_418),
.C(n_423),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_432),
.A2(n_355),
.B(n_325),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_325),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_461),
.C(n_414),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_425),
.C(n_411),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_310),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_400),
.C(n_457),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_426),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_426),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_471),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_403),
.A2(n_330),
.B1(n_373),
.B2(n_319),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_408),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_398),
.A2(n_319),
.B1(n_367),
.B2(n_310),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_434),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_422),
.A2(n_351),
.B1(n_383),
.B2(n_380),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_424),
.Y(n_478)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

AO22x1_ASAP7_75t_L g474 ( 
.A1(n_439),
.A2(n_427),
.B1(n_409),
.B2(n_407),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_453),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_483),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_472),
.Y(n_477)
);

BUFx4f_ASAP7_75t_SL g507 ( 
.A(n_478),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_411),
.B1(n_433),
.B2(n_427),
.Y(n_479)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_482),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_442),
.A2(n_427),
.B1(n_416),
.B2(n_413),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_498),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_461),
.Y(n_487)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_466),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_488),
.B(n_494),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_401),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_451),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_437),
.A2(n_413),
.B1(n_412),
.B2(n_420),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_490),
.A2(n_496),
.B1(n_469),
.B2(n_470),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_445),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_463),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_420),
.B1(n_400),
.B2(n_428),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_399),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_497),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_455),
.B(n_415),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_431),
.B(n_396),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_491),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_458),
.B(n_328),
.C(n_340),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_503),
.C(n_459),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_340),
.C(n_321),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_441),
.B(n_415),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_504),
.B(n_441),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_515),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_511),
.B(n_512),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_489),
.B(n_448),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_438),
.C(n_449),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_522),
.C(n_524),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_464),
.B1(n_436),
.B2(n_467),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_517),
.A2(n_519),
.B1(n_525),
.B2(n_534),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_518),
.B(n_523),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_495),
.A2(n_444),
.B1(n_448),
.B2(n_456),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_508),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_481),
.B(n_440),
.Y(n_521)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_521),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_502),
.C(n_492),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_505),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_471),
.C(n_452),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_475),
.A2(n_468),
.B1(n_454),
.B2(n_450),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_443),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_483),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_505),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_528),
.B(n_499),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_529),
.A2(n_531),
.B1(n_478),
.B2(n_474),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_470),
.C(n_396),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_533),
.C(n_485),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_491),
.A2(n_470),
.B(n_421),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_497),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_501),
.B(n_309),
.C(n_295),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_475),
.A2(n_421),
.B1(n_419),
.B2(n_383),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_496),
.A2(n_419),
.B1(n_343),
.B2(n_295),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_535),
.A2(n_481),
.B1(n_478),
.B2(n_493),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_536),
.A2(n_518),
.B1(n_519),
.B2(n_509),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_541),
.B(n_550),
.Y(n_566)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_542),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_490),
.C(n_479),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_543),
.B(n_530),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_544),
.B(n_545),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_520),
.B(n_474),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_527),
.Y(n_546)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_546),
.Y(n_580)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_547),
.Y(n_565)
);

FAx1_ASAP7_75t_SL g548 ( 
.A(n_512),
.B(n_511),
.CI(n_516),
.CON(n_548),
.SN(n_548)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_548),
.B(n_524),
.Y(n_562)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_500),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_552),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_526),
.B(n_497),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_553),
.A2(n_555),
.B1(n_560),
.B2(n_525),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_513),
.B(n_485),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_557),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_514),
.B(n_484),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_517),
.B(n_476),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_558),
.Y(n_564)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_559),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_237),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_575),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_510),
.C(n_532),
.Y(n_567)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_569),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_556),
.A2(n_531),
.B1(n_507),
.B2(n_534),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_570),
.A2(n_571),
.B1(n_581),
.B2(n_561),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_539),
.A2(n_536),
.B1(n_555),
.B2(n_558),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_538),
.B(n_480),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_540),
.B(n_535),
.C(n_480),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_SL g588 ( 
.A(n_576),
.B(n_579),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_540),
.B(n_507),
.C(n_293),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_539),
.A2(n_507),
.B1(n_343),
.B2(n_293),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_544),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_583),
.B(n_594),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_543),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_586),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_585),
.A2(n_597),
.B1(n_571),
.B2(n_581),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_566),
.B(n_541),
.C(n_551),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_578),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_587),
.B(n_591),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_566),
.B(n_550),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_580),
.Y(n_592)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_552),
.B1(n_548),
.B2(n_545),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_593),
.B(n_596),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_537),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_568),
.A2(n_537),
.B1(n_326),
.B2(n_307),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_595),
.B(n_574),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_327),
.C(n_313),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_576),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_599),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_579),
.B(n_313),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_582),
.A2(n_570),
.B(n_564),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_605),
.A2(n_610),
.B1(n_326),
.B2(n_282),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_589),
.B(n_573),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_606),
.B(n_609),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_607),
.B(n_599),
.Y(n_616)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_608),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_590),
.B(n_565),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_597),
.A2(n_564),
.B(n_577),
.Y(n_610)
);

AOI21xp33_ASAP7_75t_L g611 ( 
.A1(n_595),
.A2(n_565),
.B(n_574),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_611),
.A2(n_596),
.B(n_594),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_586),
.A2(n_588),
.B(n_583),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_613),
.A2(n_300),
.B(n_307),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_600),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_614),
.A2(n_615),
.B1(n_620),
.B2(n_621),
.Y(n_624)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_616),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_592),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_617),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_327),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_623),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_247),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_623),
.A2(n_612),
.B(n_300),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_SL g627 ( 
.A1(n_619),
.A2(n_605),
.B(n_610),
.C(n_607),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_627),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_618),
.B(n_602),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_628),
.A2(n_630),
.B(n_617),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_629),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_633),
.B(n_634),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_625),
.A2(n_608),
.B1(n_612),
.B2(n_18),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_632),
.A2(n_626),
.B(n_624),
.Y(n_636)
);

AOI31xp33_ASAP7_75t_L g637 ( 
.A1(n_636),
.A2(n_631),
.A3(n_627),
.B(n_18),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_637),
.A2(n_635),
.B(n_3),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_2),
.C(n_4),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g640 ( 
.A(n_639),
.Y(n_640)
);


endmodule