module fake_netlist_6_2108_n_971 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_33, n_27, n_3, n_14, n_0, n_32, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_971);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_0;
input n_32;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_971;

wire n_52;
wire n_591;
wire n_435;
wire n_91;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_63;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_828;
wire n_161;
wire n_208;
wire n_462;
wire n_68;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_50;
wire n_694;
wire n_933;
wire n_740;
wire n_703;
wire n_578;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_77;
wire n_820;
wire n_951;
wire n_783;
wire n_106;
wire n_725;
wire n_952;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_131;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_78;
wire n_84;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_142;
wire n_874;
wire n_724;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_62;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_67;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_38;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_59;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_108;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_65;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_71;
wire n_74;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_72;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_111;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_35;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_79;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_56;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_119;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_39;
wire n_344;
wire n_73;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_101;
wire n_167;
wire n_631;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_842;
wire n_758;
wire n_943;
wire n_611;
wire n_156;
wire n_491;
wire n_878;
wire n_145;
wire n_42;
wire n_133;
wire n_656;
wire n_772;
wire n_96;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_129;
wire n_705;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_122;
wire n_930;
wire n_888;
wire n_45;
wire n_454;
wire n_218;
wire n_638;
wire n_70;
wire n_234;
wire n_910;
wire n_37;
wire n_486;
wire n_911;
wire n_381;
wire n_82;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_112;
wire n_172;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_58;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_118;
wire n_224;
wire n_48;
wire n_926;
wire n_927;
wire n_93;
wire n_839;
wire n_80;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_107;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_89;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_103;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_69;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_53;
wire n_370;
wire n_44;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_46;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_83;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_813;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_92;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_105;
wire n_916;
wire n_227;
wire n_132;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_102;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_811;
wire n_312;
wire n_394;
wire n_66;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_630;
wire n_958;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_61;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_548;
wire n_905;
wire n_94;
wire n_282;
wire n_436;
wire n_833;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_40;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_139;
wire n_319;
wire n_41;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_95;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_123;
wire n_136;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_43;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_49;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_90;
wire n_347;
wire n_812;
wire n_459;
wire n_54;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_85;
wire n_99;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_47;
wire n_690;
wire n_850;
wire n_75;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_110;
wire n_151;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_81;
wire n_660;
wire n_965;
wire n_36;
wire n_55;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_64;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_135;
wire n_165;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_60;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_57;
wire n_169;
wire n_51;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

INVxp33_ASAP7_75t_SL g80 ( 
.A(n_41),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_55),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_40),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_40),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_56),
.B1(n_59),
.B2(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_66),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_56),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_43),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

OR2x6_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_47),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_39),
.B1(n_52),
.B2(n_55),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NOR2x1p5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_53),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_67),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_43),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_47),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_62),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_61),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_59),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

OR2x6_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_34),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_100),
.Y(n_159)
);

AO22x2_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_102),
.B1(n_101),
.B2(n_94),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

OR2x6_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_106),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_89),
.B1(n_88),
.B2(n_109),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_102),
.B1(n_101),
.B2(n_99),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_102),
.B1(n_89),
.B2(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_109),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

OAI221xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_109),
.B1(n_92),
.B2(n_58),
.C(n_44),
.Y(n_179)
);

OAI221xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_92),
.B1(n_45),
.B2(n_60),
.C(n_46),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_108),
.B1(n_97),
.B2(n_92),
.Y(n_181)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_107),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_123),
.B1(n_142),
.B2(n_147),
.Y(n_183)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_52),
.B1(n_107),
.B2(n_106),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_108),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_138),
.B(n_97),
.Y(n_186)
);

AO22x2_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_107),
.B1(n_106),
.B2(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_50),
.B1(n_49),
.B2(n_107),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_27),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_129),
.Y(n_190)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_149),
.B1(n_145),
.B2(n_126),
.Y(n_191)
);

NAND2x1p5_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

NAND2x1p5_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_107),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_107),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_106),
.Y(n_201)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_106),
.B1(n_2),
.B2(n_4),
.Y(n_202)
);

AO22x2_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_106),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_128),
.B(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

AO22x2_ASAP7_75t_L g210 ( 
.A1(n_126),
.A2(n_106),
.B1(n_6),
.B2(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_157),
.B(n_0),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g214 ( 
.A1(n_145),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_214)
);

NAND2x1p5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_24),
.Y(n_215)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_13),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_122),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

OAI221xp5_ASAP7_75t_L g228 ( 
.A1(n_156),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.C(n_122),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_164),
.B(n_157),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_164),
.B(n_157),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_196),
.B(n_157),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_199),
.B(n_157),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_185),
.B(n_127),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_161),
.B(n_127),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_169),
.B(n_127),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_169),
.B(n_127),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_150),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_155),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_150),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_139),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_188),
.B(n_150),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_188),
.B(n_150),
.Y(n_245)
);

NAND2x1p5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_219),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_182),
.B(n_148),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_182),
.B(n_125),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_192),
.B(n_125),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_139),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_192),
.B(n_119),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_144),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_195),
.B(n_130),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_139),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_195),
.B(n_130),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_SL g256 ( 
.A(n_218),
.B(n_144),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_155),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_155),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g259 ( 
.A(n_211),
.B(n_220),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_220),
.B(n_144),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_190),
.B(n_130),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_176),
.B(n_141),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_186),
.B(n_141),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_141),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_163),
.B(n_137),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_163),
.B(n_137),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_SL g267 ( 
.A(n_189),
.B(n_137),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_181),
.B(n_120),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_181),
.B(n_120),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_209),
.B(n_120),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_189),
.B(n_155),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_209),
.B(n_112),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_221),
.B(n_112),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_132),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_222),
.B(n_113),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_183),
.B(n_132),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_224),
.B(n_136),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_225),
.B(n_136),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_226),
.B(n_206),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_206),
.B(n_155),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_193),
.B(n_132),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_216),
.B(n_136),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_194),
.B(n_132),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_174),
.B(n_115),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_216),
.B(n_136),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_183),
.B(n_204),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_158),
.B(n_121),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_215),
.B(n_136),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_162),
.B(n_115),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_215),
.B(n_115),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_115),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_175),
.B(n_115),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_177),
.B(n_178),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_212),
.B(n_173),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_212),
.B(n_171),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_165),
.B(n_208),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_160),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_264),
.A2(n_167),
.B(n_159),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_160),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_243),
.A2(n_191),
.B(n_168),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_248),
.A2(n_168),
.B(n_191),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_249),
.A2(n_168),
.B(n_179),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_170),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_180),
.C(n_179),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_251),
.B(n_244),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_170),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

OAI21x1_ASAP7_75t_SL g310 ( 
.A1(n_276),
.A2(n_203),
.B(n_202),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_187),
.B(n_203),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_245),
.A2(n_187),
.B(n_202),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_238),
.A2(n_239),
.B(n_247),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_234),
.A2(n_228),
.B(n_174),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_228),
.B(n_210),
.C(n_184),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_184),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_253),
.A2(n_210),
.B(n_214),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_250),
.A2(n_223),
.B(n_214),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_258),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_223),
.B(n_254),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_R g324 ( 
.A(n_233),
.B(n_252),
.Y(n_324)
);

AO31x2_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_292),
.A3(n_291),
.B(n_287),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_255),
.A2(n_236),
.B(n_263),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_241),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_258),
.B(n_270),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_246),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_268),
.B(n_269),
.Y(n_332)
);

NOR2x1_ASAP7_75t_SL g333 ( 
.A(n_282),
.B(n_285),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_240),
.A2(n_242),
.B1(n_278),
.B2(n_277),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_275),
.B(n_273),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_262),
.A2(n_259),
.B(n_296),
.Y(n_336)
);

O2A1O1Ixp5_ASAP7_75t_L g337 ( 
.A1(n_260),
.A2(n_267),
.B(n_271),
.C(n_280),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_281),
.A2(n_283),
.B(n_272),
.Y(n_339)
);

NAND3x1_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_295),
.C(n_265),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_164),
.Y(n_341)
);

OAI21x1_ASAP7_75t_L g342 ( 
.A1(n_264),
.A2(n_206),
.B(n_243),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_248),
.A2(n_127),
.B(n_229),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_276),
.A2(n_286),
.B(n_239),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_230),
.B(n_164),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_241),
.B(n_257),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_238),
.A2(n_164),
.B(n_239),
.Y(n_348)
);

BUFx8_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

AO31x2_ASAP7_75t_L g350 ( 
.A1(n_276),
.A2(n_286),
.A3(n_220),
.B(n_137),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_241),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_230),
.B(n_164),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_238),
.A2(n_164),
.B(n_239),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_238),
.A2(n_164),
.B1(n_131),
.B2(n_239),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_238),
.A2(n_229),
.B(n_131),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_241),
.B(n_257),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_241),
.B(n_257),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_246),
.Y(n_358)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_241),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_276),
.A2(n_286),
.B(n_239),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_230),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_264),
.A2(n_206),
.B(n_243),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_248),
.A2(n_127),
.B(n_229),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_276),
.A2(n_286),
.B(n_239),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_230),
.B(n_164),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_248),
.A2(n_127),
.B(n_229),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_300),
.B1(n_328),
.B2(n_313),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_348),
.A2(n_353),
.B(n_312),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

AO21x2_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_302),
.B(n_303),
.Y(n_371)
);

OR2x6_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_339),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_365),
.B1(n_352),
.B2(n_361),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_297),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_305),
.A2(n_341),
.B(n_307),
.C(n_337),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_298),
.A2(n_342),
.B(n_362),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_301),
.A2(n_326),
.B(n_366),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

AO31x2_ASAP7_75t_L g380 ( 
.A1(n_316),
.A2(n_354),
.A3(n_299),
.B(n_333),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_329),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_357),
.B1(n_356),
.B2(n_347),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_336),
.B(n_319),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_319),
.A2(n_315),
.B(n_321),
.Y(n_387)
);

OAI21x1_ASAP7_75t_SL g388 ( 
.A1(n_310),
.A2(n_304),
.B(n_308),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_309),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_356),
.A2(n_357),
.B(n_316),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_351),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_320),
.A2(n_309),
.B1(n_359),
.B2(n_331),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_338),
.A2(n_330),
.B(n_327),
.C(n_334),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_331),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_309),
.A2(n_330),
.B1(n_327),
.B2(n_358),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_325),
.B(n_364),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_343),
.A2(n_363),
.B(n_335),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_358),
.A2(n_331),
.B1(n_360),
.B2(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

OAI21x1_ASAP7_75t_SL g401 ( 
.A1(n_344),
.A2(n_364),
.B(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_340),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_311),
.A2(n_350),
.B(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

OR2x6_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_355),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_306),
.A2(n_317),
.B1(n_323),
.B2(n_311),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_340),
.A2(n_323),
.B1(n_317),
.B2(n_324),
.Y(n_410)
);

AO21x2_ASAP7_75t_L g411 ( 
.A1(n_324),
.A2(n_350),
.B(n_323),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_361),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_164),
.Y(n_415)
);

AO21x2_ASAP7_75t_L g416 ( 
.A1(n_314),
.A2(n_302),
.B(n_348),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_322),
.A2(n_164),
.B1(n_300),
.B2(n_328),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

OAI211xp5_ASAP7_75t_L g420 ( 
.A1(n_345),
.A2(n_89),
.B(n_88),
.C(n_169),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_106),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_297),
.B(n_308),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_341),
.A2(n_164),
.B(n_352),
.C(n_345),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_298),
.A2(n_314),
.B(n_342),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_318),
.B(n_346),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_341),
.B(n_164),
.C(n_148),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_SL g430 ( 
.A(n_341),
.B(n_152),
.C(n_129),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_298),
.A2(n_314),
.B(n_342),
.Y(n_431)
);

OAI21x1_ASAP7_75t_SL g432 ( 
.A1(n_387),
.A2(n_388),
.B(n_368),
.Y(n_432)
);

AO21x2_ASAP7_75t_L g433 ( 
.A1(n_401),
.A2(n_376),
.B(n_405),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

CKINVDCx6p67_ASAP7_75t_R g435 ( 
.A(n_408),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_370),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_406),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_377),
.A2(n_378),
.B(n_427),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_429),
.B1(n_402),
.B2(n_424),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_428),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_380),
.Y(n_442)
);

NAND4xp25_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_430),
.C(n_420),
.D(n_414),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_422),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_408),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_406),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_411),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_377),
.A2(n_431),
.B(n_427),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_372),
.B(n_406),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_416),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx4_ASAP7_75t_SL g470 ( 
.A(n_406),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_428),
.B(n_380),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_380),
.B(n_424),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_458),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_413),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_R g476 ( 
.A(n_436),
.B(n_412),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_436),
.Y(n_479)
);

OR2x4_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_394),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_373),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g482 ( 
.A(n_449),
.B(n_412),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_413),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_444),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_369),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_R g488 ( 
.A(n_450),
.B(n_369),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_419),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_439),
.B(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_385),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_419),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_385),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_382),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_382),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_446),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_R g499 ( 
.A(n_450),
.B(n_369),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_462),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_439),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_443),
.B(n_391),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_384),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_450),
.B(n_381),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_SL g508 ( 
.A(n_437),
.B(n_392),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_418),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_450),
.B(n_390),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_R g511 ( 
.A(n_450),
.B(n_423),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_418),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_456),
.B(n_426),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_456),
.B(n_383),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_372),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_R g516 ( 
.A(n_460),
.B(n_372),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_389),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_R g522 ( 
.A(n_460),
.B(n_397),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_437),
.B(n_398),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_456),
.B(n_367),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_460),
.B(n_397),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_470),
.B(n_407),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_390),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_457),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_496),
.B(n_457),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_501),
.A2(n_432),
.B1(n_460),
.B2(n_434),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_496),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_494),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_515),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_454),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_457),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_515),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_512),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_512),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_476),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_491),
.Y(n_545)
);

BUFx2_ASAP7_75t_SL g546 ( 
.A(n_517),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_493),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_493),
.B(n_467),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g551 ( 
.A(n_490),
.B(n_468),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_479),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_481),
.B(n_454),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_510),
.B(n_460),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_514),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_454),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_455),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_513),
.B(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_521),
.B(n_464),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_527),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_528),
.B(n_464),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_464),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_464),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_526),
.B(n_463),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_474),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_511),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_483),
.B(n_461),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_L g575 ( 
.A(n_506),
.B(n_445),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_504),
.A2(n_434),
.B1(n_442),
.B2(n_421),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_475),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_500),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_484),
.B(n_447),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_530),
.B(n_442),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_530),
.B(n_568),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_563),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_530),
.B(n_433),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_538),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_548),
.B(n_467),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_433),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_555),
.B(n_470),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_538),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_541),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_532),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_548),
.B(n_467),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_568),
.B(n_433),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_532),
.Y(n_598)
);

NOR2x1_ASAP7_75t_L g599 ( 
.A(n_551),
.B(n_502),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_532),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_563),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_572),
.A2(n_508),
.B1(n_503),
.B2(n_482),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_529),
.B(n_433),
.Y(n_606)
);

NAND2x1_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_517),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_552),
.B(n_505),
.Y(n_608)
);

OA21x2_ASAP7_75t_L g609 ( 
.A1(n_577),
.A2(n_438),
.B(n_459),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_580),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_548),
.B(n_468),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_544),
.A2(n_477),
.B1(n_410),
.B2(n_437),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_535),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_535),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_546),
.B(n_453),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_545),
.B(n_469),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_572),
.B(n_473),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_468),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_529),
.B(n_433),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_549),
.B(n_469),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_571),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_577),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

INVx3_ASAP7_75t_SL g625 ( 
.A(n_555),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_529),
.B(n_465),
.Y(n_626)
);

AND2x4_ASAP7_75t_SL g627 ( 
.A(n_555),
.B(n_497),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_535),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_577),
.A2(n_487),
.B1(n_497),
.B2(n_388),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_539),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_574),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_465),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_571),
.A2(n_393),
.B(n_399),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

OAI211xp5_ASAP7_75t_SL g636 ( 
.A1(n_544),
.A2(n_451),
.B(n_445),
.C(n_453),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_573),
.B(n_465),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_539),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_539),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_573),
.B(n_466),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_580),
.B(n_519),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_585),
.B(n_574),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_549),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_622),
.B(n_542),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_585),
.B(n_625),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_584),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_608),
.B(n_542),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_610),
.B(n_542),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_594),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_549),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_619),
.B(n_623),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_599),
.B(n_553),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_564),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_625),
.B(n_564),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_601),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_582),
.B(n_588),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_592),
.B(n_564),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_595),
.B(n_565),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_594),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_595),
.B(n_555),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_598),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_598),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_606),
.B(n_550),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_600),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_632),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_627),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_626),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_600),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_543),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_626),
.B(n_543),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_601),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_595),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_550),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_586),
.B(n_543),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_612),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_612),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_604),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_565),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_565),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_545),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_642),
.B(n_566),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_586),
.B(n_545),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_620),
.B(n_550),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_614),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_620),
.B(n_562),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_603),
.A2(n_553),
.B1(n_559),
.B2(n_531),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_618),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_602),
.B(n_554),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_602),
.B(n_554),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_591),
.B(n_536),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_587),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_614),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_624),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_604),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_602),
.B(n_557),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_642),
.B(n_566),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_587),
.B(n_566),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_668),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_644),
.B(n_627),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_649),
.B(n_590),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_690),
.B(n_591),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_SL g705 ( 
.A(n_668),
.B(n_632),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_672),
.B(n_590),
.Y(n_706)
);

INVx3_ASAP7_75t_SL g707 ( 
.A(n_669),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_691),
.B(n_597),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_692),
.B(n_591),
.Y(n_709)
);

NOR2x1p5_ASAP7_75t_L g710 ( 
.A(n_647),
.B(n_607),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_SL g711 ( 
.A(n_669),
.B(n_607),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_643),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_646),
.Y(n_713)
);

OAI221xp5_ASAP7_75t_L g714 ( 
.A1(n_689),
.A2(n_629),
.B1(n_599),
.B2(n_613),
.C(n_531),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_647),
.B(n_591),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_SL g716 ( 
.A(n_693),
.B(n_488),
.Y(n_716)
);

AO221x2_ASAP7_75t_L g717 ( 
.A1(n_698),
.A2(n_613),
.B1(n_576),
.B2(n_567),
.C(n_570),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_650),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_653),
.B(n_597),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_644),
.A2(n_499),
.B1(n_516),
.B2(n_553),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_663),
.B(n_632),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_654),
.A2(n_553),
.B1(n_559),
.B2(n_536),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_677),
.B(n_683),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_643),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_654),
.A2(n_559),
.B1(n_567),
.B2(n_541),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_685),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_654),
.A2(n_559),
.B1(n_541),
.B2(n_575),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_700),
.B(n_547),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_700),
.B(n_547),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_648),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_673),
.B(n_547),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_660),
.B(n_547),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_663),
.B(n_627),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_660),
.B(n_557),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_645),
.Y(n_735)
);

AO221x2_ASAP7_75t_L g736 ( 
.A1(n_648),
.A2(n_576),
.B1(n_651),
.B2(n_696),
.C(n_695),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_666),
.B(n_583),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_663),
.B(n_593),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_666),
.B(n_583),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_676),
.B(n_686),
.Y(n_740)
);

CKINVDCx8_ASAP7_75t_R g741 ( 
.A(n_663),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_SL g742 ( 
.A(n_659),
.B(n_523),
.Y(n_742)
);

OAI221xp5_ASAP7_75t_L g743 ( 
.A1(n_675),
.A2(n_581),
.B1(n_593),
.B2(n_569),
.C(n_570),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_651),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_676),
.B(n_518),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_686),
.A2(n_541),
.B1(n_575),
.B2(n_616),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_645),
.B(n_652),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_652),
.B(n_633),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_670),
.B(n_633),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_SL g750 ( 
.A1(n_655),
.A2(n_634),
.B(n_636),
.Y(n_750)
);

OAI221xp5_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_675),
.B1(n_581),
.B2(n_569),
.C(n_659),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_750),
.B(n_546),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_711),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_726),
.B(n_688),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_716),
.A2(n_717),
.B1(n_714),
.B2(n_736),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_713),
.B(n_688),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_707),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_740),
.B(n_662),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_712),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_724),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_710),
.B(n_675),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_701),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_730),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_718),
.B(n_655),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_744),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_736),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_733),
.B(n_656),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_722),
.B(n_662),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_733),
.B(n_656),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_747),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_721),
.B(n_694),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_735),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_717),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_742),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_715),
.B(n_694),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_705),
.B(n_699),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_737),
.B(n_664),
.Y(n_777)
);

NOR2x1_ASAP7_75t_L g778 ( 
.A(n_725),
.B(n_727),
.Y(n_778)
);

INVx3_ASAP7_75t_SL g779 ( 
.A(n_715),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_702),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_745),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_720),
.B(n_699),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_704),
.B(n_661),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_732),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_739),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_734),
.B(n_706),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_728),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_738),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_703),
.B(n_661),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_741),
.B(n_681),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_738),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_729),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_709),
.B(n_681),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_708),
.B(n_682),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_755),
.A2(n_746),
.B(n_743),
.Y(n_795)
);

OAI31xp33_ASAP7_75t_L g796 ( 
.A1(n_766),
.A2(n_719),
.A3(n_682),
.B(n_684),
.Y(n_796)
);

AOI222xp33_ASAP7_75t_L g797 ( 
.A1(n_773),
.A2(n_749),
.B1(n_731),
.B2(n_748),
.C1(n_556),
.C2(n_561),
.Y(n_797)
);

OAI21xp33_ASAP7_75t_L g798 ( 
.A1(n_778),
.A2(n_766),
.B(n_768),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_760),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_760),
.Y(n_800)
);

OAI321xp33_ASAP7_75t_L g801 ( 
.A1(n_752),
.A2(n_616),
.A3(n_537),
.B1(n_561),
.B2(n_556),
.C(n_617),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_762),
.B(n_684),
.Y(n_802)
);

NOR4xp25_ASAP7_75t_L g803 ( 
.A(n_751),
.B(n_664),
.C(n_696),
.D(n_695),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_757),
.B(n_578),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_763),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_SL g806 ( 
.A1(n_774),
.A2(n_671),
.B(n_687),
.C(n_665),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_763),
.Y(n_807)
);

NAND2x1_ASAP7_75t_L g808 ( 
.A(n_761),
.B(n_616),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_765),
.Y(n_809)
);

OA211x2_ASAP7_75t_L g810 ( 
.A1(n_776),
.A2(n_617),
.B(n_537),
.C(n_558),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_781),
.B(n_665),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_765),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_759),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_772),
.A2(n_678),
.B1(n_687),
.B2(n_667),
.C(n_679),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_768),
.A2(n_667),
.B(n_671),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_785),
.B(n_678),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_753),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_759),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_SL g819 ( 
.A(n_753),
.B(n_679),
.C(n_639),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_756),
.B(n_657),
.Y(n_820)
);

AOI322xp5_ASAP7_75t_L g821 ( 
.A1(n_778),
.A2(n_640),
.A3(n_637),
.B1(n_639),
.B2(n_635),
.C1(n_628),
.C2(n_624),
.Y(n_821)
);

OAI33xp33_ASAP7_75t_L g822 ( 
.A1(n_772),
.A2(n_635),
.A3(n_628),
.B1(n_589),
.B2(n_621),
.B3(n_596),
.Y(n_822)
);

OA21x2_ASAP7_75t_L g823 ( 
.A1(n_788),
.A2(n_680),
.B(n_674),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_759),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_791),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_SL g826 ( 
.A(n_782),
.B(n_697),
.C(n_680),
.Y(n_826)
);

AOI21xp33_ASAP7_75t_SL g827 ( 
.A1(n_752),
.A2(n_616),
.B(n_522),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_799),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_800),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_817),
.B(n_780),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_805),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_807),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_825),
.B(n_770),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_809),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_798),
.B(n_779),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_815),
.A2(n_752),
.B(n_761),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_795),
.B(n_779),
.Y(n_837)
);

NOR2x1_ASAP7_75t_L g838 ( 
.A(n_819),
.B(n_752),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_802),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_812),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_821),
.B(n_752),
.C(n_797),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_813),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_808),
.B(n_791),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_818),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_824),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_804),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_R g848 ( 
.A(n_827),
.B(n_790),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_820),
.B(n_779),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_816),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_823),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_803),
.B(n_770),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_826),
.B(n_764),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_823),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_796),
.B(n_767),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_814),
.B(n_767),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_810),
.B(n_769),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_826),
.B(n_769),
.Y(n_858)
);

XNOR2x1_ASAP7_75t_L g859 ( 
.A(n_801),
.B(n_790),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_843),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_845),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_846),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_828),
.Y(n_863)
);

INVxp33_ASAP7_75t_L g864 ( 
.A(n_835),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_829),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_831),
.Y(n_866)
);

INVx8_ASAP7_75t_L g867 ( 
.A(n_844),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_832),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_854),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_841),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_833),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_830),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_839),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_851),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_854),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_837),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_844),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_852),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_844),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_844),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_858),
.Y(n_882)
);

INVx3_ASAP7_75t_SL g883 ( 
.A(n_837),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_840),
.B(n_806),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_850),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_849),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_858),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_847),
.Y(n_888)
);

BUFx4f_ASAP7_75t_SL g889 ( 
.A(n_857),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_856),
.Y(n_890)
);

NAND4xp25_ASAP7_75t_SL g891 ( 
.A(n_879),
.B(n_842),
.C(n_838),
.D(n_836),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_884),
.A2(n_859),
.B(n_835),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_877),
.B(n_856),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_853),
.C(n_819),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_870),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_874),
.B(n_853),
.C(n_855),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_870),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_SL g898 ( 
.A(n_883),
.B(n_857),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_878),
.B(n_855),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_884),
.A2(n_859),
.B(n_848),
.C(n_788),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_L g901 ( 
.A1(n_890),
.A2(n_822),
.B1(n_848),
.B2(n_770),
.C(n_792),
.Y(n_901)
);

OAI211xp5_ASAP7_75t_SL g902 ( 
.A1(n_873),
.A2(n_788),
.B(n_792),
.C(n_787),
.Y(n_902)
);

NOR3x1_ASAP7_75t_L g903 ( 
.A(n_887),
.B(n_787),
.C(n_754),
.Y(n_903)
);

NOR4xp75_ASAP7_75t_L g904 ( 
.A(n_882),
.B(n_771),
.C(n_783),
.D(n_786),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_878),
.B(n_771),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_882),
.B(n_793),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_SL g907 ( 
.A(n_864),
.B(n_775),
.C(n_758),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_SL g908 ( 
.A1(n_886),
.A2(n_784),
.B1(n_775),
.B2(n_794),
.C(n_758),
.Y(n_908)
);

NOR3x1_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_784),
.C(n_777),
.Y(n_909)
);

AOI222xp33_ASAP7_75t_L g910 ( 
.A1(n_889),
.A2(n_864),
.B1(n_883),
.B2(n_872),
.C1(n_867),
.C2(n_878),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_880),
.B(n_793),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_900),
.A2(n_867),
.B(n_878),
.C(n_880),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_892),
.A2(n_896),
.B(n_910),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_895),
.Y(n_914)
);

AOI211xp5_ASAP7_75t_L g915 ( 
.A1(n_891),
.A2(n_881),
.B(n_876),
.C(n_875),
.Y(n_915)
);

AOI211xp5_ASAP7_75t_L g916 ( 
.A1(n_894),
.A2(n_899),
.B(n_898),
.C(n_905),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_897),
.Y(n_917)
);

AO22x2_ASAP7_75t_L g918 ( 
.A1(n_894),
.A2(n_881),
.B1(n_893),
.B2(n_866),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_904),
.B(n_876),
.C(n_863),
.Y(n_919)
);

NOR2x1_ASAP7_75t_L g920 ( 
.A(n_907),
.B(n_860),
.Y(n_920)
);

XNOR2xp5_ASAP7_75t_L g921 ( 
.A(n_911),
.B(n_865),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_901),
.A2(n_871),
.B(n_869),
.Y(n_922)
);

AOI222xp33_ASAP7_75t_L g923 ( 
.A1(n_906),
.A2(n_889),
.B1(n_867),
.B2(n_868),
.C1(n_862),
.C2(n_861),
.Y(n_923)
);

INVx4_ASAP7_75t_SL g924 ( 
.A(n_909),
.Y(n_924)
);

AOI211xp5_ASAP7_75t_SL g925 ( 
.A1(n_902),
.A2(n_777),
.B(n_794),
.C(n_789),
.Y(n_925)
);

OAI221xp5_ASAP7_75t_L g926 ( 
.A1(n_908),
.A2(n_822),
.B1(n_546),
.B2(n_616),
.C(n_657),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_903),
.B(n_697),
.Y(n_927)
);

OAI221xp5_ASAP7_75t_SL g928 ( 
.A1(n_900),
.A2(n_578),
.B1(n_579),
.B2(n_674),
.C(n_658),
.Y(n_928)
);

AOI221xp5_ASAP7_75t_L g929 ( 
.A1(n_891),
.A2(n_658),
.B1(n_615),
.B2(n_638),
.C(n_605),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_924),
.B(n_920),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_917),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_914),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_921),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_916),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_918),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_918),
.B(n_922),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_SL g937 ( 
.A1(n_915),
.A2(n_395),
.B1(n_638),
.B2(n_630),
.C(n_604),
.Y(n_937)
);

XOR2xp5_ASAP7_75t_L g938 ( 
.A(n_919),
.B(n_927),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_924),
.Y(n_939)
);

AO211x2_ASAP7_75t_L g940 ( 
.A1(n_913),
.A2(n_540),
.B(n_560),
.C(n_558),
.Y(n_940)
);

NAND2x1p5_ASAP7_75t_L g941 ( 
.A(n_923),
.B(n_912),
.Y(n_941)
);

XNOR2xp5_ASAP7_75t_L g942 ( 
.A(n_929),
.B(n_926),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_928),
.B(n_489),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_930),
.B(n_925),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_939),
.B(n_398),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_SL g946 ( 
.A(n_936),
.B(n_560),
.C(n_540),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_934),
.B(n_605),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_933),
.B(n_398),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_935),
.B(n_605),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_SL g950 ( 
.A(n_936),
.B(n_495),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_932),
.B(n_398),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_SL g952 ( 
.A(n_931),
.B(n_489),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_SL g953 ( 
.A1(n_944),
.A2(n_938),
.B1(n_941),
.B2(n_942),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_947),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_949),
.B(n_941),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_950),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_945),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_952),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_946),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_955),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_956),
.A2(n_937),
.B(n_943),
.C(n_940),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_958),
.B(n_937),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_954),
.A2(n_948),
.B(n_951),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_960),
.B(n_959),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_962),
.A2(n_953),
.B1(n_957),
.B2(n_492),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_964),
.A2(n_963),
.B1(n_961),
.B2(n_495),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_L g967 ( 
.A1(n_966),
.A2(n_965),
.B(n_609),
.Y(n_967)
);

OAI22x1_ASAP7_75t_L g968 ( 
.A1(n_967),
.A2(n_492),
.B1(n_638),
.B2(n_615),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_968),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_969),
.A2(n_615),
.B1(n_630),
.B2(n_534),
.C(n_562),
.Y(n_970)
);

AOI211xp5_ASAP7_75t_L g971 ( 
.A1(n_970),
.A2(n_630),
.B(n_596),
.C(n_611),
.Y(n_971)
);


endmodule