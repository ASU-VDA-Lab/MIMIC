module fake_jpeg_30929_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_1),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_63),
.B(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_85),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_82),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_47),
.B1(n_54),
.B2(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_59),
.B1(n_62),
.B2(n_61),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_24),
.B(n_44),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_49),
.B1(n_54),
.B2(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_60),
.B1(n_50),
.B2(n_58),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_12),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_1),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_5),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_5),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_6),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_27),
.B(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_7),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OR2x4_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_26),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_97),
.B(n_37),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_79),
.B1(n_9),
.B2(n_10),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_112),
.B1(n_120),
.B2(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_13),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_34),
.B1(n_40),
.B2(n_39),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_12),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_13),
.C(n_14),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_18),
.B1(n_38),
.B2(n_16),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_126),
.Y(n_136)
);

XOR2x1_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_116),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_129),
.B(n_132),
.Y(n_141)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_105),
.CON(n_129),
.SN(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_120),
.Y(n_138)
);

CKINVDCx10_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_135),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_17),
.B1(n_36),
.B2(n_41),
.Y(n_134)
);

AOI22x1_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_112),
.B1(n_118),
.B2(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_148),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_140),
.C(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_149),
.C(n_151),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_136),
.B(n_128),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_123),
.Y(n_157)
);


endmodule