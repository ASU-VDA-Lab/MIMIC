module fake_jpeg_8356_n_100 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_12),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_11),
.B(n_19),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_32),
.A3(n_36),
.B1(n_12),
.B2(n_19),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_20),
.B1(n_14),
.B2(n_11),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_21),
.A2(n_20),
.B1(n_14),
.B2(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_49),
.B(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_31),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_15),
.B(n_19),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_23),
.C(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_45),
.B1(n_41),
.B2(n_46),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_16),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_48),
.B1(n_39),
.B2(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_23),
.B(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_22),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_59),
.C(n_55),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_74),
.C(n_77),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_54),
.C(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_69),
.B1(n_63),
.B2(n_62),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_54),
.C(n_50),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_66),
.A3(n_71),
.B1(n_51),
.B2(n_24),
.C1(n_27),
.C2(n_9),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_2),
.C(n_3),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_1),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_42),
.B1(n_24),
.B2(n_9),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_82),
.B(n_0),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_79),
.B(n_81),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_81),
.C(n_6),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.C(n_89),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_93),
.C(n_7),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_4),
.B(n_8),
.Y(n_99)
);


endmodule