module fake_jpeg_20309_n_229 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.C(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_31),
.B1(n_14),
.B2(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_20),
.B1(n_18),
.B2(n_30),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_53),
.B1(n_35),
.B2(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_26),
.CI(n_15),
.CON(n_48),
.SN(n_48)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_31),
.B1(n_37),
.B2(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_33),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_69),
.B1(n_37),
.B2(n_33),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_35),
.C(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_53),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_35),
.B(n_25),
.C(n_24),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_58),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_53),
.B(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_49),
.B1(n_33),
.B2(n_37),
.Y(n_82)
);

AND2x4_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_69),
.B1(n_70),
.B2(n_33),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_71),
.B1(n_78),
.B2(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_89),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_88),
.B(n_40),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_53),
.B(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_16),
.C(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_76),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_85),
.B1(n_82),
.B2(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_63),
.C(n_70),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_77),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_118),
.B1(n_41),
.B2(n_40),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_62),
.C(n_65),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_85),
.C(n_81),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_93),
.B(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_93),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_61),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_33),
.B1(n_75),
.B2(n_61),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_125),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_137),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_112),
.B1(n_103),
.B2(n_101),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_129),
.B1(n_138),
.B2(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_21),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_88),
.B1(n_82),
.B2(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_88),
.C(n_79),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_110),
.B(n_111),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_18),
.A3(n_40),
.B1(n_56),
.B2(n_54),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_111),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_10),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_75),
.B1(n_47),
.B2(n_45),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_109),
.B1(n_104),
.B2(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_133),
.B1(n_134),
.B2(n_142),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_29),
.C(n_28),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_40),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_118),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_150),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_163),
.B1(n_133),
.B2(n_122),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_101),
.B(n_103),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_161),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_103),
.B(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_139),
.B1(n_120),
.B2(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_23),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_28),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_21),
.B(n_16),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_134),
.B1(n_127),
.B2(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_143),
.C(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_153),
.B1(n_146),
.B2(n_155),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_141),
.C(n_29),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_157),
.C(n_149),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_28),
.C(n_29),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_176),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_151),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_147),
.B(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_57),
.B1(n_3),
.B2(n_4),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_155),
.B1(n_162),
.B2(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_185),
.B1(n_167),
.B2(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_174),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_50),
.B1(n_41),
.B2(n_29),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_166),
.C(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_178),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_57),
.C(n_41),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_198),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_57),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_199),
.B(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_207),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_12),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_182),
.B1(n_189),
.B2(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_41),
.C(n_12),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_189),
.B(n_196),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_206),
.A2(n_197),
.B(n_5),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_213),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_214),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_13),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_202),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_13),
.B(n_6),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_206),
.B(n_19),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_19),
.B(n_6),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_223),
.B(n_224),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_0),
.B(n_6),
.C(n_7),
.Y(n_224)
);

NAND4xp25_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_217),
.C(n_221),
.D(n_218),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_0),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_13),
.C2(n_225),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_7),
.B(n_8),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_7),
.Y(n_229)
);


endmodule