module fake_jpeg_2917_n_397 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_70),
.Y(n_111)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_55),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_56),
.B(n_79),
.Y(n_154)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_0),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_95),
.Y(n_134)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_20),
.B(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_27),
.B(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_5),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_R g123 ( 
.A(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_6),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_81),
.B(n_88),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_9),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_82),
.B(n_87),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_21),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g141 ( 
.A(n_84),
.Y(n_141)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_11),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_15),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_46),
.Y(n_91)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_15),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_100),
.Y(n_153)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_26),
.B(n_18),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_38),
.B(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_106),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_18),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_32),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_52),
.B1(n_26),
.B2(n_34),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_116),
.A2(n_118),
.B1(n_130),
.B2(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_32),
.B1(n_34),
.B2(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_56),
.B(n_15),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_59),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_140),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_81),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_108),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_61),
.A2(n_29),
.B1(n_39),
.B2(n_41),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_157),
.A2(n_142),
.B1(n_137),
.B2(n_146),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_33),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_48),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_173),
.Y(n_180)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_48),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_62),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_76),
.A2(n_77),
.B(n_110),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_157),
.B(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_182),
.B(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_183),
.B(n_192),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

AO22x1_ASAP7_75t_SL g185 ( 
.A1(n_134),
.A2(n_63),
.B1(n_64),
.B2(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_113),
.Y(n_186)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_114),
.B(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_189),
.B(n_191),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_134),
.A2(n_160),
.B(n_154),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_193),
.B(n_178),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_135),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_193),
.B(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_158),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_196),
.Y(n_241)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_129),
.C(n_138),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_214),
.C(n_179),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_144),
.B(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_202),
.Y(n_235)
);

OR2x4_ASAP7_75t_L g200 ( 
.A(n_127),
.B(n_141),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_231),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_170),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_121),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_213),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_112),
.A2(n_148),
.B1(n_164),
.B2(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_204),
.A2(n_215),
.B1(n_220),
.B2(n_200),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_150),
.B(n_151),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_208),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_150),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_112),
.A2(n_152),
.B1(n_159),
.B2(n_124),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_209),
.A2(n_197),
.B1(n_184),
.B2(n_201),
.Y(n_271)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_211),
.Y(n_268)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_124),
.B(n_162),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_148),
.A2(n_161),
.B1(n_165),
.B2(n_136),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_139),
.B(n_126),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_132),
.B(n_172),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_136),
.A2(n_143),
.B1(n_167),
.B2(n_127),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_221),
.A2(n_204),
.B1(n_211),
.B2(n_224),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_142),
.B(n_146),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_120),
.B(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_230),
.Y(n_232)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_228),
.Y(n_270)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_229),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_185),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_256),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_251),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_253),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_180),
.B(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_177),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_252),
.B(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_210),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_196),
.A2(n_212),
.B(n_221),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_188),
.B(n_216),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_220),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_253),
.B(n_258),
.Y(n_293)
);

AOI32xp33_ASAP7_75t_L g264 ( 
.A1(n_195),
.A2(n_206),
.A3(n_225),
.B1(n_205),
.B2(n_215),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_258),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_260),
.B1(n_232),
.B2(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_226),
.C(n_230),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_300),
.C(n_303),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_285),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_187),
.B1(n_228),
.B2(n_254),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_278),
.B1(n_287),
.B2(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_246),
.B1(n_240),
.B2(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_288),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_241),
.A2(n_232),
.B1(n_258),
.B2(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_294),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_259),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_260),
.B(n_247),
.Y(n_311)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_266),
.B(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_243),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_244),
.C(n_252),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_261),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_310),
.B(n_303),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_314),
.B(n_318),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_278),
.B(n_281),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_275),
.A2(n_235),
.B(n_236),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_276),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_264),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_262),
.B(n_247),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_322),
.A2(n_324),
.B(n_302),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_270),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_300),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_296),
.B(n_301),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_272),
.C(n_270),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_273),
.C(n_290),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_334),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_327),
.B(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_304),
.B(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_335),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_336),
.C(n_339),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_289),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_309),
.B(n_297),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_325),
.C(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_310),
.B(n_266),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_315),
.Y(n_338)
);

INVx13_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_296),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_320),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_340),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_343),
.B1(n_316),
.B2(n_318),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_316),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_307),
.A2(n_269),
.B1(n_284),
.B2(n_295),
.Y(n_343)
);

XNOR2x2_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_307),
.Y(n_345)
);

AOI21xp33_ASAP7_75t_SL g367 ( 
.A1(n_345),
.A2(n_328),
.B(n_317),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_341),
.A2(n_324),
.B(n_311),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_349),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_348),
.A2(n_342),
.B1(n_329),
.B2(n_338),
.Y(n_359)
);

NOR3xp33_ASAP7_75t_SL g349 ( 
.A(n_330),
.B(n_304),
.C(n_306),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_355),
.A2(n_316),
.B(n_344),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_361),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_367),
.B(n_355),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_347),
.A2(n_343),
.B1(n_335),
.B2(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_368),
.Y(n_371)
);

AOI321xp33_ASAP7_75t_L g363 ( 
.A1(n_356),
.A2(n_322),
.A3(n_313),
.B1(n_339),
.B2(n_327),
.C(n_340),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_348),
.A2(n_332),
.B1(n_334),
.B2(n_319),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_364),
.B(n_366),
.Y(n_375)
);

OAI322xp33_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_326),
.A3(n_313),
.B1(n_337),
.B2(n_306),
.C1(n_336),
.C2(n_331),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_346),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_312),
.B1(n_308),
.B2(n_317),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_357),
.C(n_352),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_376),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_374),
.B(n_320),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_351),
.B(n_345),
.C(n_349),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_357),
.C(n_352),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_372),
.A2(n_361),
.B(n_354),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_378),
.A2(n_380),
.B(n_382),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_368),
.C(n_321),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_381),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_375),
.A2(n_363),
.B(n_350),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_350),
.Y(n_381)
);

NAND4xp25_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_321),
.C(n_353),
.D(n_312),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_383),
.A2(n_381),
.B(n_379),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_373),
.C(n_371),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_234),
.C(n_250),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_245),
.Y(n_390)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_377),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_245),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_391),
.B(n_387),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_392),
.B1(n_250),
.B2(n_265),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g391 ( 
.A(n_384),
.B(n_234),
.CI(n_272),
.CON(n_391),
.SN(n_391)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_390),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_392),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_396),
.Y(n_397)
);


endmodule