module fake_netlist_1_5087_n_461 (n_20, n_12, n_56, n_47, n_52, n_67, n_50, n_7, n_1, n_60, n_16, n_22, n_3, n_19, n_10, n_34, n_40, n_68, n_25, n_30, n_36, n_9, n_13, n_53, n_26, n_11, n_64, n_69, n_39, n_43, n_62, n_38, n_23, n_0, n_33, n_4, n_59, n_24, n_35, n_6, n_32, n_8, n_15, n_57, n_61, n_51, n_44, n_66, n_70, n_46, n_45, n_42, n_21, n_2, n_37, n_48, n_27, n_63, n_18, n_17, n_54, n_28, n_41, n_58, n_65, n_55, n_49, n_5, n_29, n_14, n_31, n_461, n_501);
input n_20;
input n_12;
input n_56;
input n_47;
input n_52;
input n_67;
input n_50;
input n_7;
input n_1;
input n_60;
input n_16;
input n_22;
input n_3;
input n_19;
input n_10;
input n_34;
input n_40;
input n_68;
input n_25;
input n_30;
input n_36;
input n_9;
input n_13;
input n_53;
input n_26;
input n_11;
input n_64;
input n_69;
input n_39;
input n_43;
input n_62;
input n_38;
input n_23;
input n_0;
input n_33;
input n_4;
input n_59;
input n_24;
input n_35;
input n_6;
input n_32;
input n_8;
input n_15;
input n_57;
input n_61;
input n_51;
input n_44;
input n_66;
input n_70;
input n_46;
input n_45;
input n_42;
input n_21;
input n_2;
input n_37;
input n_48;
input n_27;
input n_63;
input n_18;
input n_17;
input n_54;
input n_28;
input n_41;
input n_58;
input n_65;
input n_55;
input n_49;
input n_5;
input n_29;
input n_14;
input n_31;
output n_461;
output n_501;
wire n_107;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_180;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_357;
wire n_74;
wire n_308;
wire n_44;
wire n_394;
wire n_189;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_316;
wire n_285;
wire n_471;
wire n_47;
wire n_475;
wire n_281;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_368;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_176;
wire n_436;
wire n_438;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_223;
wire n_405;
wire n_19;
wire n_409;
wire n_482;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_303;
wire n_468;
wire n_159;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_378;
wire n_246;
wire n_191;
wire n_143;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_135;
wire n_481;
wire n_315;
wire n_397;
wire n_53;
wire n_213;
wire n_196;
wire n_293;
wire n_127;
wire n_312;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_186;
wire n_137;
wire n_334;
wire n_164;
wire n_433;
wire n_120;
wire n_392;
wire n_155;
wire n_162;
wire n_114;
wire n_50;
wire n_3;
wire n_331;
wire n_330;
wire n_231;
wire n_9;
wire n_428;
wire n_178;
wire n_478;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_329;
wire n_6;
wire n_8;
wire n_187;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_441;
wire n_425;
wire n_314;
wire n_307;
wire n_215;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_351;
wire n_1;
wire n_16;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_228;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_362;
wire n_485;
wire n_396;
wire n_354;
wire n_152;
wire n_70;
wire n_458;
wire n_375;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_491;
wire n_388;
wire n_266;
wire n_80;
wire n_326;
wire n_275;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_38;
wire n_272;
wire n_100;
wire n_299;
wire n_280;
wire n_141;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_193;
wire n_232;
wire n_344;
wire n_147;
wire n_185;
wire n_367;
wire n_267;
wire n_171;
wire n_450;
wire n_140;
wire n_111;
wire n_212;
wire n_30;
wire n_13;
wire n_254;
wire n_435;
wire n_64;
wire n_69;
wire n_248;
wire n_407;
wire n_83;
wire n_200;
wire n_262;
wire n_119;
wire n_339;
wire n_347;
wire n_124;
wire n_79;
wire n_129;
wire n_157;
wire n_103;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_273;
wire n_325;
wire n_163;
wire n_348;
wire n_96;
wire n_72;
wire n_77;
wire n_90;
wire n_214;
wire n_167;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_413;
wire n_65;
wire n_5;
wire n_496;
wire n_393;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_290;
wire n_217;
wire n_201;
wire n_277;
wire n_259;
wire n_244;
wire n_276;
wire n_297;
wire n_225;
wire n_350;
wire n_208;
wire n_419;
wire n_252;
wire n_168;
wire n_271;
wire n_94;
wire n_194;
wire n_282;
wire n_58;
wire n_113;
wire n_242;
wire n_498;
wire n_284;
wire n_321;
wire n_302;
wire n_116;
wire n_292;
wire n_118;
wire n_233;
wire n_257;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_146;
wire n_337;
wire n_32;
wire n_93;
wire n_406;
wire n_372;
wire n_467;
wire n_41;
wire n_417;
wire n_451;
wire n_445;
wire n_500;
wire n_10;
wire n_390;
wire n_75;
wire n_82;
wire n_183;
wire n_132;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_360;
wire n_363;
wire n_427;
wire n_106;
wire n_296;
wire n_42;
wire n_21;
wire n_437;
wire n_89;
wire n_480;
wire n_130;
wire n_310;
wire n_341;
wire n_14;
wire n_236;
wire n_136;
wire n_260;
wire n_222;
wire n_381;
wire n_34;
wire n_142;
wire n_385;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_268;
wire n_190;
wire n_62;
wire n_4;
wire n_59;
wire n_323;
wire n_376;
wire n_240;
wire n_459;
wire n_88;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_380;
wire n_87;
wire n_466;
wire n_349;
wire n_207;
wire n_197;
wire n_81;
wire n_298;
wire n_112;
wire n_78;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_36;
wire n_416;
wire n_432;
wire n_465;
wire n_414;
wire n_369;
wire n_469;
wire n_361;
wire n_237;
wire n_15;
wire n_429;
wire n_256;
wire n_398;
wire n_117;
wire n_238;
wire n_365;
wire n_294;
wire n_2;
wire n_338;
wire n_391;
wire n_209;
wire n_241;
wire n_20;
wire n_84;
wire n_449;
wire n_12;
wire n_56;
wire n_412;
wire n_455;
wire n_67;
wire n_456;
wire n_22;
wire n_479;
wire n_311;
wire n_401;
wire n_383;
wire n_202;
wire n_319;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_486;
wire n_24;
wire n_35;
wire n_472;
wire n_490;
wire n_400;
wire n_457;
wire n_134;
wire n_48;
wire n_255;
wire n_55;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_488;
wire n_382;
wire n_60;
wire n_138;
wire n_462;
wire n_474;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_92;
wire n_313;
wire n_333;
wire n_358;
wire n_175;
wire n_128;
wire n_306;
wire n_415;
wire n_0;
wire n_258;
wire n_234;
wire n_184;
wire n_265;
wire n_57;
wire n_51;
wire n_411;
wire n_287;
wire n_144;
wire n_403;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_177;
wire n_28;
wire n_448;
wire n_49;
wire n_206;
wire n_31;
INVx1_ASAP7_75t_L g71 ( .A(n_17), .Y(n_71) );
INVx2_ASAP7_75t_L g72 ( .A(n_51), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_29), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_47), .Y(n_74) );
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_42), .Y(n_75) );
CKINVDCx14_ASAP7_75t_R g76 ( .A(n_19), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_15), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_66), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_45), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_46), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_50), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
BUFx2_ASAP7_75t_L g83 ( .A(n_39), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_20), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_17), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_36), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_61), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_37), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_23), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_25), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
NOR2xp67_ASAP7_75t_L g93 ( .A(n_63), .B(n_10), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_11), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_4), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_55), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_1), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_24), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_30), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_62), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_77), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_77), .Y(n_107) );
AND3x2_ASAP7_75t_L g108 ( .A(n_83), .B(n_0), .C(n_1), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_83), .B(n_0), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_92), .B(n_2), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_103), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_103), .B(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_95), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_75), .B(n_3), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_98), .B(n_5), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_85), .B(n_6), .Y(n_121) );
NAND2xp33_ASAP7_75t_R g122 ( .A(n_74), .B(n_33), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_97), .Y(n_125) );
NAND2xp33_ASAP7_75t_L g126 ( .A(n_103), .B(n_34), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_75), .B(n_6), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_121), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
NOR2x1p5_ASAP7_75t_L g130 ( .A(n_111), .B(n_95), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_124), .B(n_76), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_105), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_110), .B(n_71), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_105), .Y(n_136) );
NAND2xp33_ASAP7_75t_L g137 ( .A(n_110), .B(n_103), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_124), .B(n_101), .Y(n_138) );
OR2x2_ASAP7_75t_SL g139 ( .A(n_111), .B(n_71), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_121), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_113), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_121), .B(n_82), .Y(n_143) );
AO22x2_ASAP7_75t_L g144 ( .A1(n_121), .A2(n_104), .B1(n_102), .B2(n_73), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_127), .B(n_104), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_118), .B(n_101), .Y(n_147) );
INVx1_ASAP7_75t_SL g148 ( .A(n_127), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_109), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_117), .B(n_89), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_118), .B(n_89), .Y(n_152) );
NAND2x1p5_ASAP7_75t_L g153 ( .A(n_117), .B(n_90), .Y(n_153) );
INVx2_ASAP7_75t_SL g154 ( .A(n_130), .Y(n_154) );
AOI22xp5_ASAP7_75t_SL g155 ( .A1(n_148), .A2(n_91), .B1(n_81), .B2(n_120), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_131), .B(n_120), .Y(n_156) );
OR2x4_ASAP7_75t_L g157 ( .A(n_139), .B(n_82), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx1_ASAP7_75t_SL g159 ( .A(n_145), .Y(n_159) );
INVxp33_ASAP7_75t_SL g160 ( .A(n_144), .Y(n_160) );
AND2x6_ASAP7_75t_L g161 ( .A(n_128), .B(n_78), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_134), .B(n_78), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_134), .B(n_118), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_140), .B(n_79), .Y(n_165) );
AND2x4_ASAP7_75t_SL g166 ( .A(n_134), .B(n_94), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_145), .B(n_100), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_151), .B(n_108), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_136), .A2(n_112), .B(n_125), .C(n_123), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_151), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_135), .A2(n_99), .B1(n_94), .B2(n_107), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_153), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
BUFx5_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_153), .B(n_106), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_153), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_144), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_144), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_160), .A2(n_144), .B1(n_139), .B2(n_150), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_178), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_184), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_184), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_175), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_151), .B1(n_137), .B2(n_152), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_168), .B(n_149), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_170), .B(n_141), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_168), .B(n_108), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_168), .B(n_93), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_186), .A2(n_137), .B1(n_116), .B2(n_138), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_185), .A2(n_141), .B1(n_112), .B2(n_125), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_154), .B(n_116), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_164), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_181), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_172), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_172), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_166), .Y(n_216) );
BUFx8_ASAP7_75t_SL g217 ( .A(n_173), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_114), .B1(n_147), .B2(n_99), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_195), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_206), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_206), .B(n_179), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_216), .B(n_183), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_190), .A2(n_156), .B(n_163), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_193), .B(n_166), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_187), .A2(n_165), .B1(n_161), .B2(n_181), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_193), .B(n_182), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_187), .A2(n_161), .B1(n_165), .B2(n_162), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_207), .A2(n_177), .B(n_174), .C(n_162), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_209), .B(n_176), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_188), .B(n_177), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_190), .A2(n_174), .B(n_171), .C(n_88), .Y(n_234) );
INVxp33_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_196), .B(n_181), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_191), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_191), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_189), .Y(n_240) );
NAND2x1p5_ASAP7_75t_L g241 ( .A(n_212), .B(n_175), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_203), .A2(n_165), .B1(n_161), .B2(n_181), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_196), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_227), .A2(n_203), .B1(n_230), .B2(n_243), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g247 ( .A1(n_230), .A2(n_157), .B1(n_194), .B2(n_212), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_244), .B(n_212), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_244), .B(n_212), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g251 ( .A1(n_231), .A2(n_194), .B1(n_218), .B2(n_213), .C(n_210), .Y(n_251) );
OAI33xp33_ASAP7_75t_L g252 ( .A1(n_233), .A2(n_115), .A3(n_106), .B1(n_107), .B2(n_119), .B3(n_123), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_226), .A2(n_199), .B(n_201), .C(n_198), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_226), .A2(n_192), .B(n_197), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_233), .A2(n_199), .B1(n_204), .B2(n_210), .C(n_213), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_227), .A2(n_199), .B1(n_165), .B2(n_161), .Y(n_256) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_221), .A2(n_198), .B1(n_165), .B2(n_161), .C1(n_199), .C2(n_119), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_198), .B1(n_181), .B2(n_201), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_204), .B1(n_176), .B2(n_157), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_195), .B1(n_112), .B2(n_125), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_221), .A2(n_198), .B1(n_115), .B2(n_214), .C(n_215), .Y(n_262) );
AOI211xp5_ASAP7_75t_L g263 ( .A1(n_223), .A2(n_93), .B(n_88), .C(n_90), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_245), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_258), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_264), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_246), .A2(n_245), .B1(n_227), .B2(n_220), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_247), .A2(n_224), .B1(n_220), .B2(n_235), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
OAI31xp33_ASAP7_75t_L g273 ( .A1(n_260), .A2(n_225), .A3(n_232), .B(n_242), .Y(n_273) );
OAI221xp5_ASAP7_75t_L g274 ( .A1(n_263), .A2(n_242), .B1(n_220), .B2(n_234), .C(n_241), .Y(n_274) );
NAND2x1p5_ASAP7_75t_SL g275 ( .A(n_248), .B(n_222), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_254), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_249), .B(n_239), .Y(n_277) );
OAI322xp33_ASAP7_75t_L g278 ( .A1(n_265), .A2(n_79), .A3(n_96), .B1(n_102), .B2(n_86), .C1(n_80), .C2(n_97), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_249), .B(n_239), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_260), .A2(n_229), .B1(n_232), .B2(n_220), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_266), .B(n_222), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_256), .A2(n_229), .B1(n_232), .B2(n_238), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_250), .B(n_238), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_282), .Y(n_289) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_269), .B(n_266), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g291 ( .A(n_273), .B(n_263), .C(n_261), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_271), .A2(n_252), .B1(n_257), .B2(n_251), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_284), .A2(n_253), .B1(n_261), .B2(n_255), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
NAND2x1p5_ASAP7_75t_SL g295 ( .A(n_288), .B(n_250), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_269), .B(n_238), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_284), .A2(n_257), .B1(n_232), .B2(n_262), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_288), .B(n_80), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_267), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_272), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_274), .B(n_103), .C(n_96), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_276), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_281), .B(n_229), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_277), .B(n_229), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_279), .B(n_97), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_278), .B(n_240), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_279), .B(n_103), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_268), .B(n_236), .Y(n_310) );
AO211x2_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_7), .B(n_8), .C(n_9), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_283), .B(n_241), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_268), .B(n_236), .Y(n_313) );
OAI31xp33_ASAP7_75t_L g314 ( .A1(n_270), .A2(n_241), .A3(n_259), .B(n_84), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
OAI211xp5_ASAP7_75t_L g317 ( .A1(n_269), .A2(n_87), .B(n_215), .C(n_214), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_295), .B(n_275), .Y(n_319) );
NOR2xp67_ASAP7_75t_L g320 ( .A(n_302), .B(n_269), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_295), .B(n_285), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_280), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_303), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_315), .B(n_282), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_294), .B(n_299), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_307), .B(n_278), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_286), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_300), .B(n_286), .Y(n_329) );
NOR3xp33_ASAP7_75t_SL g330 ( .A(n_291), .B(n_122), .C(n_287), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_282), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_301), .B(n_309), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
NAND5xp2_ASAP7_75t_L g334 ( .A(n_297), .B(n_7), .C(n_8), .D(n_10), .E(n_11), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_285), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_315), .B(n_113), .Y(n_337) );
OAI332xp33_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .C1(n_18), .C2(n_19), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_298), .B(n_12), .Y(n_339) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_290), .B(n_211), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_298), .B(n_13), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_316), .B(n_113), .Y(n_342) );
NAND4xp25_ASAP7_75t_L g343 ( .A(n_291), .B(n_14), .C(n_16), .D(n_18), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
BUFx2_ASAP7_75t_SL g345 ( .A(n_296), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_316), .B(n_113), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_295), .B(n_219), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_308), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_306), .B(n_219), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_292), .A2(n_181), .B1(n_192), .B2(n_197), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_318), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_289), .B(n_180), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_296), .B(n_21), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_306), .B(n_22), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
OAI31xp33_ASAP7_75t_SL g360 ( .A1(n_302), .A2(n_197), .A3(n_192), .B(n_27), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_332), .B(n_304), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
NOR2xp67_ASAP7_75t_SL g363 ( .A(n_345), .B(n_317), .Y(n_363) );
OAI32xp33_ASAP7_75t_L g364 ( .A1(n_343), .A2(n_312), .A3(n_305), .B1(n_311), .B2(n_310), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_328), .B(n_290), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_325), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_332), .B(n_313), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_336), .B(n_313), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_336), .B(n_310), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_328), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_360), .A2(n_312), .B(n_126), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_359), .B(n_314), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_359), .B(n_311), .Y(n_375) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_343), .A2(n_211), .B(n_202), .C(n_205), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_320), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_333), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_328), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_335), .B(n_26), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_321), .B(n_28), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_328), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_327), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_335), .B(n_31), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_329), .B(n_32), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_345), .B(n_38), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_331), .B(n_40), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_323), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_338), .A2(n_133), .B1(n_142), .B2(n_146), .C(n_208), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_338), .B(n_41), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_331), .B(n_43), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_321), .B(n_44), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_324), .B(n_48), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_322), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_326), .B(n_49), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_344), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_344), .Y(n_397) );
XOR2x2_ASAP7_75t_L g398 ( .A(n_320), .B(n_53), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_360), .B(n_133), .C(n_142), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_334), .B(n_202), .C(n_211), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_324), .B(n_54), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_324), .B(n_56), .Y(n_402) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_340), .B(n_211), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_334), .B(n_57), .Y(n_404) );
NOR2xp33_ASAP7_75t_R g405 ( .A(n_319), .B(n_58), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_340), .A2(n_202), .B(n_208), .Y(n_406) );
INVxp67_ASAP7_75t_R g407 ( .A(n_386), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_362), .Y(n_408) );
OAI32xp33_ASAP7_75t_L g409 ( .A1(n_377), .A2(n_319), .A3(n_357), .B1(n_349), .B2(n_339), .Y(n_409) );
XNOR2x1_ASAP7_75t_L g410 ( .A(n_398), .B(n_357), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g412 ( .A1(n_389), .A2(n_341), .B(n_330), .C(n_353), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_370), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_372), .Y(n_416) );
XOR2x2_ASAP7_75t_L g417 ( .A(n_398), .B(n_358), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_395), .B(n_349), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
XNOR2xp5_ASAP7_75t_L g420 ( .A(n_367), .B(n_358), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_399), .A2(n_353), .B(n_342), .Y(n_421) );
AND2x2_ASAP7_75t_SL g422 ( .A(n_365), .B(n_337), .Y(n_422) );
AOI211x1_ASAP7_75t_L g423 ( .A1(n_364), .A2(n_342), .B(n_347), .C(n_351), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_379), .B(n_352), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_394), .B(n_352), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_361), .B(n_350), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
NOR3xp33_ASAP7_75t_SL g429 ( .A(n_390), .B(n_346), .C(n_354), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_377), .A2(n_354), .B(n_346), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_405), .A2(n_390), .B(n_375), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_403), .B(n_355), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_404), .B(n_356), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_382), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_363), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
BUFx12f_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_365), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_404), .A2(n_355), .B(n_356), .Y(n_440) );
AOI21xp33_ASAP7_75t_SL g441 ( .A1(n_381), .A2(n_348), .B(n_65), .Y(n_441) );
XNOR2x1_ASAP7_75t_L g442 ( .A(n_402), .B(n_348), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_405), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_373), .B(n_64), .Y(n_444) );
AOI21xp33_ASAP7_75t_SL g445 ( .A1(n_392), .A2(n_67), .B(n_69), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_400), .A2(n_202), .B(n_205), .Y(n_446) );
OAI221xp5_ASAP7_75t_SL g447 ( .A1(n_371), .A2(n_200), .B1(n_205), .B2(n_146), .C(n_133), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_400), .A2(n_200), .B(n_180), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_391), .Y(n_449) );
OAI31xp33_ASAP7_75t_L g450 ( .A1(n_401), .A2(n_200), .A3(n_146), .B(n_142), .Y(n_450) );
AOI31xp33_ASAP7_75t_L g451 ( .A1(n_380), .A2(n_180), .A3(n_142), .B(n_146), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_387), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_384), .A2(n_142), .B(n_146), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_385), .B(n_406), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
AOI221x1_ASAP7_75t_L g456 ( .A1(n_399), .A2(n_343), .B1(n_334), .B2(n_371), .C(n_375), .Y(n_456) );
OAI21xp5_ASAP7_75t_SL g457 ( .A1(n_399), .A2(n_377), .B(n_376), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_362), .Y(n_458) );
XOR2xp5_ASAP7_75t_SL g459 ( .A(n_398), .B(n_319), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_374), .Y(n_460) );
UNKNOWN g461 ( );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_364), .B(n_343), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_368), .B(n_369), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g464 ( .A1(n_462), .A2(n_436), .B(n_431), .C(n_423), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_459), .B(n_410), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_411), .B(n_424), .Y(n_466) );
NOR2x1p5_ASAP7_75t_L g467 ( .A(n_438), .B(n_449), .Y(n_467) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_443), .A2(n_462), .B1(n_420), .B2(n_435), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_456), .A2(n_457), .B(n_448), .Y(n_470) );
NAND2x1_ASAP7_75t_SL g471 ( .A(n_414), .B(n_425), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_408), .B(n_458), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g473 ( .A1(n_422), .A2(n_435), .B1(n_415), .B2(n_417), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_415), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_429), .B(n_455), .C(n_444), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_470), .B(n_444), .C(n_412), .Y(n_479) );
AOI322xp5_ASAP7_75t_L g480 ( .A1(n_465), .A2(n_440), .A3(n_433), .B1(n_463), .B2(n_439), .C1(n_418), .C2(n_413), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_472), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_464), .B(n_419), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_473), .A2(n_409), .B1(n_440), .B2(n_416), .C(n_452), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_470), .A2(n_432), .B1(n_446), .B2(n_439), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g485 ( .A1(n_477), .A2(n_407), .B(n_441), .C(n_445), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g486 ( .A1(n_471), .A2(n_421), .B(n_450), .C(n_414), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_476), .A2(n_430), .B1(n_421), .B2(n_437), .C(n_425), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_484), .A2(n_467), .B1(n_468), .B2(n_475), .Y(n_488) );
OAI211xp5_ASAP7_75t_L g489 ( .A1(n_479), .A2(n_483), .B(n_480), .C(n_485), .Y(n_489) );
AND4x1_ASAP7_75t_L g490 ( .A(n_487), .B(n_461), .C(n_466), .D(n_453), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_481), .B(n_474), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_482), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_490), .B(n_442), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_489), .B(n_486), .C(n_447), .D(n_454), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_491), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_494), .A2(n_488), .B1(n_492), .B2(n_469), .Y(n_496) );
AND3x4_ASAP7_75t_L g497 ( .A(n_493), .B(n_460), .C(n_432), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g498 ( .A(n_497), .B(n_495), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_498), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_499), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_500), .A2(n_496), .B1(n_451), .B2(n_478), .C(n_472), .Y(n_501) );
endmodule