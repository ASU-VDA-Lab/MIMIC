module real_aes_15899_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_876, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_876;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_769;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_0), .Y(n_597) );
AND2x4_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g143 ( .A(n_2), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_3), .A2(n_5), .B1(n_261), .B2(n_262), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_4), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_6), .A2(n_23), .B1(n_162), .B2(n_174), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_7), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_8), .A2(n_53), .B1(n_194), .B2(n_195), .Y(n_193) );
BUFx3_ASAP7_75t_L g554 ( .A(n_9), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_10), .A2(n_16), .B1(n_171), .B2(n_211), .Y(n_226) );
INVx1_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_12), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_13), .B(n_218), .Y(n_539) );
OR2x2_ASAP7_75t_L g110 ( .A(n_14), .B(n_32), .Y(n_110) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_15), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_17), .A2(n_85), .B1(n_521), .B2(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_17), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_18), .B(n_201), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_19), .B(n_239), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_20), .A2(n_87), .B1(n_174), .B2(n_201), .Y(n_603) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_21), .A2(n_49), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_22), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_24), .B(n_162), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_25), .B(n_169), .Y(n_285) );
INVx4_ASAP7_75t_R g247 ( .A(n_26), .Y(n_247) );
AO32x2_ASAP7_75t_L g600 ( .A1(n_27), .A2(n_180), .A3(n_181), .B1(n_601), .B2(n_604), .Y(n_600) );
AO32x1_ASAP7_75t_L g637 ( .A1(n_27), .A2(n_180), .A3(n_181), .B1(n_601), .B2(n_604), .Y(n_637) );
INVx1_ASAP7_75t_L g266 ( .A(n_28), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_29), .B(n_162), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_30), .A2(n_171), .B(n_172), .C(n_175), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_31), .A2(n_46), .B1(n_171), .B2(n_229), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_33), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_34), .A2(n_52), .B1(n_162), .B2(n_248), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_35), .A2(n_92), .B1(n_174), .B2(n_229), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_36), .B(n_541), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_37), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_37), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_38), .B(n_576), .Y(n_626) );
INVx1_ASAP7_75t_L g288 ( .A(n_39), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_40), .B(n_171), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_41), .A2(n_69), .B1(n_229), .B2(n_609), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_42), .Y(n_212) );
INVx2_ASAP7_75t_L g132 ( .A(n_43), .Y(n_132) );
BUFx3_ASAP7_75t_L g109 ( .A(n_44), .Y(n_109) );
INVx1_ASAP7_75t_L g125 ( .A(n_44), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_45), .B(n_628), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_47), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_48), .A2(n_86), .B1(n_171), .B2(n_229), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_50), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_51), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_54), .A2(n_79), .B1(n_203), .B2(n_576), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_55), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_56), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_56), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_57), .A2(n_83), .B1(n_174), .B2(n_201), .Y(n_550) );
INVx1_ASAP7_75t_L g157 ( .A(n_58), .Y(n_157) );
AND2x4_ASAP7_75t_L g177 ( .A(n_59), .B(n_178), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_60), .A2(n_91), .B1(n_229), .B2(n_259), .Y(n_258) );
AO22x1_ASAP7_75t_L g199 ( .A1(n_61), .A2(n_74), .B1(n_200), .B2(n_202), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_62), .B(n_174), .Y(n_538) );
INVx1_ASAP7_75t_L g178 ( .A(n_63), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_64), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_65), .B(n_180), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_66), .A2(n_191), .B(n_194), .C(n_596), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_67), .B(n_174), .C(n_543), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_68), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_70), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_71), .B(n_194), .Y(n_219) );
AND2x2_ASAP7_75t_L g598 ( .A(n_72), .B(n_252), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_73), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_75), .B(n_162), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_76), .A2(n_97), .B1(n_201), .B2(n_203), .Y(n_578) );
INVx2_ASAP7_75t_L g169 ( .A(n_77), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_78), .B(n_214), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_80), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_81), .B(n_180), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_82), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_84), .B(n_155), .Y(n_197) );
INVx1_ASAP7_75t_L g521 ( .A(n_85), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_88), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_89), .A2(n_102), .B1(n_229), .B2(n_248), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_90), .B(n_576), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_93), .B(n_180), .Y(n_208) );
INVx1_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_94), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_95), .B(n_239), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_96), .A2(n_194), .B(n_231), .C(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g251 ( .A(n_98), .B(n_252), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g136 ( .A(n_99), .Y(n_136) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_100), .B(n_218), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_101), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_116), .B(n_872), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx6f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_106), .Y(n_874) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g871 ( .A(n_108), .B(n_860), .Y(n_871) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g515 ( .A(n_109), .Y(n_515) );
INVx1_ASAP7_75t_L g126 ( .A(n_110), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
AND3x2_ASAP7_75t_L g138 ( .A(n_112), .B(n_126), .C(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g860 ( .A(n_113), .Y(n_860) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_127), .Y(n_116) );
INVx1_ASAP7_75t_L g134 ( .A(n_117), .Y(n_134) );
NOR2xp67_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx8_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_125), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_126), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_509), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g513 ( .A(n_132), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_132), .B(n_870), .Y(n_869) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .C(n_505), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .C(n_140), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_136), .B(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_137), .Y(n_507) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g508 ( .A(n_140), .Y(n_508) );
XNOR2x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_147), .Y(n_140) );
AOI22x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_143), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_146), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_147), .A2(n_524), .B1(n_859), .B2(n_861), .Y(n_523) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_405), .Y(n_147) );
NAND3xp33_ASAP7_75t_SL g148 ( .A(n_149), .B(n_307), .C(n_367), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_182), .B1(n_294), .B2(n_300), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g364 ( .A(n_151), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_151), .B(n_281), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_151), .B(n_327), .Y(n_475) );
AND2x2_ASAP7_75t_L g481 ( .A(n_151), .B(n_306), .Y(n_481) );
INVxp67_ASAP7_75t_L g486 ( .A(n_151), .Y(n_486) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g298 ( .A(n_152), .Y(n_298) );
AOI21x1_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_158), .B(n_179), .Y(n_152) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_153), .A2(n_257), .A3(n_263), .B(n_265), .Y(n_256) );
BUFx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_154), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g252 ( .A(n_154), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_154), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_154), .B(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_154), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI21xp33_ASAP7_75t_L g205 ( .A1(n_155), .A2(n_176), .B(n_197), .Y(n_205) );
INVx2_ASAP7_75t_L g232 ( .A(n_155), .Y(n_232) );
INVx2_ASAP7_75t_L g240 ( .A(n_155), .Y(n_240) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_170), .B(n_176), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_164), .B(n_167), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_162), .A2(n_248), .B1(n_592), .B2(n_593), .Y(n_591) );
INVx2_ASAP7_75t_L g609 ( .A(n_162), .Y(n_609) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g165 ( .A(n_163), .Y(n_165) );
INVx3_ASAP7_75t_L g171 ( .A(n_163), .Y(n_171) );
INVx2_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
INVx1_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
INVx1_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_163), .Y(n_218) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
INVx1_ASAP7_75t_L g248 ( .A(n_163), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx2_ASAP7_75t_L g262 ( .A(n_165), .Y(n_262) );
O2A1O1Ixp5_ASAP7_75t_L g558 ( .A1(n_167), .A2(n_262), .B(n_559), .C(n_560), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_167), .A2(n_175), .B1(n_602), .B2(n_603), .Y(n_601) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_168), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g543 ( .A(n_168), .Y(n_543) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx8_ASAP7_75t_L g175 ( .A(n_169), .Y(n_175) );
INVx2_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
INVx1_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
INVx4_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_SL g576 ( .A(n_174), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_175), .B(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_175), .A2(n_217), .B(n_219), .Y(n_216) );
INVx6_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_175), .A2(n_189), .B(n_199), .C(n_205), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_175), .A2(n_538), .B(n_539), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_175), .A2(n_227), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_176), .A2(n_590), .B(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx10_ASAP7_75t_L g222 ( .A(n_177), .Y(n_222) );
BUFx10_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
INVx1_ASAP7_75t_L g264 ( .A(n_177), .Y(n_264) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_177), .A2(n_573), .A3(n_607), .B(n_611), .Y(n_606) );
NOR2x1_ASAP7_75t_L g220 ( .A(n_180), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g335 ( .A(n_180), .Y(n_335) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g292 ( .A(n_181), .B(n_222), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_181), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g556 ( .A(n_181), .Y(n_556) );
BUFx3_ASAP7_75t_L g573 ( .A(n_181), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_181), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g620 ( .A(n_181), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_253), .B(n_267), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_223), .Y(n_184) );
INVx1_ASAP7_75t_L g402 ( .A(n_185), .Y(n_402) );
AND2x2_ASAP7_75t_L g431 ( .A(n_185), .B(n_393), .Y(n_431) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_206), .Y(n_185) );
AND2x2_ASAP7_75t_L g324 ( .A(n_186), .B(n_237), .Y(n_324) );
INVx1_ASAP7_75t_L g380 ( .A(n_186), .Y(n_380) );
AND2x2_ASAP7_75t_L g430 ( .A(n_186), .B(n_236), .Y(n_430) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g304 ( .A(n_187), .B(n_236), .Y(n_304) );
AND2x4_ASAP7_75t_L g449 ( .A(n_187), .B(n_237), .Y(n_449) );
AOI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_198), .B(n_204), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_193), .B(n_197), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_190), .A2(n_290), .B(n_291), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_190), .A2(n_227), .B1(n_333), .B2(n_334), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_190), .A2(n_227), .B1(n_608), .B2(n_610), .Y(n_607) );
AOI21x1_ASAP7_75t_L g622 ( .A1(n_190), .A2(n_623), .B(n_624), .Y(n_622) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g215 ( .A(n_192), .Y(n_215) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_196), .B(n_244), .Y(n_243) );
INVxp67_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g628 ( .A(n_201), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g284 ( .A1(n_202), .A2(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_203), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g374 ( .A(n_206), .Y(n_374) );
AND2x2_ASAP7_75t_L g443 ( .A(n_206), .B(n_237), .Y(n_443) );
AND2x2_ASAP7_75t_L g450 ( .A(n_206), .B(n_275), .Y(n_450) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
BUFx3_ASAP7_75t_L g306 ( .A(n_207), .Y(n_306) );
AND2x2_ASAP7_75t_L g317 ( .A(n_207), .B(n_303), .Y(n_317) );
AND2x2_ASAP7_75t_L g381 ( .A(n_207), .B(n_224), .Y(n_381) );
AND2x2_ASAP7_75t_L g386 ( .A(n_207), .B(n_237), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_216), .B(n_220), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .C(n_214), .Y(n_210) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_215), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_218), .A2(n_247), .B1(n_248), .B2(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AO31x2_ASAP7_75t_L g331 ( .A1(n_222), .A2(n_332), .A3(n_335), .B(n_336), .Y(n_331) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_222), .A2(n_537), .B(n_540), .Y(n_536) );
AOI31xp67_ASAP7_75t_L g548 ( .A1(n_222), .A2(n_335), .A3(n_549), .B(n_552), .Y(n_548) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_222), .A2(n_558), .B(n_561), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_223), .B(n_392), .Y(n_494) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_236), .Y(n_223) );
INVx2_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
OR2x2_ASAP7_75t_L g278 ( .A(n_224), .B(n_237), .Y(n_278) );
INVx2_ASAP7_75t_L g303 ( .A(n_224), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_224), .B(n_273), .Y(n_319) );
AND2x2_ASAP7_75t_L g393 ( .A(n_224), .B(n_237), .Y(n_393) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_232), .A3(n_233), .B(n_234), .Y(n_224) );
OAI22x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B1(n_228), .B2(n_230), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_230), .B1(n_258), .B2(n_260), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_227), .A2(n_575), .B1(n_577), .B2(n_578), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_227), .A2(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_229), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g541 ( .A(n_229), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_230), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_SL g577 ( .A(n_231), .Y(n_577) );
INVx1_ASAP7_75t_L g594 ( .A(n_231), .Y(n_594) );
INVx2_ASAP7_75t_L g535 ( .A(n_232), .Y(n_535) );
INVx2_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_241), .B(n_251), .Y(n_237) );
AOI21x1_ASAP7_75t_L g588 ( .A1(n_238), .A2(n_589), .B(n_598), .Y(n_588) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B(n_250), .Y(n_241) );
INVx1_ASAP7_75t_L g563 ( .A(n_248), .Y(n_563) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_254), .B(n_356), .Y(n_502) );
BUFx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g293 ( .A(n_256), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_256), .B(n_281), .Y(n_299) );
INVx1_ASAP7_75t_L g348 ( .A(n_256), .Y(n_348) );
OR2x2_ASAP7_75t_L g353 ( .A(n_256), .B(n_331), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_256), .B(n_331), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_256), .B(n_330), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_256), .B(n_298), .Y(n_438) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_263), .A2(n_573), .A3(n_574), .B(n_579), .Y(n_572) );
INVx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_SL g604 ( .A(n_264), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_276), .B(n_279), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
OR2x2_ASAP7_75t_L g277 ( .A(n_270), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g429 ( .A(n_270), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g459 ( .A(n_270), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_271), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g427 ( .A(n_271), .Y(n_427) );
OR2x2_ASAP7_75t_L g340 ( .A(n_272), .B(n_341), .Y(n_340) );
INVxp33_ASAP7_75t_L g458 ( .A(n_272), .Y(n_458) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx2_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI221xp5_ASAP7_75t_SL g424 ( .A1(n_277), .A2(n_349), .B1(n_354), .B2(n_425), .C(n_428), .Y(n_424) );
OR2x2_ASAP7_75t_L g411 ( .A(n_278), .B(n_362), .Y(n_411) );
INVx2_ASAP7_75t_L g460 ( .A(n_278), .Y(n_460) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g360 ( .A(n_280), .Y(n_360) );
OR2x2_ASAP7_75t_L g363 ( .A(n_280), .B(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_280), .Y(n_404) );
OR2x2_ASAP7_75t_L g417 ( .A(n_280), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_293), .Y(n_280) );
NAND2x1p5_ASAP7_75t_SL g312 ( .A(n_281), .B(n_297), .Y(n_312) );
INVx3_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_281), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_281), .Y(n_351) );
AND2x2_ASAP7_75t_L g432 ( .A(n_281), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g439 ( .A(n_281), .B(n_346), .Y(n_439) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_289), .B(n_292), .Y(n_283) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_299), .Y(n_294) );
AND2x2_ASAP7_75t_L g491 ( .A(n_295), .B(n_350), .Y(n_491) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g395 ( .A(n_297), .B(n_365), .Y(n_395) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g329 ( .A(n_298), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g356 ( .A(n_298), .B(n_331), .Y(n_356) );
AND2x4_ASAP7_75t_L g453 ( .A(n_299), .B(n_423), .Y(n_453) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g372 ( .A(n_304), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_305), .B(n_393), .Y(n_477) );
AND2x2_ASAP7_75t_L g484 ( .A(n_305), .B(n_444), .Y(n_484) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g409 ( .A(n_306), .Y(n_409) );
AOI321xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_321), .A3(n_338), .B1(n_339), .B2(n_342), .C(n_357), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_309), .B(n_318), .Y(n_308) );
AOI21xp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_314), .B(n_316), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI21xp33_ASAP7_75t_L g321 ( .A1(n_311), .A2(n_322), .B(n_325), .Y(n_321) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OR2x2_ASAP7_75t_L g421 ( .A(n_312), .B(n_353), .Y(n_421) );
INVx1_ASAP7_75t_L g413 ( .A(n_313), .Y(n_413) );
INVx2_ASAP7_75t_L g398 ( .A(n_314), .Y(n_398) );
OAI32xp33_ASAP7_75t_L g501 ( .A1(n_314), .A2(n_463), .A3(n_474), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g416 ( .A(n_315), .Y(n_416) );
INVx1_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_SL g454 ( .A(n_317), .B(n_361), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_318), .B(n_322), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_318), .A2(n_395), .B1(n_456), .B2(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g444 ( .A(n_319), .Y(n_444) );
INVx1_ASAP7_75t_L g341 ( .A(n_320), .Y(n_341) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g426 ( .A(n_324), .Y(n_426) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_325), .B(n_343), .C(n_349), .D(n_354), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVxp67_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
AND2x2_ASAP7_75t_L g447 ( .A(n_326), .B(n_356), .Y(n_447) );
OR2x2_ASAP7_75t_L g456 ( .A(n_326), .B(n_329), .Y(n_456) );
AND2x2_ASAP7_75t_L g480 ( .A(n_326), .B(n_352), .Y(n_480) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g394 ( .A(n_327), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g401 ( .A(n_327), .B(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g465 ( .A(n_328), .Y(n_465) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g373 ( .A(n_329), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g423 ( .A(n_329), .Y(n_423) );
INVx1_ASAP7_75t_L g365 ( .A(n_330), .Y(n_365) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g346 ( .A(n_331), .Y(n_346) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x4_ASAP7_75t_L g359 ( .A(n_345), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_347), .Y(n_464) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g418 ( .A(n_356), .Y(n_418) );
AND2x2_ASAP7_75t_L g461 ( .A(n_356), .B(n_401), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B(n_363), .C(n_366), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g472 ( .A(n_361), .B(n_450), .Y(n_472) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g376 ( .A(n_364), .Y(n_376) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_382), .C(n_396), .Y(n_367) );
OAI21xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_371), .A2(n_479), .B(n_482), .Y(n_478) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g392 ( .A(n_374), .Y(n_392) );
AND2x2_ASAP7_75t_L g452 ( .A(n_374), .B(n_449), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g471 ( .A(n_379), .Y(n_471) );
AND2x2_ASAP7_75t_L g497 ( .A(n_379), .B(n_460), .Y(n_497) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g385 ( .A(n_380), .Y(n_385) );
INVx2_ASAP7_75t_L g436 ( .A(n_381), .Y(n_436) );
NAND2x1_ASAP7_75t_L g470 ( .A(n_381), .B(n_471), .Y(n_470) );
AOI33xp33_ASAP7_75t_L g488 ( .A1(n_381), .A2(n_401), .A3(n_439), .B1(n_449), .B2(n_481), .B3(n_876), .Y(n_488) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_387), .B1(n_390), .B2(n_394), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g415 ( .A(n_386), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_387), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g500 ( .A(n_389), .B(n_434), .Y(n_500) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OAI22xp33_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_399), .B1(n_402), .B2(n_403), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_400), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_400), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_401), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g487 ( .A(n_401), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_466), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_424), .C(n_445), .D(n_462), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_412), .B1(n_414), .B2(n_417), .C(n_419), .Y(n_407) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_408), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g495 ( .A(n_411), .Y(n_495) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_415), .A2(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B(n_432), .C(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g474 ( .A(n_434), .B(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_SL g498 ( .A(n_434), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B1(n_440), .B2(n_442), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_451), .C(n_457), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_449), .A2(n_497), .B1(n_498), .B2(n_499), .C(n_501), .Y(n_496) );
INVx3_ASAP7_75t_L g504 ( .A(n_449), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_451) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_461), .Y(n_457) );
INVx1_ASAP7_75t_L g463 ( .A(n_460), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_489), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B(n_473), .C(n_476), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_472), .B(n_493), .C(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B(n_496), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_516), .B(n_865), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx6_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x6_ASAP7_75t_SL g512 ( .A(n_513), .B(n_514), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_769), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_526), .B(n_674), .C(n_701), .D(n_737), .Y(n_525) );
AOI221x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_585), .B1(n_613), .B2(n_649), .C(n_653), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_566), .C(n_583), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_546), .Y(n_530) );
INVx2_ASAP7_75t_L g614 ( .A(n_531), .Y(n_614) );
AND2x2_ASAP7_75t_L g787 ( .A(n_531), .B(n_731), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_531), .B(n_584), .Y(n_796) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g802 ( .A(n_532), .Y(n_802) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g647 ( .A(n_533), .Y(n_647) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g730 ( .A(n_534), .B(n_582), .Y(n_730) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_545), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_535), .A2(n_536), .B(n_545), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_544), .Y(n_540) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_546), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_546), .B(n_758), .Y(n_757) );
INVxp67_ASAP7_75t_L g800 ( .A(n_546), .Y(n_800) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_555), .Y(n_546) );
AND2x2_ASAP7_75t_L g584 ( .A(n_547), .B(n_572), .Y(n_584) );
INVx2_ASAP7_75t_L g656 ( .A(n_547), .Y(n_656) );
AND2x2_ASAP7_75t_L g721 ( .A(n_547), .B(n_659), .Y(n_721) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g582 ( .A(n_548), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g648 ( .A(n_555), .Y(n_648) );
AND2x2_ASAP7_75t_L g658 ( .A(n_555), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g720 ( .A(n_555), .B(n_572), .Y(n_720) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_565), .Y(n_555) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_556), .A2(n_557), .B(n_565), .Y(n_569) );
INVx1_ASAP7_75t_L g685 ( .A(n_566), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_568), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_568), .B(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_568), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_568), .B(n_755), .Y(n_762) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g731 ( .A(n_569), .B(n_706), .Y(n_731) );
OR2x2_ASAP7_75t_L g733 ( .A(n_569), .B(n_659), .Y(n_733) );
INVx1_ASAP7_75t_L g792 ( .A(n_569), .Y(n_792) );
BUFx2_ASAP7_75t_L g806 ( .A(n_569), .Y(n_806) );
OR2x2_ASAP7_75t_L g834 ( .A(n_569), .B(n_572), .Y(n_834) );
INVx1_ASAP7_75t_L g853 ( .A(n_570), .Y(n_853) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
OR2x2_ASAP7_75t_L g713 ( .A(n_571), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g732 ( .A(n_571), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_581), .Y(n_571) );
INVx2_ASAP7_75t_L g652 ( .A(n_572), .Y(n_652) );
AND2x2_ASAP7_75t_L g668 ( .A(n_572), .B(n_581), .Y(n_668) );
INVx1_ASAP7_75t_L g706 ( .A(n_572), .Y(n_706) );
INVx1_ASAP7_75t_L g749 ( .A(n_572), .Y(n_749) );
AND2x2_ASAP7_75t_L g791 ( .A(n_572), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g847 ( .A(n_583), .Y(n_847) );
AND2x4_ASAP7_75t_L g785 ( .A(n_584), .B(n_645), .Y(n_785) );
INVx2_ASAP7_75t_L g814 ( .A(n_584), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_584), .B(n_806), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_585), .B(n_804), .Y(n_803) );
AND2x4_ASAP7_75t_L g585 ( .A(n_586), .B(n_599), .Y(n_585) );
AND2x2_ASAP7_75t_L g725 ( .A(n_586), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g746 ( .A(n_586), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g617 ( .A(n_587), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g672 ( .A(n_587), .Y(n_672) );
AND2x2_ASAP7_75t_L g712 ( .A(n_587), .B(n_605), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_587), .B(n_696), .Y(n_753) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g665 ( .A(n_588), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_594), .Y(n_590) );
INVx3_ASAP7_75t_L g631 ( .A(n_599), .Y(n_631) );
AND2x2_ASAP7_75t_L g676 ( .A(n_599), .B(n_671), .Y(n_676) );
AND2x2_ASAP7_75t_L g831 ( .A(n_599), .B(n_635), .Y(n_831) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .Y(n_599) );
INVx1_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
AND2x2_ASAP7_75t_L g710 ( .A(n_600), .B(n_618), .Y(n_710) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_604), .A2(n_622), .B(n_625), .Y(n_621) );
AND2x4_ASAP7_75t_L g663 ( .A(n_605), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g636 ( .A(n_606), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g673 ( .A(n_606), .B(n_637), .Y(n_673) );
AND2x2_ASAP7_75t_L g683 ( .A(n_606), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_606), .B(n_618), .Y(n_735) );
AND2x2_ASAP7_75t_L g741 ( .A(n_606), .B(n_665), .Y(n_741) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_632), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_614), .A2(n_775), .B(n_779), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_614), .B(n_805), .Y(n_852) );
NAND2x1_ASAP7_75t_SL g615 ( .A(n_616), .B(n_630), .Y(n_615) );
INVx1_ASAP7_75t_L g858 ( .A(n_616), .Y(n_858) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g635 ( .A(n_618), .Y(n_635) );
INVx2_ASAP7_75t_L g640 ( .A(n_618), .Y(n_640) );
INVxp67_ASAP7_75t_L g661 ( .A(n_618), .Y(n_661) );
AND2x2_ASAP7_75t_L g681 ( .A(n_618), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g692 ( .A(n_618), .B(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g696 ( .A(n_618), .Y(n_696) );
INVx1_ASAP7_75t_L g714 ( .A(n_618), .Y(n_714) );
OR2x2_ASAP7_75t_L g747 ( .A(n_618), .B(n_682), .Y(n_747) );
INVx1_ASAP7_75t_L g818 ( .A(n_618), .Y(n_818) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B(n_629), .Y(n_619) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_638), .B(n_643), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_634), .A2(n_757), .B1(n_759), .B2(n_762), .Y(n_756) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_635), .B(n_683), .Y(n_717) );
BUFx2_ASAP7_75t_L g776 ( .A(n_635), .Y(n_776) );
INVx2_ASAP7_75t_L g726 ( .A(n_636), .Y(n_726) );
OR2x2_ASAP7_75t_L g810 ( .A(n_636), .B(n_640), .Y(n_810) );
INVx1_ASAP7_75t_L g642 ( .A(n_637), .Y(n_642) );
INVx1_ASAP7_75t_L g691 ( .A(n_637), .Y(n_691) );
NOR2x1p5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_640), .Y(n_761) );
OR2x2_ASAP7_75t_L g845 ( .A(n_640), .B(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g848 ( .A(n_640), .B(n_683), .Y(n_848) );
INVxp67_ASAP7_75t_SL g811 ( .A(n_641), .Y(n_811) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_645), .B(n_705), .Y(n_767) );
AND2x2_ASAP7_75t_L g857 ( .A(n_645), .B(n_655), .Y(n_857) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g766 ( .A(n_646), .B(n_655), .Y(n_766) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g723 ( .A(n_647), .B(n_656), .Y(n_723) );
AND2x2_ASAP7_75t_L g758 ( .A(n_647), .B(n_652), .Y(n_758) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g677 ( .A(n_650), .B(n_658), .Y(n_677) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g817 ( .A(n_652), .B(n_818), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_660), .B1(n_666), .B2(n_669), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g854 ( .A1(n_654), .A2(n_855), .B(n_856), .C(n_858), .Y(n_854) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g705 ( .A(n_656), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g773 ( .A(n_656), .Y(n_773) );
OR2x2_ASAP7_75t_L g820 ( .A(n_657), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g675 ( .A(n_661), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g778 ( .A(n_664), .Y(n_778) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g684 ( .A(n_665), .Y(n_684) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
INVx1_ASAP7_75t_L g765 ( .A(n_665), .Y(n_765) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g821 ( .A(n_668), .Y(n_821) );
AND2x2_ASAP7_75t_L g843 ( .A(n_668), .B(n_806), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_669), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g695 ( .A(n_673), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g751 ( .A(n_673), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g846 ( .A(n_673), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_678), .B2(n_685), .C(n_686), .Y(n_674) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx2_ASAP7_75t_L g768 ( .A(n_681), .Y(n_768) );
BUFx2_ASAP7_75t_L g788 ( .A(n_683), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_694), .B(n_697), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g830 ( .A(n_689), .B(n_752), .Y(n_830) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g736 ( .A(n_691), .Y(n_736) );
AND2x2_ASAP7_75t_L g826 ( .A(n_691), .B(n_696), .Y(n_826) );
INVx1_ASAP7_75t_L g709 ( .A(n_693), .Y(n_709) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_715), .C(n_727), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B1(n_711), .B2(n_713), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
BUFx2_ASAP7_75t_L g743 ( .A(n_710), .Y(n_743) );
AND2x2_ASAP7_75t_L g836 ( .A(n_710), .B(n_778), .Y(n_836) );
OAI21xp33_ASAP7_75t_L g839 ( .A1(n_711), .A2(n_840), .B(n_842), .Y(n_839) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B1(n_722), .B2(n_724), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_718), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AND2x4_ASAP7_75t_L g790 ( .A(n_723), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g777 ( .A(n_726), .B(n_778), .Y(n_777) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_726), .Y(n_793) );
AOI21xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_732), .B(n_734), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
AND2x2_ASAP7_75t_L g804 ( .A(n_729), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g841 ( .A(n_729), .B(n_806), .Y(n_841) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g755 ( .A(n_730), .Y(n_755) );
OR2x2_ASAP7_75t_L g833 ( .A(n_730), .B(n_834), .Y(n_833) );
OR2x2_ASAP7_75t_L g748 ( .A(n_733), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g780 ( .A(n_733), .Y(n_780) );
OR2x2_ASAP7_75t_L g813 ( .A(n_733), .B(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g784 ( .A(n_734), .Y(n_784) );
OR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_756), .C(n_763), .Y(n_737) );
OAI322xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_742), .A3(n_744), .B1(n_746), .B2(n_748), .C1(n_750), .C2(n_754), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_740), .A2(n_780), .B(n_816), .C(n_819), .Y(n_815) );
BUFx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g760 ( .A(n_741), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g797 ( .A(n_741), .Y(n_797) );
AND2x4_ASAP7_75t_L g825 ( .A(n_741), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI32xp33_ASAP7_75t_L g794 ( .A1(n_743), .A2(n_781), .A3(n_795), .B1(n_797), .B2(n_798), .Y(n_794) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g781 ( .A(n_747), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_749), .B(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_767), .C(n_768), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_770), .B(n_827), .Y(n_769) );
AOI211xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_774), .B(n_782), .C(n_807), .Y(n_770) );
INVxp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_SL g849 ( .A1(n_775), .A2(n_850), .B(n_851), .C(n_853), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
OAI31xp33_ASAP7_75t_L g829 ( .A1(n_777), .A2(n_830), .A3(n_831), .B(n_832), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g789 ( .A(n_781), .Y(n_789) );
NAND4xp25_ASAP7_75t_SL g782 ( .A(n_783), .B(n_786), .C(n_794), .D(n_803), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
AOI32xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .A3(n_789), .B1(n_790), .B2(n_793), .Y(n_786) );
INVx1_ASAP7_75t_L g838 ( .A(n_790), .Y(n_838) );
INVx1_ASAP7_75t_L g850 ( .A(n_793), .Y(n_850) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_815), .C(n_822), .Y(n_807) );
OAI21xp5_ASAP7_75t_SL g808 ( .A1(n_809), .A2(n_811), .B(n_812), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_816), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NOR4xp25_ASAP7_75t_L g827 ( .A(n_828), .B(n_839), .C(n_849), .D(n_854), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_835), .Y(n_828) );
OAI21xp33_ASAP7_75t_L g835 ( .A1(n_830), .A2(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_847), .B2(n_848), .Y(n_842) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_846), .Y(n_855) );
INVxp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx8_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_860), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx12f_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx5_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx10_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_SL g872 ( .A(n_873), .B(n_874), .Y(n_872) );
endmodule