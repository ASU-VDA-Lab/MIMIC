module fake_netlist_1_2348_n_704 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_704);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_704;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g79 ( .A(n_7), .Y(n_79) );
INVx3_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_12), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_14), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_72), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_44), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_55), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_45), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_30), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_78), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_70), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_28), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_49), .B(n_51), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_25), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_50), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_43), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_4), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_31), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_58), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_35), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_68), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_32), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_24), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_38), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_19), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_15), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_42), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_82), .B(n_1), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_112), .B(n_1), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_121), .B(n_2), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_118), .B(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_90), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_79), .B(n_3), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_92), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_122), .B(n_4), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
NAND2xp33_ASAP7_75t_SL g154 ( .A(n_86), .B(n_5), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_79), .B(n_5), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_97), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_97), .A2(n_29), .B(n_75), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_113), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_113), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_110), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_117), .Y(n_168) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_119), .A2(n_26), .B(n_71), .Y(n_169) );
INVx5_ASAP7_75t_L g170 ( .A(n_119), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_139), .B(n_90), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_133), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_139), .B(n_84), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_136), .B(n_120), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_141), .B(n_98), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_136), .B(n_96), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_136), .B(n_124), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_136), .B(n_124), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_128), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_134), .B(n_84), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_128), .B(n_122), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_146), .B(n_103), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_144), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_146), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_128), .B(n_108), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_128), .B(n_83), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_128), .B(n_83), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_146), .B(n_102), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_134), .B(n_109), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_127), .B(n_111), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_144), .Y(n_206) );
INVxp67_ASAP7_75t_SL g207 ( .A(n_127), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_129), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_135), .B(n_107), .Y(n_211) );
INVx5_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_157), .B(n_103), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_157), .B(n_120), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_135), .B(n_106), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_131), .B(n_116), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_129), .Y(n_219) );
OR2x2_ASAP7_75t_SL g220 ( .A(n_162), .B(n_125), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
AOI22xp5_ASAP7_75t_SL g225 ( .A1(n_133), .A2(n_123), .B1(n_91), .B2(n_126), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_131), .B(n_125), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_157), .B(n_115), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
INVx5_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_137), .B(n_114), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_131), .B(n_105), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_137), .B(n_101), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_132), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_226), .B(n_132), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_171), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_176), .B(n_132), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_173), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_180), .A2(n_156), .B1(n_143), .B2(n_148), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_173), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_233), .A2(n_154), .B1(n_158), .B2(n_156), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
AND3x1_ASAP7_75t_L g244 ( .A(n_217), .B(n_150), .C(n_154), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_226), .B(n_150), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_187), .B(n_153), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_174), .B(n_153), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_207), .B(n_155), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_175), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_201), .B(n_155), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_190), .A2(n_152), .B1(n_143), .B2(n_142), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_191), .B(n_158), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_226), .B(n_151), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_181), .B(n_152), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_226), .B1(n_191), .B2(n_217), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_190), .A2(n_164), .B1(n_140), .B2(n_142), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_179), .Y(n_261) );
BUFx2_ASAP7_75t_SL g262 ( .A(n_180), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_148), .B1(n_151), .B2(n_160), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_190), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_175), .Y(n_266) );
NAND3xp33_ASAP7_75t_SL g267 ( .A(n_214), .B(n_100), .C(n_104), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_209), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_202), .B(n_160), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_221), .B(n_140), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_231), .B(n_205), .Y(n_273) );
NOR2xp33_ASAP7_75t_R g274 ( .A(n_180), .B(n_188), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_180), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_195), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_231), .B(n_161), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_173), .B(n_163), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_180), .A2(n_164), .B1(n_161), .B2(n_167), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_198), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_183), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_215), .B(n_167), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_183), .A2(n_163), .B1(n_129), .B2(n_130), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_215), .B(n_163), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_209), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_215), .B(n_163), .Y(n_289) );
AO22x1_ASAP7_75t_L g290 ( .A1(n_215), .A2(n_163), .B1(n_130), .B2(n_149), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_198), .Y(n_291) );
AND2x6_ASAP7_75t_SL g292 ( .A(n_225), .B(n_6), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_221), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_221), .A2(n_168), .B1(n_130), .B2(n_149), .Y(n_294) );
BUFx8_ASAP7_75t_SL g295 ( .A(n_225), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_189), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_178), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_223), .A2(n_166), .B1(n_149), .B2(n_145), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_189), .B(n_145), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_178), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_296), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_257), .B(n_234), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_257), .B(n_183), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_245), .A2(n_223), .B1(n_183), .B2(n_184), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_245), .B(n_184), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_243), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_234), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_245), .A2(n_223), .B1(n_184), .B2(n_203), .Y(n_313) );
OAI321xp33_ASAP7_75t_L g314 ( .A1(n_251), .A2(n_232), .A3(n_230), .B1(n_216), .B2(n_211), .C(n_147), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_280), .A2(n_182), .B(n_184), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_264), .B(n_223), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_261), .B(n_203), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_237), .B(n_203), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_271), .Y(n_321) );
CKINVDCx8_ASAP7_75t_R g322 ( .A(n_262), .Y(n_322) );
AND2x6_ASAP7_75t_L g323 ( .A(n_265), .B(n_188), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_243), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
BUFx12f_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_271), .Y(n_327) );
BUFx6f_ASAP7_75t_SL g328 ( .A(n_268), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_256), .B(n_203), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_249), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_243), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_276), .B(n_227), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_236), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_243), .B(n_200), .Y(n_336) );
BUFx8_ASAP7_75t_SL g337 ( .A(n_295), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_253), .Y(n_338) );
AND2x2_ASAP7_75t_SL g339 ( .A(n_253), .B(n_227), .Y(n_339) );
NOR3xp33_ASAP7_75t_L g340 ( .A(n_273), .B(n_204), .C(n_188), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_256), .B(n_200), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_275), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_248), .B(n_200), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_275), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_270), .B(n_189), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_283), .A2(n_227), .B1(n_196), .B2(n_194), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_288), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_263), .B(n_200), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_236), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_240), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_295), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_339), .A2(n_266), .B1(n_259), .B2(n_283), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_335), .Y(n_355) );
OR2x6_ASAP7_75t_SL g356 ( .A(n_352), .B(n_260), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_345), .B(n_278), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_339), .A2(n_293), .B1(n_267), .B2(n_242), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_326), .A2(n_270), .B1(n_247), .B2(n_250), .Y(n_361) );
BUFx8_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_350), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_350), .Y(n_364) );
CKINVDCx6p67_ASAP7_75t_R g365 ( .A(n_328), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_351), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_302), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_311), .A2(n_293), .B1(n_287), .B2(n_258), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_SL g370 ( .A1(n_327), .A2(n_279), .B(n_272), .C(n_255), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_321), .B(n_274), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_348), .A2(n_227), .B1(n_284), .B2(n_239), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_309), .A2(n_162), .B(n_169), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_312), .B(n_287), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_326), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_331), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_321), .A2(n_281), .B1(n_194), .B2(n_196), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_345), .B(n_240), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_321), .A2(n_194), .B1(n_196), .B2(n_291), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_316), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_312), .B(n_287), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_318), .A2(n_246), .B(n_286), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_301), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_303), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_244), .B1(n_319), .B2(n_334), .C(n_329), .Y(n_386) );
NAND4xp25_ASAP7_75t_L g387 ( .A(n_376), .B(n_340), .C(n_189), .D(n_313), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_367), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_317), .B1(n_312), .B2(n_320), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_378), .B(n_303), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_358), .B(n_306), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_383), .A2(n_325), .B1(n_341), .B2(n_314), .C(n_343), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_359), .A2(n_317), .B1(n_328), .B2(n_309), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_370), .A2(n_327), .B(n_290), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_309), .B1(n_304), .B2(n_308), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_380), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_307), .B1(n_323), .B2(n_305), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_362), .A2(n_323), .B1(n_315), .B2(n_347), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_362), .A2(n_352), .B1(n_323), .B2(n_262), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_298), .B1(n_290), .B2(n_346), .C(n_289), .Y(n_400) );
CKINVDCx6p67_ASAP7_75t_R g401 ( .A(n_365), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_362), .A2(n_323), .B1(n_347), .B2(n_338), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_381), .A2(n_285), .B(n_165), .C(n_145), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_255), .B(n_277), .C(n_291), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_381), .B(n_338), .Y(n_405) );
BUFx10_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_369), .A2(n_165), .B(n_159), .C(n_149), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_159), .B(n_165), .C(n_166), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_362), .A2(n_323), .B1(n_338), .B2(n_336), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_357), .A2(n_159), .B(n_166), .C(n_280), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_372), .A2(n_322), .B1(n_277), .B2(n_269), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_385), .A2(n_323), .B1(n_336), .B2(n_342), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_405), .B(n_380), .Y(n_414) );
OAI33xp33_ASAP7_75t_L g415 ( .A1(n_387), .A2(n_379), .A3(n_166), .B1(n_372), .B2(n_377), .B3(n_360), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_388), .B(n_380), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_391), .B(n_357), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_386), .A2(n_385), .B1(n_365), .B2(n_360), .Y(n_419) );
OAI21x1_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_373), .B(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_409), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_409), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_405), .B(n_363), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_389), .A2(n_392), .B1(n_393), .B2(n_390), .Y(n_424) );
AOI33xp33_ASAP7_75t_L g425 ( .A1(n_395), .A2(n_356), .A3(n_294), .B1(n_199), .B2(n_224), .B3(n_218), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_390), .B(n_375), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_406), .A2(n_375), .B1(n_405), .B2(n_412), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_396), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_396), .B(n_363), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_406), .B(n_354), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_356), .B1(n_379), .B2(n_355), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_410), .B(n_354), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_399), .A2(n_382), .B(n_371), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_354), .Y(n_436) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_404), .A2(n_373), .B(n_355), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_404), .B(n_355), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_413), .B(n_364), .Y(n_439) );
AOI322xp5_ASAP7_75t_L g440 ( .A1(n_398), .A2(n_337), .A3(n_7), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_402), .A2(n_382), .B(n_374), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_407), .A2(n_377), .B1(n_374), .B2(n_147), .C(n_364), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_411), .A2(n_364), .B1(n_322), .B2(n_382), .Y(n_443) );
OAI211xp5_ASAP7_75t_SL g444 ( .A1(n_408), .A2(n_337), .B(n_224), .C(n_199), .Y(n_444) );
OAI21x1_ASAP7_75t_L g445 ( .A1(n_400), .A2(n_384), .B(n_169), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_403), .A2(n_162), .B(n_169), .C(n_147), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_401), .B(n_384), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_388), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_448), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_434), .B(n_384), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g453 ( .A(n_440), .B(n_374), .C(n_219), .D(n_10), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_415), .A2(n_219), .B1(n_170), .B2(n_11), .C1(n_12), .C2(n_13), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_421), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_448), .B(n_169), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_423), .Y(n_458) );
OAI31xp33_ASAP7_75t_L g459 ( .A1(n_433), .A2(n_336), .A3(n_252), .B(n_235), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_423), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_428), .A2(n_366), .B1(n_349), .B2(n_220), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_430), .B(n_169), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_162), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_427), .B(n_6), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_423), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_429), .Y(n_468) );
OAI33xp33_ASAP7_75t_L g469 ( .A1(n_418), .A2(n_218), .A3(n_228), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_424), .A2(n_162), .B1(n_170), .B2(n_349), .C(n_210), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_425), .B(n_208), .C(n_170), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_426), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_414), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_431), .B(n_9), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_419), .B(n_14), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_416), .B(n_208), .C(n_170), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_431), .B(n_366), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_438), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_414), .B(n_439), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
AND4x1_ASAP7_75t_L g483 ( .A(n_442), .B(n_16), .C(n_18), .D(n_19), .Y(n_483) );
OAI33xp33_ASAP7_75t_L g484 ( .A1(n_447), .A2(n_228), .A3(n_18), .B1(n_20), .B2(n_21), .B3(n_222), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_414), .B(n_366), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_437), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_434), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_432), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_429), .B(n_447), .C(n_441), .D(n_435), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_436), .B(n_366), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_434), .B(n_20), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_437), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_439), .B(n_366), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_420), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_445), .B(n_366), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_475), .B(n_445), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_451), .B(n_443), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_453), .A2(n_444), .B1(n_446), .B2(n_420), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_491), .B(n_21), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_481), .B(n_349), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_489), .B(n_22), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_490), .B(n_493), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_449), .B(n_349), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_458), .B(n_349), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_453), .B(n_210), .C(n_213), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_468), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_491), .B(n_213), .C(n_222), .D(n_192), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_452), .B(n_170), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_476), .B(n_220), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_455), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_458), .B(n_33), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_462), .B(n_37), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_462), .B(n_39), .Y(n_523) );
OAI21xp33_ASAP7_75t_SL g524 ( .A1(n_459), .A2(n_40), .B(n_47), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_492), .B(n_48), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_450), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_52), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_457), .B(n_170), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_466), .B(n_454), .C(n_494), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_492), .B(n_473), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_461), .B(n_170), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_474), .B(n_54), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_484), .B(n_197), .C(n_192), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_471), .A2(n_170), .B(n_177), .Y(n_536) );
AOI211xp5_ASAP7_75t_L g537 ( .A1(n_463), .A2(n_208), .B(n_186), .C(n_177), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_482), .Y(n_538) );
OR2x6_ASAP7_75t_L g539 ( .A(n_473), .B(n_342), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_475), .B(n_479), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_482), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_459), .B(n_206), .C(n_197), .D(n_193), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_478), .B(n_56), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g544 ( .A(n_480), .B(n_206), .C(n_193), .D(n_254), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_480), .B(n_59), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_483), .B(n_208), .C(n_186), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_485), .B(n_60), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g548 ( .A(n_479), .B(n_297), .C(n_300), .D(n_67), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_472), .B(n_62), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_489), .B(n_63), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_472), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_496), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_483), .B(n_208), .C(n_186), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_496), .Y(n_554) );
NAND4xp25_ASAP7_75t_SL g555 ( .A(n_471), .B(n_77), .C(n_332), .D(n_324), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_450), .B(n_186), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_535), .B(n_450), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_505), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_513), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_516), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_507), .B(n_450), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_540), .B(n_495), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_535), .B(n_495), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_510), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_503), .B(n_469), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_503), .A2(n_470), .B1(n_488), .B2(n_487), .C(n_486), .Y(n_570) );
XOR2xp5_ASAP7_75t_L g571 ( .A(n_554), .B(n_477), .Y(n_571) );
OAI33xp33_ASAP7_75t_L g572 ( .A1(n_529), .A2(n_497), .A3(n_488), .B1(n_486), .B2(n_487), .B3(n_477), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_556), .B(n_465), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_526), .B(n_552), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_512), .A2(n_498), .B1(n_464), .B2(n_465), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_519), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_498), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_521), .B(n_464), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_512), .B(n_497), .C(n_488), .D(n_456), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_526), .B(n_456), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_554), .B(n_186), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_509), .B(n_344), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_510), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_531), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_504), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_509), .B(n_212), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_501), .B(n_212), .Y(n_587) );
NAND2xp33_ASAP7_75t_R g588 ( .A(n_520), .B(n_300), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_526), .B(n_212), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_538), .B(n_212), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_499), .B(n_212), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_499), .B(n_212), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_511), .B(n_229), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_551), .B(n_229), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_506), .Y(n_597) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_524), .A2(n_229), .B(n_344), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_518), .B(n_229), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_514), .B(n_297), .C(n_238), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_506), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_506), .Y(n_602) );
AOI31xp33_ASAP7_75t_L g603 ( .A1(n_546), .A2(n_238), .A3(n_241), .B(n_344), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_344), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_SL g606 ( .A1(n_553), .A2(n_241), .B(n_344), .C(n_342), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_557), .B(n_229), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_539), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_557), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_569), .B(n_560), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_559), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_577), .B(n_550), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_574), .B(n_550), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_569), .A2(n_518), .B1(n_548), .B2(n_502), .C(n_527), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_606), .A2(n_555), .B(n_537), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_562), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_608), .A2(n_544), .B1(n_533), .B2(n_536), .C(n_545), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_568), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_566), .B(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_608), .B(n_525), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_576), .B(n_547), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_603), .B(n_549), .Y(n_623) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_574), .B(n_539), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_585), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_573), .B(n_539), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_596), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_596), .B(n_523), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_571), .B(n_522), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_609), .B(n_532), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_584), .B(n_528), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_565), .B(n_515), .Y(n_634) );
NAND2x1_ASAP7_75t_L g635 ( .A(n_594), .B(n_534), .Y(n_635) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_564), .B(n_534), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_609), .B(n_542), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_578), .B(n_229), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_588), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_583), .B(n_342), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_583), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_591), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_592), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_563), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_301), .B(n_310), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_558), .Y(n_647) );
OA22x2_ASAP7_75t_L g648 ( .A1(n_575), .A2(n_301), .B1(n_310), .B2(n_324), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_579), .A2(n_301), .B1(n_310), .B2(n_324), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_570), .A2(n_310), .B1(n_324), .B2(n_332), .C(n_602), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_594), .B(n_310), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_581), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_580), .B(n_324), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_580), .B(n_332), .Y(n_654) );
XNOR2x1_ASAP7_75t_L g655 ( .A(n_607), .B(n_332), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_597), .B(n_332), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_607), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_601), .B(n_604), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_599), .A2(n_570), .B1(n_586), .B2(n_593), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_600), .B(n_587), .C(n_606), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_590), .Y(n_662) );
AO22x2_ASAP7_75t_L g663 ( .A1(n_572), .A2(n_600), .B1(n_605), .B2(n_589), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_595), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_572), .B(n_566), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_560), .B(n_513), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_559), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_610), .B(n_665), .C(n_614), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_610), .A2(n_636), .B1(n_663), .B2(n_627), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_663), .A2(n_636), .B(n_658), .Y(n_670) );
NOR2xp33_ASAP7_75t_R g671 ( .A(n_666), .B(n_631), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_640), .A2(n_617), .B(n_621), .C(n_623), .Y(n_672) );
OA22x2_ASAP7_75t_L g673 ( .A1(n_624), .A2(n_625), .B1(n_621), .B2(n_630), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_635), .A2(n_660), .B(n_661), .Y(n_674) );
AOI211x1_ASAP7_75t_SL g675 ( .A1(n_661), .A2(n_637), .B(n_615), .C(n_623), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g676 ( .A1(n_647), .A2(n_648), .B(n_612), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_659), .A2(n_664), .B1(n_629), .B2(n_630), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_657), .A2(n_612), .B1(n_620), .B2(n_648), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g679 ( .A(n_613), .B(n_662), .C(n_634), .D(n_654), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_613), .A2(n_657), .A3(n_667), .B1(n_611), .B2(n_619), .C1(n_616), .C2(n_639), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_655), .A2(n_632), .B1(n_652), .B2(n_628), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_670), .B(n_638), .C(n_650), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_668), .B(n_628), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_675), .B(n_646), .C(n_633), .D(n_653), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_677), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g686 ( .A1(n_674), .A2(n_649), .B(n_646), .C(n_622), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_669), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_672), .A2(n_642), .B1(n_644), .B2(n_643), .C(n_626), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_673), .A2(n_626), .B(n_645), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_685), .B(n_678), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_688), .B(n_676), .Y(n_691) );
NOR2x2_ASAP7_75t_L g692 ( .A(n_687), .B(n_679), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_684), .B(n_656), .C(n_641), .Y(n_693) );
NAND2x1_ASAP7_75t_L g694 ( .A(n_683), .B(n_681), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_693), .B(n_682), .Y(n_695) );
AND3x2_ASAP7_75t_L g696 ( .A(n_692), .B(n_686), .C(n_671), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_690), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_696), .B(n_694), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
XOR2xp5_ASAP7_75t_L g700 ( .A(n_699), .B(n_695), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_698), .A2(n_691), .B1(n_689), .B2(n_680), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
BUFx4_ASAP7_75t_R g703 ( .A(n_702), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_701), .B1(n_651), .B2(n_632), .C(n_618), .Y(n_704) );
endmodule