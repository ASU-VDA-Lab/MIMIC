module fake_jpeg_2280_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_1),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_2),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_50),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_63),
.B(n_68),
.C(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OR2x4_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_52),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_52),
.C(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_67),
.B1(n_51),
.B2(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_70),
.B1(n_57),
.B2(n_76),
.Y(n_96)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_60),
.B(n_68),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_67),
.B1(n_53),
.B2(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_56),
.B1(n_66),
.B2(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_87),
.B1(n_84),
.B2(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_54),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_110),
.B1(n_86),
.B2(n_92),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_54),
.B(n_55),
.C(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_95),
.B1(n_51),
.B2(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_115),
.B1(n_121),
.B2(n_122),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_65),
.B1(n_55),
.B2(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_124),
.B1(n_102),
.B2(n_9),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_12),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_62),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_5),
.B(n_7),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_11),
.B(n_12),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_7),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_24),
.C(n_47),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_30),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_26),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_144),
.B1(n_147),
.B2(n_152),
.C(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_8),
.Y(n_138)
);

OAI211xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_140),
.B(n_143),
.C(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_11),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_29),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_23),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_156),
.A2(n_122),
.B1(n_16),
.B2(n_17),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_164),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_34),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_167),
.B(n_173),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_14),
.B(n_18),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_147),
.B1(n_144),
.B2(n_136),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_19),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_22),
.B(n_31),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_142),
.C(n_145),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_183),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_163),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_36),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_38),
.C(n_41),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_43),
.C(n_44),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_188),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_169),
.B1(n_167),
.B2(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_175),
.C(n_181),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_177),
.B(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_195),
.B1(n_164),
.B2(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_165),
.B1(n_161),
.B2(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_196),
.A3(n_190),
.B1(n_198),
.B2(n_161),
.C1(n_165),
.C2(n_174),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_184),
.C(n_46),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_49),
.Y(n_204)
);


endmodule