module fake_jpeg_22099_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_16),
.B1(n_24),
.B2(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_61),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_39),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_37),
.B1(n_31),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_78),
.B1(n_81),
.B2(n_19),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_42),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_80),
.B1(n_32),
.B2(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_24),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_21),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_25),
.B1(n_19),
.B2(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_24),
.B1(n_37),
.B2(n_21),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_99),
.B1(n_102),
.B2(n_110),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_24),
.B1(n_36),
.B2(n_48),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_93),
.A2(n_62),
.B1(n_57),
.B2(n_72),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_104),
.B1(n_82),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_112),
.B1(n_85),
.B2(n_60),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_50),
.B1(n_47),
.B2(n_35),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_47),
.A3(n_44),
.B1(n_55),
.B2(n_40),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_108),
.B1(n_70),
.B2(n_72),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_22),
.B1(n_26),
.B2(n_32),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_35),
.B1(n_32),
.B2(n_22),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_40),
.A3(n_17),
.B1(n_27),
.B2(n_23),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_66),
.B1(n_26),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_29),
.B1(n_30),
.B2(n_25),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_83),
.Y(n_120)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_118),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_116),
.B(n_120),
.Y(n_154)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_99),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_127),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_131),
.B1(n_133),
.B2(n_138),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_141),
.B1(n_84),
.B2(n_89),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_140),
.Y(n_171)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_139),
.B1(n_113),
.B2(n_91),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_108),
.B(n_89),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_40),
.B(n_17),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_85),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_77),
.B1(n_65),
.B2(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_84),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_93),
.B(n_91),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_143),
.A2(n_152),
.B(n_173),
.Y(n_205)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_147),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_88),
.B1(n_112),
.B2(n_96),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_150),
.B1(n_133),
.B2(n_124),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_88),
.B1(n_96),
.B2(n_103),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_88),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_162),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_90),
.B1(n_105),
.B2(n_107),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_23),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_105),
.B1(n_30),
.B2(n_28),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_163),
.B(n_165),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_115),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_17),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_100),
.B(n_15),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_100),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_164),
.B(n_15),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_126),
.B(n_142),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_28),
.C(n_27),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_116),
.C(n_121),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_28),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_175),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_15),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_28),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_200),
.B1(n_203),
.B2(n_148),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_189),
.C(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_181),
.Y(n_217)
);

AO22x2_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_131),
.B1(n_23),
.B2(n_27),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_147),
.B1(n_169),
.B2(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_124),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_191),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_137),
.C(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_151),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_194),
.B(n_196),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_117),
.B1(n_15),
.B2(n_2),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_207),
.B(n_13),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_145),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_1),
.C(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_3),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_230),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_214),
.B1(n_215),
.B2(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_223),
.B1(n_231),
.B2(n_201),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_183),
.A2(n_171),
.B1(n_168),
.B2(n_143),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_150),
.B1(n_167),
.B2(n_162),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_175),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_14),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_13),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_227),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_4),
.C(n_6),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_229),
.C(n_206),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_12),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_11),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_195),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_179),
.B1(n_197),
.B2(n_182),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_185),
.C(n_177),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_192),
.C(n_205),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_205),
.C(n_179),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_179),
.C(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_247),
.Y(n_254)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_249),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

XNOR2x2_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_200),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_226),
.B(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_252),
.B(n_213),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_187),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_222),
.B(n_219),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_269),
.B(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_231),
.B1(n_204),
.B2(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_214),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_221),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_228),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_241),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_203),
.B(n_198),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_239),
.C(n_255),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_280),
.B1(n_281),
.B2(n_203),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_276),
.B(n_279),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_265),
.B1(n_259),
.B2(n_262),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_203),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_256),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_267),
.B1(n_260),
.B2(n_234),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_294),
.B1(n_275),
.B2(n_11),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_6),
.C(n_7),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_291),
.B(n_293),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_280),
.B(n_270),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_264),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_278),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_241),
.B1(n_11),
.B2(n_8),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_10),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_291),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_309),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_295),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_305),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_310),
.Y(n_316)
);

AOI321xp33_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_308),
.C(n_310),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_9),
.Y(n_319)
);


endmodule