module real_jpeg_29920_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_23),
.B1(n_26),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_0),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_0),
.A2(n_28),
.B1(n_32),
.B2(n_109),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_0),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_0),
.A2(n_59),
.B1(n_61),
.B2(n_109),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_1),
.B(n_27),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_32),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_32),
.B(n_209),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_168),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_1),
.A2(n_56),
.B(n_59),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_76),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_1),
.A2(n_97),
.B1(n_113),
.B2(n_257),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_49),
.B1(n_59),
.B2(n_61),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_67),
.Y(n_72)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_170),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_170),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_59),
.B1(n_61),
.B2(n_170),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_9),
.A2(n_28),
.B1(n_32),
.B2(n_135),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_135),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_9),
.A2(n_59),
.B1(n_61),
.B2(n_135),
.Y(n_249)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_25),
.B1(n_59),
.B2(n_61),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_23),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_38),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_38),
.B1(n_59),
.B2(n_61),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_118)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_15),
.A2(n_23),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_15),
.A2(n_28),
.B1(n_32),
.B2(n_47),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_15),
.A2(n_47),
.B1(n_59),
.B2(n_61),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_340),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_81),
.B(n_338),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_20),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_21),
.A2(n_45),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_22),
.A2(n_34),
.B(n_80),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_340)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_30),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_30),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_23),
.B(n_168),
.CON(n_167),
.SN(n_167)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_27),
.A2(n_34),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_28),
.A2(n_35),
.B1(n_167),
.B2(n_181),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_28),
.A2(n_54),
.A3(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_30),
.B(n_32),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_33),
.A2(n_46),
.B(n_50),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_34),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_40),
.B(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_73),
.C(n_78),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_41),
.A2(n_42),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.C(n_64),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_43),
.A2(n_44),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_45),
.A2(n_50),
.B1(n_108),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_45),
.A2(n_50),
.B1(n_134),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_51),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_51),
.A2(n_64),
.B1(n_306),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_62),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_52),
.A2(n_101),
.B(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_52),
.A2(n_62),
.B(n_117),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_52),
.A2(n_58),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_52),
.A2(n_141),
.B(n_217),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_52),
.A2(n_58),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_52),
.A2(n_58),
.B1(n_216),
.B2(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_55),
.B(n_207),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_55),
.A2(n_57),
.B(n_168),
.C(n_236),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_100),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_58),
.B(n_168),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_61),
.B(n_261),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_63),
.B(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_65),
.A2(n_75),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_70),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_66),
.A2(n_71),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_66),
.A2(n_71),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_66),
.A2(n_71),
.B1(n_164),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_66),
.A2(n_71),
.B1(n_192),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_76),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_75),
.A2(n_77),
.B(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_75),
.A2(n_131),
.B(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_78),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_331),
.B(n_337),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_301),
.A3(n_323),
.B1(n_329),
.B2(n_330),
.C(n_342),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_153),
.B(n_300),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_136),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_85),
.B(n_136),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_110),
.C(n_121),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_86),
.A2(n_87),
.B1(n_110),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_102),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_104),
.C(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_89),
.B(n_99),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_90),
.A2(n_183),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_91),
.A2(n_98),
.B(n_126),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_91),
.A2(n_96),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_95),
.A2(n_113),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_97),
.A2(n_113),
.B1(n_124),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_110),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_120),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_112),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_116),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_112),
.A2(n_147),
.B(n_150),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_113),
.A2(n_196),
.B1(n_249),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_121),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.C(n_132),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_122),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_127),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_130),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_151),
.B2(n_152),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_139),
.B(n_146),
.C(n_152),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B(n_145),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_142),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_144),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_145),
.B(n_303),
.C(n_313),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_145),
.A2(n_303),
.B1(n_304),
.B2(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_145),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_294),
.B(n_299),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_197),
.B(n_280),
.C(n_293),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_184),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_156),
.B(n_184),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_171),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_158),
.B(n_159),
.C(n_171),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_173),
.B(n_177),
.C(n_179),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_185),
.A2(n_186),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_195),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_279),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_272),
.B(n_278),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_227),
.B(n_271),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_218),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_201),
.B(n_218),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_211),
.C(n_214),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_202),
.A2(n_203),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_205),
.Y(n_225)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_225),
.C(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_265),
.B(n_270),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_245),
.B(n_264),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_230),
.B(n_237),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_253),
.B(n_263),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_251),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_262),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_291),
.B2(n_292),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.C(n_292),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_315),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_312),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_321),
.C(n_322),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_314),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_322),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);


endmodule