module fake_netlist_6_3081_n_1234 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1234);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1234;

wire n_992;
wire n_801;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;

INVxp67_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_24),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_69),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_93),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_44),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_49),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_5),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_48),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_22),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_78),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_15),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_148),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_79),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_143),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_140),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_56),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_8),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_18),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_47),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_102),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_106),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_213),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_222),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_185),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_186),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_216),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_191),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_195),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_212),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_215),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_217),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_221),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_240),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g273 ( 
.A(n_242),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_249),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_245),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_258),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_206),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_260),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_237),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_243),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_242),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_243),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_179),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_273),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_272),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_275),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_300),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_270),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_274),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_306),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_278),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_274),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_269),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_290),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_284),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_205),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_292),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_283),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_193),
.Y(n_369)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_193),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_315),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_368),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_271),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_220),
.Y(n_375)
);

BUFx12f_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_291),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_231),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_289),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_327),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_329),
.B(n_225),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_312),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_203),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_298),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_203),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_299),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_313),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_314),
.Y(n_399)
);

BUFx8_ASAP7_75t_SL g400 ( 
.A(n_346),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_320),
.B(n_276),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_276),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_312),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g405 ( 
.A(n_334),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

BUFx12f_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_365),
.B(n_310),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_292),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_308),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_282),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_308),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_364),
.B1(n_343),
.B2(n_340),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_317),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_386),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_402),
.A2(n_321),
.B1(n_367),
.B2(n_346),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_374),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_305),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_312),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_382),
.A2(n_340),
.B1(n_364),
.B2(n_343),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_376),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_317),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_334),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_398),
.A2(n_307),
.B(n_224),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_411),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_390),
.A2(n_37),
.B(n_35),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_382),
.B(n_338),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_338),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_388),
.B(n_342),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_342),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_398),
.A2(n_226),
.B(n_223),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_400),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_387),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_398),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_377),
.A2(n_353),
.B1(n_180),
.B2(n_339),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_353),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_379),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_382),
.B(n_227),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_296),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_371),
.A2(n_309),
.B1(n_296),
.B2(n_228),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_375),
.B(n_230),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_309),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_391),
.B(n_181),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_405),
.A2(n_321),
.B1(n_367),
.B2(n_277),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_369),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_277),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_375),
.B(n_181),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_406),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_182),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_412),
.B(n_369),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_395),
.B(n_185),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_182),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_369),
.B(n_236),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_375),
.B(n_184),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_375),
.B(n_389),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_373),
.Y(n_492)
);

OAI22x1_ASAP7_75t_R g493 ( 
.A1(n_385),
.A2(n_180),
.B1(n_207),
.B2(n_202),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_373),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_399),
.B(n_185),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_410),
.A2(n_210),
.B1(n_192),
.B2(n_233),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_373),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_385),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_389),
.B(n_184),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_390),
.B(n_234),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_389),
.A2(n_236),
.B1(n_235),
.B2(n_234),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_393),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_453),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_453),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_436),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_459),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_459),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_444),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_444),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_466),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_454),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_466),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_455),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_471),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_458),
.B(n_393),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_491),
.B(n_393),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_465),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_469),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_R g531 ( 
.A(n_419),
.B(n_397),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_480),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_471),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_491),
.B(n_393),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_433),
.B(n_396),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_429),
.B(n_385),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_432),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_434),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_434),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_505),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_431),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_470),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_489),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_489),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_489),
.Y(n_549)
);

AND2x2_ASAP7_75t_SL g550 ( 
.A(n_419),
.B(n_396),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_492),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_494),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_428),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_431),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_473),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_435),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_429),
.B(n_385),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_447),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_484),
.B(n_502),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_500),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_450),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_467),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_448),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_423),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_506),
.Y(n_572)
);

BUFx8_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_456),
.C(n_423),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_532),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_564),
.Y(n_579)
);

AOI21x1_ASAP7_75t_L g580 ( 
.A1(n_537),
.A2(n_437),
.B(n_424),
.Y(n_580)
);

AO21x2_ASAP7_75t_L g581 ( 
.A1(n_561),
.A2(n_437),
.B(n_424),
.Y(n_581)
);

AND3x2_ASAP7_75t_L g582 ( 
.A(n_539),
.B(n_420),
.C(n_461),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_564),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_562),
.B(n_458),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_511),
.A2(n_441),
.B(n_452),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_509),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_564),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_509),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_551),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_551),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_526),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_528),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_552),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_542),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_529),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_546),
.B(n_438),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_570),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_571),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_536),
.B(n_438),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_521),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_538),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_548),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_578),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_575),
.A2(n_385),
.B1(n_496),
.B2(n_485),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_590),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_L g620 ( 
.A(n_585),
.B(n_456),
.C(n_472),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_606),
.B(n_566),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_482),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_578),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_610),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_590),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_612),
.A2(n_385),
.B1(n_496),
.B2(n_485),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_449),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_603),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_583),
.B(n_569),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_574),
.B(n_510),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_576),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_576),
.B(n_449),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_596),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_583),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_543),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_583),
.B(n_516),
.Y(n_638)
);

AO21x2_ASAP7_75t_L g639 ( 
.A1(n_587),
.A2(n_580),
.B(n_531),
.Y(n_639)
);

BUFx6f_ASAP7_75t_SL g640 ( 
.A(n_583),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_598),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_517),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_593),
.B(n_518),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

INVx6_ASAP7_75t_L g645 ( 
.A(n_593),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_577),
.B(n_414),
.Y(n_646)
);

BUFx6f_ASAP7_75t_SL g647 ( 
.A(n_593),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_612),
.B(n_519),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_604),
.B(n_414),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_579),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_577),
.B(n_414),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_579),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_608),
.B(n_426),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_605),
.B(n_426),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_609),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_605),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_609),
.B(n_607),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_613),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_613),
.B(n_426),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_592),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_609),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_579),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_592),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_611),
.B(n_558),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_590),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_591),
.B(n_544),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_579),
.B(n_558),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_592),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_590),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_597),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_586),
.B(n_588),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_586),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_601),
.B(n_573),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_588),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_597),
.B(n_555),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_582),
.A2(n_522),
.B1(n_524),
.B2(n_520),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_594),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_SL g686 ( 
.A1(n_601),
.A2(n_500),
.B1(n_553),
.B2(n_556),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_602),
.B(n_547),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_588),
.A2(n_553),
.B1(n_550),
.B2(n_556),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_602),
.B(n_472),
.C(n_481),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_597),
.B(n_560),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_599),
.B(n_550),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_599),
.B(n_559),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_581),
.A2(n_496),
.B1(n_485),
.B2(n_497),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_600),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_597),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_615),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_624),
.B(n_600),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_635),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_641),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_655),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_660),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_621),
.B(n_534),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_687),
.B(n_573),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_637),
.B(n_557),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_648),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_627),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_636),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_663),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_638),
.Y(n_710)
);

XOR2xp5_ASAP7_75t_L g711 ( 
.A(n_686),
.B(n_515),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_643),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_689),
.A2(n_620),
.B(n_617),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_658),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_689),
.A2(n_525),
.B(n_461),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_664),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_687),
.B(n_573),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_673),
.B(n_545),
.Y(n_718)
);

INVxp33_ASAP7_75t_L g719 ( 
.A(n_642),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_665),
.Y(n_720)
);

XOR2x2_ASAP7_75t_SL g721 ( 
.A(n_686),
.B(n_507),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_670),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_681),
.B(n_557),
.Y(n_723)
);

XOR2xp5_ASAP7_75t_L g724 ( 
.A(n_684),
.B(n_565),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_630),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_616),
.B(n_427),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_645),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_624),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_672),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_640),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_657),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_657),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_631),
.B(n_525),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_645),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_657),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_640),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_659),
.Y(n_737)
);

XOR2xp5_ASAP7_75t_L g738 ( 
.A(n_668),
.B(n_565),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_683),
.B(n_600),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_SL g740 ( 
.A(n_647),
.B(n_549),
.Y(n_740)
);

BUFx5_ASAP7_75t_L g741 ( 
.A(n_692),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_647),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_690),
.B(n_540),
.Y(n_743)
);

INVxp33_ASAP7_75t_L g744 ( 
.A(n_671),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_644),
.B(n_488),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_639),
.A2(n_487),
.B(n_476),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_666),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_629),
.B(n_488),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_633),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_654),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_633),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_688),
.B(n_563),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_676),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_680),
.Y(n_754)
);

XOR2xp5_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_541),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_682),
.Y(n_756)
);

BUFx5_ASAP7_75t_L g757 ( 
.A(n_692),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_622),
.B(n_485),
.Y(n_758)
);

XOR2xp5_ASAP7_75t_L g759 ( 
.A(n_693),
.B(n_563),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_616),
.B(n_430),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_694),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_679),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_625),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_679),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_619),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_695),
.B(n_430),
.Y(n_766)
);

XOR2xp5_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_563),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_614),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_618),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_507),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_623),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_662),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_625),
.Y(n_773)
);

XNOR2xp5_ASAP7_75t_L g774 ( 
.A(n_669),
.B(n_501),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_625),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_527),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_667),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_705),
.B(n_728),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_744),
.B(n_634),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_629),
.B(n_661),
.C(n_479),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_710),
.B(n_632),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_750),
.B(n_632),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_733),
.A2(n_485),
.B1(n_496),
.B2(n_527),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_696),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_697),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_712),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_719),
.B(n_654),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_699),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_739),
.B(n_629),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_731),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_700),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_770),
.B(n_691),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_701),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_758),
.B(n_490),
.C(n_479),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_706),
.B(n_235),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_748),
.B(n_675),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_776),
.B(n_490),
.C(n_468),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_749),
.B(n_674),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_751),
.B(n_677),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_743),
.B(n_194),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_702),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_715),
.A2(n_496),
.B(n_468),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_707),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_721),
.B(n_646),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_734),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_725),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_732),
.B(n_581),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_737),
.B(n_685),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_704),
.A2(n_717),
.B(n_752),
.C(n_740),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_734),
.B(n_646),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_714),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_755),
.A2(n_194),
.B1(n_200),
.B2(n_487),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_703),
.B(n_718),
.C(n_745),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_729),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_709),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_734),
.B(n_652),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_716),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_720),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_769),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_698),
.B(n_652),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_740),
.A2(n_493),
.B(n_445),
.C(n_484),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_762),
.B(n_678),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_753),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_711),
.A2(n_194),
.B1(n_200),
.B2(n_568),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_727),
.B(n_695),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_200),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_754),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_764),
.B(n_678),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_723),
.A2(n_527),
.B1(n_535),
.B2(n_501),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_771),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_727),
.B(n_649),
.Y(n_832)
);

BUFx8_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_730),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_723),
.B(n_650),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_736),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_777),
.B(n_656),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_735),
.B(n_675),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_756),
.B(n_651),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_L g840 ( 
.A(n_742),
.B(n_460),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_761),
.B(n_768),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_759),
.B(n_653),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_775),
.B(n_650),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_708),
.B(n_535),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_763),
.B(n_650),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_814),
.B(n_765),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_810),
.B(n_765),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_813),
.A2(n_767),
.B1(n_774),
.B2(n_724),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_813),
.A2(n_747),
.B1(n_760),
.B2(n_726),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_782),
.B(n_779),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_826),
.B(n_773),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_843),
.B(n_781),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_843),
.B(n_741),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_796),
.B(n_773),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_786),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_800),
.B(n_0),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_789),
.B(n_741),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_833),
.B(n_834),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_783),
.B(n_741),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_778),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_792),
.B(n_741),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_835),
.B(n_746),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_793),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_820),
.B(n_757),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_812),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_757),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_827),
.B(n_1),
.Y(n_868)
);

BUFx8_ASAP7_75t_L g869 ( 
.A(n_836),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_833),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_797),
.B(n_757),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_832),
.B(n_757),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_831),
.B(n_757),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_805),
.B(n_766),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_802),
.A2(n_619),
.B(n_587),
.C(n_580),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_790),
.B(n_452),
.Y(n_877)
);

BUFx5_ASAP7_75t_L g878 ( 
.A(n_818),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_787),
.B(n_2),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_832),
.B(n_535),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_788),
.B(n_692),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_785),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_825),
.B(n_370),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_788),
.B(n_692),
.Y(n_884)
);

AND2x6_ASAP7_75t_SL g885 ( 
.A(n_795),
.B(n_460),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_803),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_809),
.B(n_2),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_804),
.A2(n_840),
.B1(n_825),
.B2(n_842),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_794),
.A2(n_370),
.B(n_503),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_791),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_845),
.B(n_3),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_809),
.B(n_4),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_844),
.B(n_584),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_842),
.B(n_5),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_838),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_822),
.A2(n_503),
.B(n_554),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_801),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_821),
.B(n_6),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_815),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_819),
.B(n_7),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_816),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_824),
.B(n_7),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_828),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_806),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_811),
.B(n_8),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_841),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_780),
.A2(n_584),
.B(n_475),
.C(n_440),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_807),
.Y(n_908)
);

INVx8_ASAP7_75t_L g909 ( 
.A(n_839),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_846),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_817),
.B(n_430),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_9),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_829),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_798),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_837),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_838),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_878),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_867),
.B(n_799),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_851),
.B(n_913),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_861),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_857),
.B(n_808),
.C(n_830),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_878),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_914),
.B(n_10),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_883),
.A2(n_440),
.B1(n_475),
.B2(n_378),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_848),
.B(n_559),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_885),
.B(n_10),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_559),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_873),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_878),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_443),
.B(n_417),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_915),
.B(n_11),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_870),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_853),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_457),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_859),
.B(n_457),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_882),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_910),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_871),
.A2(n_476),
.B(n_451),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_847),
.B(n_457),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_890),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_848),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_909),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_856),
.B(n_11),
.Y(n_943)
);

NOR2x1_ASAP7_75t_R g944 ( 
.A(n_898),
.B(n_451),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_879),
.B(n_12),
.C(n_13),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_897),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_906),
.B(n_895),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_899),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_916),
.B(n_12),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_886),
.B(n_13),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_910),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_903),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_864),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_888),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_869),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_863),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_907),
.A2(n_896),
.B(n_849),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_893),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_862),
.B(n_463),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_866),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_904),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_894),
.A2(n_378),
.B(n_498),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_875),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_852),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_861),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_901),
.B(n_14),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_SL g968 ( 
.A1(n_868),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_912),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_928),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_941),
.B(n_905),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_918),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_918),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_956),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_933),
.B(n_947),
.Y(n_976)
);

BUFx8_ASAP7_75t_SL g977 ( 
.A(n_932),
.Y(n_977)
);

BUFx12f_ASAP7_75t_SL g978 ( 
.A(n_932),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_940),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_SL g980 ( 
.A(n_955),
.B(n_850),
.C(n_891),
.Y(n_980)
);

INVx3_ASAP7_75t_SL g981 ( 
.A(n_932),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_919),
.B(n_969),
.Y(n_982)
);

AND3x1_ASAP7_75t_SL g983 ( 
.A(n_968),
.B(n_17),
.C(n_19),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_949),
.B(n_855),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_946),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_965),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_948),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_966),
.B(n_858),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_942),
.B(n_872),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_958),
.A2(n_860),
.B1(n_880),
.B2(n_863),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_964),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_925),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_941),
.B(n_854),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_936),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_942),
.B(n_909),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_937),
.Y(n_996)
);

AO22x1_ASAP7_75t_L g997 ( 
.A1(n_958),
.A2(n_880),
.B1(n_860),
.B2(n_887),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_957),
.B(n_877),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_925),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_957),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_953),
.B(n_892),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_957),
.B(n_925),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_964),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_968),
.B(n_865),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_959),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_SL g1006 ( 
.A(n_955),
.B(n_902),
.C(n_900),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_937),
.B(n_874),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_937),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_954),
.B(n_860),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_961),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_920),
.B(n_881),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_962),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_967),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_927),
.B(n_893),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_952),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_927),
.B(n_917),
.Y(n_1016)
);

CKINVDCx14_ASAP7_75t_R g1017 ( 
.A(n_926),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_967),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_960),
.B(n_884),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_952),
.B(n_875),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_945),
.B(n_889),
.C(n_911),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_945),
.B(n_19),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_952),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_922),
.Y(n_1024)
);

AND3x1_ASAP7_75t_SL g1025 ( 
.A(n_943),
.B(n_20),
.C(n_21),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_950),
.B(n_20),
.C(n_21),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_939),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_939),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_951),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_929),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_970),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_981),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_990),
.A2(n_963),
.B1(n_924),
.B2(n_935),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1000),
.B(n_972),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_1000),
.B(n_921),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_970),
.B(n_931),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_1026),
.A2(n_963),
.B(n_924),
.C(n_923),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_997),
.A2(n_944),
.B(n_934),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_1022),
.A2(n_944),
.B(n_938),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_980),
.A2(n_930),
.B1(n_504),
.B2(n_443),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_991),
.B(n_23),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_980),
.A2(n_504),
.B1(n_417),
.B2(n_451),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1022),
.A2(n_23),
.B(n_24),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1004),
.A2(n_25),
.B(n_26),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1000),
.B(n_451),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1013),
.B(n_25),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1017),
.A2(n_476),
.B1(n_499),
.B2(n_495),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_991),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1037),
.A2(n_1017),
.B1(n_972),
.B2(n_1021),
.Y(n_1049)
);

BUFx4f_ASAP7_75t_L g1050 ( 
.A(n_1032),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1044),
.A2(n_983),
.B1(n_1025),
.B2(n_1026),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_1032),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_1034),
.A2(n_1004),
.B(n_986),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_1031),
.A2(n_998),
.B(n_1024),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1043),
.A2(n_1006),
.B(n_993),
.Y(n_1055)
);

NAND2x1p5_ASAP7_75t_L g1056 ( 
.A(n_1035),
.B(n_1000),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1048),
.B(n_976),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1036),
.B(n_1018),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1041),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1038),
.A2(n_998),
.B(n_1024),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_1039),
.A2(n_993),
.B(n_1007),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1033),
.A2(n_1006),
.B(n_1021),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1045),
.B(n_1003),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1047),
.B(n_1029),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_1042),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_SL g1067 ( 
.A1(n_1040),
.A2(n_1003),
.B(n_982),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1034),
.A2(n_975),
.B(n_1001),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1036),
.B(n_973),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_SL g1070 ( 
.A1(n_1034),
.A2(n_983),
.B(n_1002),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1034),
.A2(n_975),
.B(n_1007),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1044),
.A2(n_1002),
.B(n_1009),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1036),
.B(n_973),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1052),
.B(n_981),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1050),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1052),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1049),
.A2(n_1051),
.B1(n_1063),
.B2(n_1070),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1050),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1059),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1056),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_1068),
.A3(n_1071),
.B(n_1061),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_1078),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_1077),
.B1(n_1051),
.B2(n_1055),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1084),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1083),
.A2(n_1077),
.B1(n_1080),
.B2(n_1075),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1076),
.A3(n_1081),
.B(n_1065),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1074),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1087),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1087),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_1089),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1090),
.B(n_1080),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_1094),
.A2(n_1091),
.B(n_1053),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1093),
.B(n_1072),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1095),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1096),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1097),
.Y(n_1099)
);

NAND2x1_ASAP7_75t_L g1100 ( 
.A(n_1098),
.B(n_1067),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1100),
.B(n_1092),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_1092),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_1102),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_1103),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_1102),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_1104),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1106),
.B(n_1062),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1105),
.B(n_1060),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1109),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_1107),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1108),
.B(n_977),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_1111),
.B(n_1064),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_977),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_1110),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1114),
.Y(n_1116)
);

AO221x2_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_978),
.B1(n_1066),
.B2(n_1058),
.C(n_1005),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_R g1118 ( 
.A(n_1116),
.B(n_26),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1117),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1120),
.B(n_1057),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_1069),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_27),
.Y(n_1123)
);

INVxp67_ASAP7_75t_SL g1124 ( 
.A(n_1122),
.Y(n_1124)
);

INVxp33_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_1073),
.B1(n_1064),
.B2(n_1008),
.Y(n_1126)
);

OAI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1124),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1125),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1126),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1129),
.B(n_28),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1128),
.B(n_29),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1132),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1131),
.B(n_1130),
.Y(n_1134)
);

AOI31xp33_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_31),
.A3(n_32),
.B(n_33),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1133),
.B(n_31),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1136),
.B(n_32),
.C(n_33),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

CKINVDCx6p67_ASAP7_75t_R g1139 ( 
.A(n_1138),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1137),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1140),
.B(n_34),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1139),
.B(n_34),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1142),
.A2(n_1015),
.B(n_1054),
.Y(n_1143)
);

NOR3xp33_ASAP7_75t_SL g1144 ( 
.A(n_1141),
.B(n_38),
.C(n_39),
.Y(n_1144)
);

INVxp33_ASAP7_75t_L g1145 ( 
.A(n_1142),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_408),
.B1(n_1023),
.B2(n_42),
.C(n_45),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_40),
.C(n_41),
.D(n_50),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1143),
.A2(n_1023),
.B1(n_53),
.B2(n_54),
.C(n_55),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1147),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_1148),
.B(n_51),
.C(n_57),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1149),
.A2(n_1146),
.B(n_61),
.C(n_62),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1150),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_SL g1153 ( 
.A(n_1152),
.B(n_59),
.C(n_63),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_1151),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1154),
.B(n_392),
.C(n_384),
.Y(n_1155)
);

OA211x2_ASAP7_75t_L g1156 ( 
.A1(n_1153),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_1156)
);

AO22x2_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1155),
.A2(n_73),
.B(n_74),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_L g1159 ( 
.A(n_1158),
.B(n_75),
.C(n_76),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1157),
.B(n_77),
.C(n_80),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_1159),
.B(n_81),
.C(n_82),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1160),
.B(n_86),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1160),
.B(n_87),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1162),
.Y(n_1164)
);

AND2x2_ASAP7_75t_SL g1165 ( 
.A(n_1163),
.B(n_1161),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_L g1166 ( 
.A(n_1163),
.B(n_88),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1164),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1165),
.Y(n_1168)
);

XNOR2xp5_ASAP7_75t_L g1169 ( 
.A(n_1168),
.B(n_1166),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1167),
.B(n_89),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1169),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1170),
.A2(n_378),
.B1(n_1025),
.B2(n_996),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1171),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1172),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1173),
.Y(n_1175)
);

XNOR2xp5_ASAP7_75t_L g1176 ( 
.A(n_1174),
.B(n_90),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1175),
.Y(n_1177)
);

OAI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1176),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.C(n_96),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1177),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1178),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1177),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1181),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1180),
.A2(n_108),
.B(n_109),
.Y(n_1183)
);

AOI21xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1179),
.A2(n_111),
.B(n_112),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_1184),
.Y(n_1185)
);

CKINVDCx14_ASAP7_75t_R g1186 ( 
.A(n_1182),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1186),
.A2(n_1183),
.B(n_378),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1185),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1188),
.A2(n_995),
.B1(n_1028),
.B2(n_1020),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1188),
.A2(n_113),
.B(n_115),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1189),
.A2(n_116),
.B(n_117),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1191),
.A2(n_118),
.B(n_119),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1190),
.A2(n_380),
.B1(n_999),
.B2(n_992),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1193),
.A2(n_1028),
.B1(n_121),
.B2(n_122),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1194),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1192),
.A2(n_380),
.B1(n_1014),
.B2(n_128),
.Y(n_1197)
);

XNOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_1197),
.B(n_126),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_127),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1195),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1197),
.A2(n_1014),
.B1(n_130),
.B2(n_131),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1196),
.A2(n_129),
.B(n_132),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1196),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_1196),
.A2(n_134),
.B(n_135),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1197),
.B(n_137),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1197),
.A2(n_138),
.B(n_141),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1197),
.B(n_142),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1197),
.A2(n_144),
.B(n_145),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1196),
.A2(n_146),
.B(n_147),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1197),
.A2(n_150),
.B(n_153),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1203),
.A2(n_1200),
.B(n_1199),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1205),
.B(n_154),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1198),
.B(n_155),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1207),
.B(n_156),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1202),
.A2(n_157),
.B(n_158),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1206),
.B(n_1210),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1209),
.A2(n_159),
.B(n_160),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1208),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1204),
.Y(n_1219)
);

AOI322xp5_ASAP7_75t_L g1220 ( 
.A1(n_1218),
.A2(n_1201),
.A3(n_164),
.B1(n_166),
.B2(n_167),
.C1(n_170),
.C2(n_171),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1211),
.A2(n_161),
.B1(n_172),
.B2(n_174),
.Y(n_1221)
);

AOI322xp5_ASAP7_75t_L g1222 ( 
.A1(n_1219),
.A2(n_175),
.A3(n_176),
.B1(n_177),
.B2(n_178),
.C1(n_1027),
.C2(n_989),
.Y(n_1222)
);

AOI222xp33_ASAP7_75t_L g1223 ( 
.A1(n_1216),
.A2(n_1027),
.B1(n_495),
.B2(n_499),
.C1(n_464),
.C2(n_463),
.Y(n_1223)
);

AOI211xp5_ASAP7_75t_L g1224 ( 
.A1(n_1212),
.A2(n_495),
.B(n_464),
.C(n_463),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1215),
.A2(n_499),
.B1(n_464),
.B2(n_384),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1214),
.A2(n_1011),
.B1(n_984),
.B2(n_1016),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1225),
.B(n_1213),
.Y(n_1227)
);

AOI21xp33_ASAP7_75t_L g1228 ( 
.A1(n_1224),
.A2(n_1217),
.B(n_1016),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1220),
.A2(n_1222),
.B(n_1226),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_L g1230 ( 
.A1(n_1229),
.A2(n_1221),
.B1(n_1223),
.B2(n_1012),
.C(n_1010),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1230),
.A2(n_1227),
.B(n_1228),
.C(n_974),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1231),
.A2(n_988),
.B1(n_974),
.B2(n_994),
.Y(n_1232)
);

AOI211xp5_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_1030),
.B(n_1019),
.C(n_979),
.Y(n_1233)
);

AOI211xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_971),
.B(n_987),
.C(n_985),
.Y(n_1234)
);


endmodule