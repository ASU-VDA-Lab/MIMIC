module fake_jpeg_10974_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_23),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_44),
.B(n_46),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_47),
.B(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_2),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_2),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_56),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_70),
.Y(n_83)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_40),
.Y(n_101)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_4),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_20),
.B(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_22),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_7),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_23),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_37),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_31),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_39),
.B1(n_38),
.B2(n_41),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_114),
.B(n_115),
.C(n_87),
.D(n_102),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_29),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_38),
.B1(n_41),
.B2(n_32),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_110),
.B1(n_117),
.B2(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_26),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_26),
.B1(n_36),
.B2(n_32),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_29),
.B1(n_40),
.B2(n_10),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_42),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_9),
.B1(n_12),
.B2(n_48),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_50),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_12),
.B(n_54),
.C(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_129),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_52),
.B1(n_61),
.B2(n_65),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_127),
.B1(n_131),
.B2(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_83),
.A2(n_54),
.B1(n_94),
.B2(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_139),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_101),
.B1(n_114),
.B2(n_100),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_91),
.B1(n_81),
.B2(n_84),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_142),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_90),
.B1(n_115),
.B2(n_95),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_129),
.B(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_95),
.B1(n_85),
.B2(n_86),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_84),
.B1(n_91),
.B2(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_116),
.B1(n_93),
.B2(n_80),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_151),
.B1(n_153),
.B2(n_130),
.Y(n_174)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_116),
.B1(n_93),
.B2(n_80),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_92),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_178),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_181),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_132),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_181),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_137),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_120),
.A2(n_146),
.B(n_145),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_156),
.C(n_163),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_138),
.B1(n_140),
.B2(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_150),
.B1(n_148),
.B2(n_144),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_149),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_168),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_133),
.C(n_135),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_166),
.C(n_180),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_151),
.B1(n_143),
.B2(n_136),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_136),
.B1(n_176),
.B2(n_174),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_167),
.C(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_156),
.B(n_164),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_161),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_209),
.B(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_213),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_167),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_166),
.B(n_160),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_197),
.B(n_190),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_170),
.C(n_157),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_204),
.B1(n_211),
.B2(n_214),
.Y(n_229)
);

AOI221xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_200),
.B1(n_189),
.B2(n_183),
.C(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_224),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_203),
.B1(n_195),
.B2(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_184),
.B(n_183),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_225),
.A2(n_192),
.B1(n_170),
.B2(n_162),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_233),
.B1(n_223),
.B2(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_202),
.B1(n_211),
.B2(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_217),
.B1(n_221),
.B2(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_213),
.C(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_187),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_233),
.A3(n_230),
.B1(n_228),
.B2(n_232),
.C1(n_229),
.C2(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_245),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_234),
.B1(n_186),
.B2(n_196),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_237),
.C(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_246),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_251),
.C(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_244),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_231),
.C(n_206),
.Y(n_254)
);


endmodule