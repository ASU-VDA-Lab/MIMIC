module fake_netlist_5_2527_n_1818 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1818);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1818;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1715;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_84),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_104),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_95),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_11),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_12),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_1),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_26),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_43),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_62),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_58),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_18),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_94),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_36),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_39),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_79),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_64),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_58),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_92),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_116),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_26),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_93),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_35),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_86),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_53),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_154),
.Y(n_229)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_40),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_21),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_38),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_106),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_99),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_0),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_151),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_83),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_70),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_111),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_98),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_43),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g249 ( 
.A(n_126),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_66),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_80),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_135),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_45),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_13),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_51),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_117),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_89),
.Y(n_266)
);

BUFx8_ASAP7_75t_SL g267 ( 
.A(n_122),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_49),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_138),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_56),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_53),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_118),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_29),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_61),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_52),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_29),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_100),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_20),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_132),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_31),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_57),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_107),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_49),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_112),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_153),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_7),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_36),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_55),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_2),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_35),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_72),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_59),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_85),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_51),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_42),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_87),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_28),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_76),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_12),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_24),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_48),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_9),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_38),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_61),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_137),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_23),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_115),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_74),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_88),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_5),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_108),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_23),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_44),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_133),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_140),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_121),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_148),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_134),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_34),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_21),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_5),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_68),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_113),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_163),
.Y(n_335)
);

BUFx4f_ASAP7_75t_SL g336 ( 
.A(n_10),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_130),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_22),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_57),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_103),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_209),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_267),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_172),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_289),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_224),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_328),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_209),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_222),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_222),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_179),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_179),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_175),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_227),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_216),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_216),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_229),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_234),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_173),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_300),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_247),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_197),
.B(n_0),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_247),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_174),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_255),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_271),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_176),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_271),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_273),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_273),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_201),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_193),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_205),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_208),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_1),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_212),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_278),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_278),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_279),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_295),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_242),
.B(n_2),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_183),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_236),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_175),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_295),
.B(n_3),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_254),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_211),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_213),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_262),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_296),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_296),
.Y(n_399)
);

BUFx6f_ASAP7_75t_SL g400 ( 
.A(n_178),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_214),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_215),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_219),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_221),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_303),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_310),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g408 ( 
.A(n_184),
.B(n_4),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_242),
.B(n_6),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_223),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_304),
.B(n_6),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_228),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_235),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_178),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_237),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_238),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_181),
.B(n_7),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_240),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_243),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

AND3x2_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_312),
.C(n_177),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_389),
.B(n_185),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_246),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_359),
.B(n_177),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_353),
.B(n_250),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_344),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_354),
.B(n_340),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_357),
.B(n_251),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_360),
.B(n_178),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_366),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_358),
.B(n_252),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_358),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_361),
.Y(n_446)
);

NOR2x1_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_249),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_364),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_417),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_342),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_370),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_365),
.B(n_258),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_378),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_342),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_350),
.Y(n_463)
);

CKINVDCx6p67_ASAP7_75t_R g464 ( 
.A(n_360),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_350),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_351),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_351),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_371),
.B(n_259),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_352),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_352),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_372),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_347),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_372),
.B(n_288),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_375),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

NAND2x1_ASAP7_75t_L g480 ( 
.A(n_376),
.B(n_207),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_377),
.B(n_263),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_384),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_385),
.B(n_266),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_356),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_363),
.B(n_332),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_356),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_387),
.B(n_312),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_398),
.B(n_275),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g497 ( 
.A1(n_398),
.A2(n_182),
.B(n_181),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_363),
.B(n_335),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_408),
.B1(n_394),
.B2(n_268),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_451),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_435),
.B(n_329),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_369),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_497),
.B1(n_434),
.B2(n_443),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_451),
.B(n_362),
.Y(n_516)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_454),
.B(n_341),
.C(n_233),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_477),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_431),
.B(n_390),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_483),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_493),
.A2(n_393),
.B1(n_285),
.B2(n_277),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_368),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_491),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

CKINVDCx6p67_ASAP7_75t_R g537 ( 
.A(n_464),
.Y(n_537)
);

AND3x1_ASAP7_75t_L g538 ( 
.A(n_490),
.B(n_277),
.C(n_197),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_443),
.A2(n_423),
.B1(n_422),
.B2(n_411),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_447),
.B(n_374),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_438),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_477),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_464),
.B(n_343),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_447),
.B(n_379),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_380),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_477),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_481),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_481),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_433),
.B(n_399),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_457),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_481),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_481),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_481),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_455),
.B(n_381),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_481),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_433),
.B(n_402),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_464),
.B(n_345),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_492),
.B(n_395),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_461),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_455),
.B(n_396),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_473),
.B(n_401),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_490),
.B(n_403),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_404),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g573 ( 
.A(n_492),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_428),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_433),
.B(n_329),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_485),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_428),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_433),
.B(n_182),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_L g580 ( 
.A(n_454),
.B(n_301),
.C(n_200),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_485),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_485),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_448),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_402),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_428),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_495),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_455),
.B(n_405),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_455),
.B(n_413),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_418),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_436),
.B(n_420),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_436),
.B(n_415),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_497),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_448),
.B(n_383),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_495),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_465),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_439),
.B(n_244),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_465),
.Y(n_605)
);

BUFx6f_ASAP7_75t_SL g606 ( 
.A(n_493),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_439),
.B(n_440),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_432),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_437),
.Y(n_610)
);

NOR2x1p5_ASAP7_75t_L g611 ( 
.A(n_440),
.B(n_393),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_465),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_444),
.B(n_400),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_480),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_444),
.B(n_400),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_465),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_437),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_458),
.B(n_281),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_442),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_465),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_458),
.B(n_287),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_407),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_442),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_445),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_445),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_441),
.A2(n_302),
.B1(n_323),
.B2(n_412),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_469),
.B(n_391),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_446),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_482),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_465),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_446),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_462),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_474),
.B(n_407),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_449),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_449),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_450),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_SL g639 ( 
.A(n_499),
.B(n_338),
.C(n_406),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_486),
.B(n_285),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_450),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_486),
.B(n_290),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_462),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_496),
.B(n_336),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_480),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_452),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_462),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_452),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_496),
.B(n_249),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_426),
.B(n_294),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_501),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_501),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_408),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_607),
.B(n_497),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_506),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_636),
.B(n_513),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_504),
.B(n_497),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_508),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_504),
.B(n_427),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_504),
.B(n_467),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_524),
.B(n_187),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_597),
.B(n_186),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_514),
.B(n_207),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_602),
.B(n_188),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_539),
.B(n_192),
.C(n_189),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_611),
.A2(n_298),
.B1(n_325),
.B2(n_337),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_453),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_593),
.B(n_318),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_597),
.A2(n_498),
.B(n_494),
.C(n_460),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_611),
.A2(n_321),
.B1(n_322),
.B2(n_260),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_604),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_619),
.B(n_207),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_609),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_515),
.B(n_230),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_609),
.Y(n_681)
);

AND2x6_ASAP7_75t_SL g682 ( 
.A(n_628),
.B(n_220),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_640),
.B(n_467),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_525),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_618),
.B(n_467),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_510),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_619),
.B(n_207),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_595),
.B(n_265),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_511),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_622),
.B(n_467),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_585),
.B(n_230),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_610),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_470),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_610),
.B(n_617),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_614),
.B(n_646),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_633),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_521),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_585),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_614),
.B(n_207),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_586),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_620),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_620),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_624),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_623),
.B(n_453),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_470),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_531),
.B(n_335),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_633),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_625),
.Y(n_711)
);

BUFx6f_ASAP7_75t_SL g712 ( 
.A(n_650),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_625),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_626),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_623),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_626),
.B(n_470),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_629),
.Y(n_717)
);

NOR2x1_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_225),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_650),
.A2(n_317),
.B1(n_190),
.B2(n_196),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_553),
.B(n_459),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_565),
.B(n_194),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_512),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_614),
.B(n_175),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_542),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_645),
.B(n_627),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_650),
.A2(n_493),
.B1(n_196),
.B2(n_319),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_650),
.A2(n_319),
.B1(n_190),
.B2(n_198),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_644),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_648),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_632),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_565),
.B(n_459),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_540),
.B(n_195),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_547),
.B(n_199),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_632),
.B(n_489),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_203),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_635),
.B(n_489),
.Y(n_736)
);

INVx8_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_512),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_206),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_538),
.B(n_335),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_635),
.B(n_489),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_599),
.A2(n_332),
.B1(n_248),
.B2(n_245),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_614),
.B(n_175),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_575),
.B(n_175),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_637),
.B(n_186),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_634),
.B(n_460),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_519),
.B(n_468),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_614),
.B(n_175),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_634),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_648),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_638),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_638),
.B(n_198),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_646),
.B(n_175),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_646),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_569),
.B(n_232),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_641),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_538),
.B(n_468),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_641),
.B(n_202),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_647),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_613),
.B(n_472),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_647),
.B(n_202),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_646),
.B(n_521),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_650),
.B(n_239),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_553),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_253),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_575),
.B(n_175),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_649),
.B(n_204),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_526),
.B(n_175),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_512),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_651),
.B(n_256),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_536),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_526),
.B(n_231),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_528),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_575),
.A2(n_297),
.B1(n_204),
.B2(n_315),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_528),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_563),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_500),
.A2(n_306),
.B1(n_245),
.B2(n_226),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_563),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_529),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_575),
.A2(n_327),
.B1(n_217),
.B2(n_218),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_573),
.B(n_472),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_532),
.A2(n_333),
.B(n_217),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_579),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_533),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_630),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_533),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_534),
.B(n_210),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_534),
.B(n_210),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_543),
.B(n_231),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_543),
.B(n_218),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_579),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_503),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_502),
.B(n_475),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_536),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_615),
.B(n_226),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_579),
.B(n_241),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_503),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_522),
.B(n_231),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_522),
.B(n_231),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_500),
.B(n_566),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_507),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_606),
.A2(n_269),
.B1(n_334),
.B2(n_333),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_574),
.B(n_241),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_507),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_575),
.A2(n_269),
.B1(n_334),
.B2(n_248),
.Y(n_807)
);

AO221x1_ASAP7_75t_L g808 ( 
.A1(n_505),
.A2(n_257),
.B1(n_280),
.B2(n_284),
.C(n_305),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_639),
.B(n_475),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_578),
.B(n_257),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_575),
.B(n_231),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_509),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_575),
.A2(n_280),
.B1(n_317),
.B2(n_326),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_509),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_578),
.B(n_284),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_518),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_527),
.B(n_476),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_587),
.B(n_305),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_517),
.B(n_476),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_516),
.B(n_261),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_666),
.A2(n_587),
.B1(n_570),
.B2(n_567),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_764),
.A2(n_560),
.B(n_549),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_775),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_700),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_696),
.A2(n_530),
.B(n_536),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_696),
.A2(n_530),
.B(n_592),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_724),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_658),
.Y(n_828)
);

OAI21xp33_ASAP7_75t_L g829 ( 
.A1(n_666),
.A2(n_580),
.B(n_270),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_505),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_669),
.B(n_505),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_669),
.B(n_558),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_656),
.A2(n_530),
.B(n_592),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_802),
.B(n_537),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_659),
.A2(n_558),
.B(n_548),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_764),
.A2(n_590),
.B(n_589),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_702),
.B(n_546),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_663),
.B(n_525),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_668),
.A2(n_530),
.B(n_592),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_668),
.A2(n_592),
.B(n_555),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_SL g841 ( 
.A(n_787),
.B(n_537),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_677),
.A2(n_591),
.B(n_548),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_672),
.B(n_558),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_706),
.B(n_518),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_677),
.A2(n_582),
.B(n_545),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_688),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_725),
.A2(n_306),
.B(n_315),
.C(n_327),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_746),
.B(n_588),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_771),
.A2(n_525),
.B(n_555),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_588),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_682),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_731),
.B(n_525),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_765),
.A2(n_326),
.B(n_288),
.C(n_331),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_676),
.B(n_588),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_722),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_678),
.B(n_594),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_687),
.A2(n_552),
.B(n_545),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_771),
.A2(n_555),
.B(n_525),
.Y(n_858)
);

CKINVDCx8_ASAP7_75t_R g859 ( 
.A(n_664),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_687),
.A2(n_550),
.B1(n_552),
.B2(n_557),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_681),
.B(n_594),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_796),
.A2(n_555),
.B(n_576),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_693),
.B(n_594),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_765),
.A2(n_331),
.B(n_487),
.C(n_478),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_665),
.A2(n_582),
.B(n_550),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_SL g866 ( 
.A1(n_779),
.A2(n_559),
.B(n_600),
.C(n_557),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_795),
.B(n_559),
.Y(n_867)
);

NOR2x1_ASAP7_75t_L g868 ( 
.A(n_809),
.B(n_546),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_747),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_796),
.A2(n_555),
.B(n_562),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_572),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_755),
.B(n_535),
.Y(n_872)
);

AOI33xp33_ASAP7_75t_L g873 ( 
.A1(n_742),
.A2(n_414),
.A3(n_410),
.B1(n_416),
.B2(n_419),
.B3(n_487),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_703),
.B(n_572),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_783),
.B(n_564),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_685),
.A2(n_562),
.B(n_576),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_756),
.A2(n_478),
.B(n_494),
.C(n_484),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_777),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_691),
.A2(n_576),
.B(n_562),
.Y(n_879)
);

CKINVDCx8_ASAP7_75t_R g880 ( 
.A(n_664),
.Y(n_880)
);

AOI21x1_ASAP7_75t_L g881 ( 
.A1(n_723),
.A2(n_748),
.B(n_743),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_704),
.B(n_581),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_715),
.B(n_749),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_766),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_705),
.B(n_581),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_679),
.B(n_554),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_759),
.A2(n_498),
.B(n_479),
.C(n_484),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_778),
.B(n_479),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_694),
.A2(n_562),
.B(n_576),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_756),
.A2(n_410),
.B(n_414),
.C(n_416),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_755),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_781),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_757),
.B(n_535),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_684),
.A2(n_576),
.B(n_562),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_692),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_785),
.A2(n_523),
.B(n_520),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_711),
.B(n_583),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_664),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_757),
.A2(n_523),
.B(n_520),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_713),
.B(n_583),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_683),
.A2(n_523),
.B(n_520),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_674),
.A2(n_596),
.B(n_600),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_721),
.B(n_332),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_732),
.A2(n_419),
.B(n_272),
.C(n_264),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_654),
.B(n_274),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_714),
.B(n_596),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_707),
.A2(n_561),
.B(n_541),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_717),
.B(n_541),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_781),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_793),
.A2(n_598),
.B1(n_551),
.B2(n_556),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_735),
.B(n_544),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_819),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_730),
.B(n_544),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_750),
.B(n_551),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_752),
.B(n_556),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_695),
.B(n_561),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_719),
.A2(n_598),
.B(n_571),
.C(n_577),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_773),
.A2(n_743),
.B(n_723),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_773),
.A2(n_523),
.B(n_520),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_786),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_817),
.A2(n_584),
.B(n_571),
.C(n_577),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_732),
.A2(n_320),
.B(n_282),
.C(n_283),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_720),
.B(n_584),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_735),
.B(n_276),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_SL g926 ( 
.A(n_737),
.B(n_286),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_758),
.B(n_603),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_780),
.A2(n_603),
.B1(n_621),
.B2(n_631),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_761),
.B(n_603),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_720),
.B(n_621),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_797),
.A2(n_601),
.B(n_616),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_748),
.A2(n_523),
.B(n_520),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_754),
.A2(n_736),
.B(n_734),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_767),
.B(n_621),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_754),
.A2(n_523),
.B(n_520),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_601),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_716),
.A2(n_605),
.B(n_631),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_745),
.A2(n_616),
.B(n_612),
.C(n_605),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_767),
.B(n_612),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_673),
.B(n_772),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_722),
.A2(n_643),
.B(n_471),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_772),
.A2(n_643),
.B1(n_231),
.B2(n_466),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_667),
.A2(n_643),
.B(n_471),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_667),
.A2(n_643),
.B(n_466),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_667),
.B(n_643),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_721),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_698),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_739),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_667),
.B(n_466),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_722),
.A2(n_463),
.B(n_456),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_722),
.A2(n_463),
.B(n_456),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_739),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_738),
.A2(n_768),
.B(n_744),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_667),
.B(n_463),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_738),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_738),
.A2(n_456),
.B(n_339),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_738),
.A2(n_811),
.B(n_741),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_794),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_762),
.B(n_753),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_701),
.A2(n_316),
.B(n_314),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_760),
.B(n_231),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_701),
.A2(n_313),
.B(n_311),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_737),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_708),
.A2(n_231),
.B(n_308),
.C(n_307),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_784),
.A2(n_309),
.B(n_299),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_698),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_820),
.B(n_293),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_794),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_712),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_709),
.Y(n_970)
);

AO21x1_ASAP7_75t_L g971 ( 
.A1(n_733),
.A2(n_231),
.B(n_9),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_718),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_733),
.A2(n_8),
.B(n_10),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_820),
.A2(n_292),
.B(n_291),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_709),
.A2(n_169),
.B(n_155),
.Y(n_975)
);

INVx11_ASAP7_75t_L g976 ( 
.A(n_798),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_670),
.B(n_8),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_740),
.B(n_13),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_710),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_710),
.A2(n_152),
.B(n_146),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_763),
.A2(n_769),
.B(n_789),
.C(n_790),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_728),
.A2(n_144),
.B(n_142),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_728),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_799),
.B(n_14),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_803),
.B(n_15),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_812),
.B(n_816),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_729),
.B(n_109),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_699),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_729),
.A2(n_105),
.B(n_101),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_751),
.A2(n_96),
.B(n_77),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_751),
.A2(n_69),
.B(n_65),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_726),
.B(n_15),
.Y(n_992)
);

O2A1O1Ixp5_ASAP7_75t_L g993 ( 
.A1(n_805),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_770),
.A2(n_19),
.B(n_20),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_806),
.B(n_22),
.Y(n_995)
);

O2A1O1Ixp5_ASAP7_75t_L g996 ( 
.A1(n_810),
.A2(n_24),
.B(n_27),
.C(n_30),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_806),
.B(n_27),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_814),
.A2(n_30),
.B(n_32),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_671),
.B(n_32),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_798),
.A2(n_712),
.B1(n_699),
.B2(n_675),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_699),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_814),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_652),
.B(n_33),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_652),
.A2(n_33),
.B(n_34),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_770),
.A2(n_37),
.B(n_40),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_953),
.A2(n_776),
.B(n_807),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_SL g1007 ( 
.A1(n_828),
.A2(n_851),
.B1(n_846),
.B2(n_948),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_957),
.A2(n_776),
.B(n_807),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_946),
.A2(n_782),
.B1(n_727),
.B2(n_804),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_911),
.B(n_792),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_869),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_833),
.A2(n_839),
.B(n_832),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_911),
.B(n_662),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_925),
.A2(n_818),
.B(n_815),
.C(n_791),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_925),
.A2(n_774),
.B(n_791),
.C(n_801),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_823),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_823),
.Y(n_1017)
);

BUFx4f_ASAP7_75t_L g1018 ( 
.A(n_837),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_878),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_952),
.B(n_657),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_913),
.Y(n_1021)
);

AOI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_940),
.A2(n_774),
.B(n_801),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_SL g1023 ( 
.A(n_969),
.B(n_800),
.C(n_808),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_830),
.B(n_653),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_883),
.B(n_813),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_883),
.B(n_699),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_998),
.A2(n_653),
.B1(n_690),
.B2(n_689),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_898),
.B(n_699),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_831),
.A2(n_680),
.B(n_657),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_824),
.B(n_686),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_867),
.B(n_798),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_907),
.A2(n_686),
.B(n_660),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_884),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_829),
.A2(n_800),
.B1(n_690),
.B2(n_689),
.C(n_680),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_923),
.A2(n_662),
.B(n_660),
.C(n_655),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_798),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_867),
.B(n_798),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_958),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_855),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_838),
.A2(n_842),
.B(n_836),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_967),
.B(n_655),
.Y(n_1041)
);

INVx6_ASAP7_75t_L g1042 ( 
.A(n_936),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_958),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_884),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_855),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_904),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_968),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_844),
.B(n_46),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_904),
.A2(n_978),
.B(n_923),
.C(n_903),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_978),
.A2(n_46),
.B(n_47),
.C(n_50),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_992),
.A2(n_50),
.B(n_52),
.C(n_54),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_919),
.A2(n_54),
.B(n_55),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_SL g1053 ( 
.A1(n_834),
.A2(n_60),
.B1(n_63),
.B2(n_827),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_912),
.B(n_60),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_826),
.A2(n_63),
.B(n_840),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_859),
.B(n_880),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_963),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_968),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_SL g1059 ( 
.A1(n_834),
.A2(n_999),
.B1(n_868),
.B2(n_895),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_895),
.B(n_905),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_825),
.A2(n_934),
.B(n_879),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_837),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_892),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_875),
.B(n_972),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_959),
.B(n_848),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_843),
.B(n_939),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_886),
.B(n_888),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_963),
.B(n_1001),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1004),
.A2(n_1000),
.B1(n_877),
.B2(n_986),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_1001),
.B(n_988),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_864),
.A2(n_987),
.B(n_877),
.C(n_853),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_977),
.Y(n_1072)
);

BUFx8_ASAP7_75t_L g1073 ( 
.A(n_888),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_909),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_841),
.B(n_926),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_855),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_970),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_876),
.A2(n_889),
.B(n_849),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_936),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_855),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_858),
.A2(n_835),
.B(n_981),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1002),
.B(n_921),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_947),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_966),
.Y(n_1084)
);

CKINVDCx14_ASAP7_75t_R g1085 ( 
.A(n_936),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_862),
.A2(n_870),
.B(n_865),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_983),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_979),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_SL g1089 ( 
.A1(n_990),
.A2(n_991),
.B(n_847),
.C(n_902),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_992),
.A2(n_864),
.B(n_853),
.C(n_985),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_891),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_974),
.A2(n_965),
.B(n_887),
.C(n_873),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_955),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_930),
.B(n_924),
.Y(n_1096)
);

CKINVDCx8_ASAP7_75t_R g1097 ( 
.A(n_955),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_845),
.A2(n_857),
.B(n_852),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_971),
.A2(n_973),
.B1(n_924),
.B2(n_984),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_988),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_891),
.Y(n_1101)
);

NAND3x1_ASAP7_75t_L g1102 ( 
.A(n_993),
.B(n_996),
.C(n_1005),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_852),
.A2(n_894),
.B(n_838),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_822),
.A2(n_917),
.B(n_933),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1003),
.Y(n_1105)
);

AO21x1_ASAP7_75t_L g1106 ( 
.A1(n_987),
.A2(n_860),
.B(n_917),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_908),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_914),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_872),
.A2(n_893),
.B(n_901),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_881),
.B(n_897),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_960),
.B(n_962),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_890),
.A2(n_866),
.B(n_995),
.C(n_997),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_871),
.B(n_900),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_890),
.A2(n_976),
.B1(n_928),
.B2(n_906),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_SL g1115 ( 
.A(n_945),
.B(n_994),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_872),
.A2(n_893),
.B(n_954),
.C(n_949),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_915),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_874),
.A2(n_885),
.B1(n_882),
.B2(n_916),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_850),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_854),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_922),
.A2(n_964),
.B(n_918),
.C(n_938),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_856),
.A2(n_929),
.B1(n_861),
.B2(n_863),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_927),
.A2(n_942),
.B1(n_821),
.B2(n_910),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_961),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_866),
.A2(n_956),
.B(n_931),
.C(n_937),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_SL g1126 ( 
.A1(n_943),
.A2(n_944),
.B(n_896),
.C(n_989),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_950),
.B(n_951),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_920),
.A2(n_932),
.B(n_935),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_941),
.B(n_975),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_899),
.A2(n_980),
.B(n_982),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_946),
.B(n_607),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_946),
.B(n_607),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_1001),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_824),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_953),
.A2(n_696),
.B(n_957),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_905),
.B(n_654),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_925),
.A2(n_666),
.B(n_658),
.C(n_940),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_925),
.A2(n_666),
.B(n_658),
.C(n_940),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_946),
.B(n_607),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_823),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_827),
.B(n_542),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_953),
.A2(n_696),
.B(n_957),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_827),
.B(n_542),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_946),
.B(n_607),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_946),
.B(n_607),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_SL g1146 ( 
.A(n_925),
.B(n_666),
.C(n_658),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_SL g1147 ( 
.A1(n_828),
.A2(n_500),
.B1(n_851),
.B2(n_846),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_907),
.A2(n_937),
.B(n_879),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_823),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_855),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_953),
.A2(n_696),
.B(n_957),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_L g1152 ( 
.A(n_925),
.B(n_539),
.C(n_666),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_946),
.B(n_948),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_925),
.B(n_666),
.C(n_658),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_824),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_828),
.B(n_658),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1032),
.A2(n_1142),
.B(n_1135),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1082),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1081),
.A2(n_1012),
.B(n_1089),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1057),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1151),
.A2(n_1148),
.B(n_1128),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1106),
.A2(n_1069),
.A3(n_1121),
.B(n_1123),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1017),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_1138),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1082),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1115),
.A2(n_1040),
.B(n_1104),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1146),
.A2(n_1152),
.B(n_1154),
.C(n_1049),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1083),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1086),
.A2(n_1113),
.B(n_1006),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1078),
.A2(n_1109),
.B(n_1029),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1069),
.A2(n_1123),
.A3(n_1110),
.B(n_1061),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1156),
.B(n_1060),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1098),
.A2(n_1102),
.B(n_1090),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1033),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1113),
.A2(n_1066),
.B(n_1126),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1097),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1084),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1072),
.B(n_1136),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1066),
.A2(n_1008),
.B(n_1010),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_1068),
.B(n_1042),
.Y(n_1182)
);

AOI221x1_ASAP7_75t_L g1183 ( 
.A1(n_1052),
.A2(n_1046),
.B1(n_1055),
.B2(n_1114),
.C(n_1094),
.Y(n_1183)
);

NAND3x1_ASAP7_75t_L g1184 ( 
.A(n_1067),
.B(n_1132),
.C(n_1145),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1103),
.A2(n_1130),
.B(n_1127),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1131),
.B(n_1139),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1013),
.A2(n_1122),
.B(n_1027),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_SL g1188 ( 
.A(n_1053),
.B(n_1018),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1027),
.A2(n_1114),
.A3(n_1122),
.B(n_1118),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1133),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1144),
.B(n_1145),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1039),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1141),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1130),
.A2(n_1127),
.B(n_1035),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1016),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1065),
.B(n_1041),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1112),
.A2(n_1125),
.B(n_1010),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1065),
.B(n_1108),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1134),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1050),
.A2(n_1153),
.B(n_1051),
.C(n_1054),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1039),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1015),
.A2(n_1071),
.B(n_1099),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1118),
.A2(n_1013),
.B(n_1014),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1037),
.A2(n_1111),
.B(n_1024),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1024),
.A2(n_1116),
.B(n_1129),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1096),
.A2(n_1009),
.B(n_1048),
.C(n_1022),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1155),
.B(n_1044),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1124),
.A2(n_1022),
.B(n_1025),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1020),
.B(n_1120),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1073),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1059),
.B(n_1011),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1048),
.A2(n_1034),
.B(n_1140),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1019),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1119),
.A2(n_1105),
.B(n_1009),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1105),
.A2(n_1064),
.B(n_1026),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1021),
.A2(n_1047),
.B(n_1038),
.C(n_1043),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1030),
.B(n_1018),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1105),
.A2(n_1026),
.B(n_1133),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1088),
.B(n_1074),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1058),
.A2(n_1149),
.A3(n_1063),
.B(n_1077),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1073),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1091),
.A2(n_1101),
.B(n_1087),
.C(n_1095),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1023),
.A2(n_1036),
.B(n_1028),
.C(n_1100),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1045),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1147),
.A2(n_1075),
.B1(n_1007),
.B2(n_1143),
.C(n_1079),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1028),
.B(n_1036),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_1070),
.B(n_1068),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_1080),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1092),
.A2(n_1042),
.B(n_1085),
.C(n_1076),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1039),
.A2(n_1080),
.B(n_1093),
.C(n_1150),
.Y(n_1232)
);

AO22x2_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_1056),
.B1(n_1092),
.B2(n_1080),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1093),
.A2(n_1138),
.B1(n_1137),
.B2(n_779),
.C(n_1050),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1093),
.A2(n_1081),
.B(n_1032),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1150),
.A2(n_1081),
.B(n_1089),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1106),
.A2(n_931),
.A3(n_1069),
.B(n_1121),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

AO32x2_ASAP7_75t_L g1241 ( 
.A1(n_1069),
.A2(n_1059),
.A3(n_1027),
.B1(n_1114),
.B2(n_1118),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1089),
.C(n_1049),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1243)
);

OAI22x1_ASAP7_75t_L g1244 ( 
.A1(n_1154),
.A2(n_828),
.B1(n_1072),
.B2(n_952),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1245)
);

BUFx8_ASAP7_75t_L g1246 ( 
.A(n_1062),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1081),
.A2(n_1032),
.B(n_1148),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1146),
.A2(n_1152),
.B1(n_1154),
.B2(n_666),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1097),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1154),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1082),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1134),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1097),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1146),
.A2(n_1152),
.B1(n_1154),
.B2(n_666),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1106),
.A2(n_931),
.A3(n_1069),
.B(n_1121),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1134),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1154),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1011),
.B(n_827),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1264)
);

AOI221xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_779),
.B2(n_1050),
.C(n_1051),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1154),
.A2(n_1137),
.B1(n_1138),
.B2(n_504),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1097),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1156),
.B(n_828),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1146),
.A2(n_1152),
.B1(n_1154),
.B2(n_666),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1089),
.C(n_1049),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1154),
.B(n_828),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1097),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1154),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1156),
.B(n_828),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1031),
.A2(n_977),
.B(n_940),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1097),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1082),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1154),
.B2(n_666),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1154),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1156),
.B(n_828),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1154),
.B2(n_666),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1146),
.A2(n_1152),
.B1(n_1154),
.B2(n_666),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1082),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1154),
.B(n_828),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1082),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1082),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1097),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1151),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1134),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1032),
.A2(n_907),
.B(n_1135),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1031),
.A2(n_977),
.B(n_940),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1069),
.A2(n_1059),
.A3(n_1027),
.B1(n_1114),
.B2(n_1118),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1097),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1161),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1209),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1200),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1200),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1179),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1284),
.A2(n_1287),
.B1(n_1253),
.B2(n_1276),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_SL g1315 ( 
.A(n_1178),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1192),
.B(n_1158),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1253),
.A2(n_1285),
.B1(n_1276),
.B2(n_1262),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1237),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1270),
.A2(n_1286),
.B1(n_1279),
.B2(n_1174),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1248),
.A2(n_1290),
.B1(n_1259),
.B2(n_1271),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1293),
.B1(n_1291),
.B2(n_1267),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1178),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1268),
.B(n_1288),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1215),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1248),
.A2(n_1290),
.B1(n_1271),
.B2(n_1259),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1196),
.Y(n_1326)
);

OAI22x1_ASAP7_75t_L g1327 ( 
.A1(n_1273),
.A2(n_1295),
.B1(n_1213),
.B2(n_1219),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1188),
.A2(n_1266),
.B1(n_1262),
.B2(n_1285),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1165),
.A2(n_1266),
.B1(n_1188),
.B2(n_1203),
.Y(n_1329)
);

BUFx10_ASAP7_75t_L g1330 ( 
.A(n_1178),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1255),
.Y(n_1331)
);

BUFx4_ASAP7_75t_R g1332 ( 
.A(n_1166),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1203),
.A2(n_1165),
.B1(n_1198),
.B2(n_1175),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_SL g1334 ( 
.A(n_1250),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1212),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1240),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1261),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1250),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1211),
.A2(n_1199),
.B1(n_1159),
.B2(n_1254),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_1244),
.B1(n_1175),
.B2(n_1167),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1283),
.A2(n_1296),
.B1(n_1299),
.B2(n_1294),
.Y(n_1341)
);

BUFx2_ASAP7_75t_SL g1342 ( 
.A(n_1256),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1180),
.A2(n_1233),
.B1(n_1306),
.B2(n_1241),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1204),
.A2(n_1216),
.B1(n_1181),
.B2(n_1171),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1256),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1225),
.A2(n_1182),
.B1(n_1184),
.B2(n_1207),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1221),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1303),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1208),
.A2(n_1182),
.B1(n_1183),
.B2(n_1176),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1177),
.A2(n_1210),
.B1(n_1208),
.B2(n_1239),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1233),
.A2(n_1241),
.B1(n_1306),
.B2(n_1307),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1269),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1194),
.A2(n_1223),
.B1(n_1182),
.B2(n_1269),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1241),
.A2(n_1306),
.B1(n_1307),
.B2(n_1282),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1201),
.A2(n_1217),
.B1(n_1169),
.B2(n_1263),
.Y(n_1355)
);

INVx6_ASAP7_75t_L g1356 ( 
.A(n_1274),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1238),
.A2(n_1281),
.B1(n_1257),
.B2(n_1302),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1227),
.A2(n_1258),
.B1(n_1300),
.B2(n_1228),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1246),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1222),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1222),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1282),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1243),
.A2(n_1245),
.B1(n_1278),
.B2(n_1289),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1222),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1282),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1307),
.A2(n_1301),
.B1(n_1265),
.B2(n_1246),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1301),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1220),
.A2(n_1301),
.B1(n_1206),
.B2(n_1229),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1193),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1292),
.A2(n_1298),
.B(n_1297),
.Y(n_1370)
);

OAI22x1_ASAP7_75t_SL g1371 ( 
.A1(n_1193),
.A2(n_1226),
.B1(n_1190),
.B2(n_1231),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1202),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1234),
.B(n_1265),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1202),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1218),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1160),
.A2(n_1214),
.B1(n_1236),
.B2(n_1205),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1280),
.Y(n_1377)
);

INVx4_ASAP7_75t_SL g1378 ( 
.A(n_1163),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1242),
.A2(n_1272),
.B1(n_1234),
.B2(n_1214),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1195),
.A2(n_1185),
.B1(n_1235),
.B2(n_1230),
.Y(n_1380)
);

INVx8_ASAP7_75t_L g1381 ( 
.A(n_1232),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1163),
.B(n_1173),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1247),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1247),
.A2(n_1189),
.B1(n_1172),
.B2(n_1157),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1305),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1224),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1162),
.A2(n_1252),
.B1(n_1277),
.B2(n_1275),
.Y(n_1387)
);

CKINVDCx6p67_ASAP7_75t_R g1388 ( 
.A(n_1168),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1173),
.B(n_1189),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1189),
.A2(n_1249),
.B1(n_1251),
.B2(n_1264),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1173),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1260),
.A2(n_1053),
.B1(n_490),
.B2(n_1188),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1304),
.A2(n_1152),
.B1(n_1146),
.B2(n_1154),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1187),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1170),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1178),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1284),
.A2(n_1152),
.B1(n_1146),
.B2(n_1154),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1194),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1170),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1270),
.A2(n_1154),
.B1(n_828),
.B2(n_1156),
.Y(n_1403)
);

BUFx12f_ASAP7_75t_L g1404 ( 
.A(n_1246),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1178),
.Y(n_1405)
);

CKINVDCx14_ASAP7_75t_R g1406 ( 
.A(n_1194),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1188),
.A2(n_1154),
.B1(n_1146),
.B2(n_828),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1194),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1255),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1284),
.A2(n_1152),
.B1(n_1146),
.B2(n_1154),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1188),
.A2(n_1053),
.B1(n_490),
.B2(n_1154),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1178),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1178),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1164),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1270),
.A2(n_1154),
.B1(n_828),
.B2(n_1156),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1194),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1255),
.Y(n_1417)
);

INVx4_ASAP7_75t_L g1418 ( 
.A(n_1178),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1188),
.A2(n_1053),
.B1(n_490),
.B2(n_1154),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1188),
.A2(n_490),
.B1(n_925),
.B2(n_666),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1188),
.A2(n_1053),
.B1(n_490),
.B2(n_1154),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1188),
.A2(n_490),
.B1(n_925),
.B2(n_666),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1284),
.A2(n_1152),
.B1(n_1146),
.B2(n_1154),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1360),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1382),
.B(n_1343),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1361),
.Y(n_1426)
);

CKINVDCx11_ASAP7_75t_R g1427 ( 
.A(n_1404),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1339),
.B(n_1321),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1364),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1339),
.B(n_1317),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1370),
.A2(n_1363),
.B(n_1357),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1391),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1411),
.A2(n_1419),
.B1(n_1421),
.B2(n_1392),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1420),
.A2(n_1422),
.B1(n_1319),
.B2(n_1355),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1393),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1318),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1344),
.A2(n_1390),
.B(n_1363),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1343),
.B(n_1351),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1336),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1317),
.B(n_1308),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1311),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1344),
.A2(n_1390),
.B(n_1357),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1395),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1411),
.A2(n_1419),
.B1(n_1421),
.B2(n_1392),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1312),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1389),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1351),
.B(n_1320),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1383),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1348),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1378),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1310),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1325),
.B(n_1340),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1387),
.A2(n_1375),
.B(n_1349),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1326),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_SL g1456 ( 
.A1(n_1407),
.A2(n_1323),
.B(n_1403),
.C(n_1415),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1349),
.A2(n_1346),
.B(n_1373),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1313),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1388),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1397),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1369),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1402),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1377),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1333),
.B(n_1316),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1376),
.A2(n_1384),
.B(n_1350),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1354),
.B(n_1333),
.Y(n_1466)
);

OAI31xp33_ASAP7_75t_L g1467 ( 
.A1(n_1407),
.A2(n_1423),
.A3(n_1410),
.B(n_1400),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1377),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1324),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1385),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1354),
.B(n_1328),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1384),
.A2(n_1380),
.B(n_1376),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1379),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1379),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1331),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1350),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1328),
.B(n_1340),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1409),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1368),
.A2(n_1314),
.B(n_1329),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1386),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1347),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1381),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1329),
.B(n_1314),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1381),
.Y(n_1485)
);

AO22x2_ASAP7_75t_L g1486 ( 
.A1(n_1366),
.A2(n_1423),
.B1(n_1400),
.B2(n_1410),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1394),
.A2(n_1341),
.B(n_1414),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1417),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1341),
.A2(n_1358),
.B(n_1366),
.Y(n_1489)
);

BUFx4f_ASAP7_75t_SL g1490 ( 
.A(n_1401),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1327),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1371),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1353),
.A2(n_1374),
.B(n_1372),
.Y(n_1493)
);

OAI21xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1322),
.A2(n_1418),
.B(n_1398),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1352),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1322),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1338),
.B(n_1365),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1315),
.A2(n_1332),
.B(n_1345),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1342),
.B(n_1365),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1428),
.B(n_1464),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1472),
.A2(n_1315),
.B(n_1413),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1498),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1491),
.B(n_1425),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1413),
.Y(n_1504)
);

AND2x2_ASAP7_75t_SL g1505 ( 
.A(n_1477),
.B(n_1367),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1425),
.B(n_1337),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1441),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1458),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_R g1509 ( 
.A(n_1470),
.B(n_1334),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1455),
.B(n_1362),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1475),
.B(n_1405),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_SL g1513 ( 
.A(n_1428),
.B(n_1406),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1479),
.A2(n_1416),
.B(n_1408),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1467),
.A2(n_1359),
.B(n_1412),
.C(n_1356),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1467),
.A2(n_1412),
.B(n_1356),
.C(n_1330),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1444),
.A2(n_1412),
.B1(n_1335),
.B2(n_1309),
.Y(n_1517)
);

OR2x6_ASAP7_75t_L g1518 ( 
.A(n_1432),
.B(n_1335),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1519)
);

AO32x2_ASAP7_75t_L g1520 ( 
.A1(n_1483),
.A2(n_1461),
.A3(n_1466),
.B1(n_1438),
.B2(n_1457),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1448),
.B(n_1478),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1460),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_1451),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1434),
.A2(n_1444),
.B1(n_1433),
.B2(n_1456),
.C(n_1453),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1464),
.B(n_1430),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1483),
.B(n_1463),
.Y(n_1526)
);

NAND4xp25_ASAP7_75t_L g1527 ( 
.A(n_1453),
.B(n_1430),
.C(n_1477),
.D(n_1484),
.Y(n_1527)
);

AO32x2_ASAP7_75t_L g1528 ( 
.A1(n_1483),
.A2(n_1466),
.A3(n_1438),
.B1(n_1457),
.B2(n_1471),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1484),
.A2(n_1471),
.B(n_1492),
.C(n_1482),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1427),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1486),
.A2(n_1473),
.B1(n_1474),
.B2(n_1440),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1445),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1450),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1487),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1439),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_R g1536 ( 
.A(n_1470),
.B(n_1480),
.Y(n_1536)
);

AND2x2_ASAP7_75t_SL g1537 ( 
.A(n_1463),
.B(n_1489),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1538)
);

OAI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1437),
.A2(n_1442),
.B(n_1476),
.Y(n_1539)
);

BUFx8_ASAP7_75t_SL g1540 ( 
.A(n_1480),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1437),
.A2(n_1442),
.B(n_1489),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1469),
.B(n_1457),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1446),
.B(n_1443),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_L g1544 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1486),
.A2(n_1489),
.B1(n_1485),
.B2(n_1482),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1459),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_SL g1547 ( 
.A1(n_1480),
.A2(n_1470),
.B(n_1497),
.C(n_1468),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1489),
.A2(n_1431),
.B(n_1487),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1486),
.A2(n_1485),
.B1(n_1482),
.B2(n_1480),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1534),
.B(n_1446),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1508),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1542),
.B(n_1472),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1541),
.B(n_1472),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1541),
.B(n_1465),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1522),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1510),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1424),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1500),
.B(n_1525),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1449),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1524),
.A2(n_1486),
.B1(n_1505),
.B2(n_1514),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1548),
.B(n_1436),
.Y(n_1564)
);

AND2x4_ASAP7_75t_SL g1565 ( 
.A(n_1523),
.B(n_1432),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1502),
.B(n_1426),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1543),
.Y(n_1567)
);

NAND2x1_ASAP7_75t_L g1568 ( 
.A(n_1502),
.B(n_1501),
.Y(n_1568)
);

INVx11_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1528),
.B(n_1429),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1543),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1528),
.B(n_1429),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1531),
.B(n_1462),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1570),
.B(n_1501),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1573),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1566),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1551),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1551),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1570),
.B(n_1528),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1551),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1570),
.B(n_1548),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1569),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1563),
.A2(n_1527),
.B1(n_1544),
.B2(n_1457),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1572),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1572),
.B(n_1503),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1572),
.B(n_1555),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1555),
.B(n_1537),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1565),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1538),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1507),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.Y(n_1593)
);

AOI211xp5_ASAP7_75t_L g1594 ( 
.A1(n_1553),
.A2(n_1514),
.B(n_1515),
.C(n_1527),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1563),
.A2(n_1517),
.B1(n_1549),
.B2(n_1545),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1558),
.B(n_1545),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1558),
.B(n_1454),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1454),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1550),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1556),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1521),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1565),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1575),
.B(n_1561),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1575),
.B(n_1599),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1580),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1582),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1580),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1583),
.A2(n_1549),
.B1(n_1504),
.B2(n_1554),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1599),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_1583),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1592),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1584),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1592),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1592),
.Y(n_1617)
);

INVxp33_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1577),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1588),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1601),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1577),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1600),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1579),
.B(n_1559),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1552),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1593),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1578),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1582),
.B(n_1568),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1593),
.B(n_1579),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1594),
.B(n_1526),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1576),
.B(n_1565),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1600),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1552),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1609),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1591),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1626),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1626),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1604),
.B(n_1622),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1635),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1591),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1636),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1606),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1628),
.B(n_1596),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1620),
.B(n_1581),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1636),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1620),
.Y(n_1655)
);

NOR3xp33_ASAP7_75t_L g1656 ( 
.A(n_1610),
.B(n_1594),
.C(n_1582),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1633),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1619),
.Y(n_1659)
);

AO21x1_ASAP7_75t_L g1660 ( 
.A1(n_1633),
.A2(n_1596),
.B(n_1581),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1613),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1574),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1574),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1610),
.A2(n_1595),
.B1(n_1529),
.B2(n_1504),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1597),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1622),
.B(n_1601),
.Y(n_1668)
);

NAND2x1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_1631),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1621),
.B(n_1557),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1613),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1597),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1611),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1610),
.A2(n_1595),
.B1(n_1504),
.B2(n_1526),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1619),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1631),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1631),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1625),
.B(n_1598),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1657),
.B(n_1582),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1618),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1659),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1655),
.B(n_1618),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1665),
.A2(n_1608),
.B(n_1606),
.C(n_1573),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1648),
.B(n_1623),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1658),
.B(n_1637),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1665),
.A2(n_1608),
.B(n_1553),
.C(n_1598),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1637),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1660),
.A2(n_1553),
.B1(n_1598),
.B2(n_1554),
.C(n_1606),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1659),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1645),
.B(n_1647),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1650),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1651),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1668),
.B(n_1624),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1662),
.Y(n_1701)
);

OAI31xp33_ASAP7_75t_L g1702 ( 
.A1(n_1650),
.A2(n_1506),
.A3(n_1554),
.B(n_1546),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1639),
.B(n_1557),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1638),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1646),
.B(n_1585),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1660),
.A2(n_1606),
.B(n_1513),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1661),
.Y(n_1710)
);

NAND2x1_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1606),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1670),
.B(n_1668),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1674),
.A2(n_1606),
.B1(n_1432),
.B2(n_1435),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1669),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1677),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1684),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1687),
.A2(n_1674),
.B1(n_1642),
.B2(n_1649),
.C(n_1654),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1707),
.B(n_1650),
.Y(n_1720)
);

INVxp67_ASAP7_75t_SL g1721 ( 
.A(n_1715),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1653),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1691),
.A2(n_1678),
.B1(n_1669),
.B2(n_1509),
.C(n_1654),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1696),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1712),
.B(n_1672),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1681),
.B(n_1682),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1713),
.A2(n_1649),
.B1(n_1519),
.B2(n_1679),
.C(n_1511),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1706),
.B(n_1569),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1696),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1695),
.A2(n_1709),
.B1(n_1703),
.B2(n_1699),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1701),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1702),
.A2(n_1644),
.B(n_1676),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1715),
.A2(n_1644),
.B1(n_1667),
.B2(n_1666),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_SL g1735 ( 
.A(n_1698),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1704),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_L g1737 ( 
.A(n_1715),
.B(n_1536),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1699),
.A2(n_1667),
.B1(n_1666),
.B2(n_1672),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1694),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1704),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1703),
.A2(n_1667),
.B1(n_1652),
.B2(n_1518),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1667),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1723),
.A2(n_1697),
.B1(n_1694),
.B2(n_1690),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1735),
.Y(n_1744)
);

NOR4xp25_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1716),
.C(n_1697),
.D(n_1641),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1742),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1730),
.A2(n_1711),
.B1(n_1708),
.B2(n_1689),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1717),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1719),
.A2(n_1689),
.B1(n_1693),
.B2(n_1711),
.Y(n_1749)
);

AOI321xp33_ASAP7_75t_L g1750 ( 
.A1(n_1719),
.A2(n_1693),
.A3(n_1714),
.B1(n_1686),
.B2(n_1683),
.C(n_1692),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1718),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1724),
.Y(n_1752)
);

AOI322xp5_ASAP7_75t_L g1753 ( 
.A1(n_1726),
.A2(n_1627),
.A3(n_1652),
.B1(n_1615),
.B2(n_1612),
.C1(n_1640),
.C2(n_1641),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1727),
.A2(n_1686),
.B(n_1683),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_SL g1755 ( 
.A(n_1727),
.B(n_1692),
.C(n_1688),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1729),
.Y(n_1756)
);

AOI222xp33_ASAP7_75t_L g1757 ( 
.A1(n_1733),
.A2(n_1640),
.B1(n_1716),
.B2(n_1562),
.C1(n_1680),
.C2(n_1627),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1739),
.B(n_1663),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1728),
.B(n_1663),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1731),
.Y(n_1760)
);

AOI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1720),
.A2(n_1688),
.B(n_1714),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1732),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1748),
.Y(n_1763)
);

AOI222xp33_ASAP7_75t_L g1764 ( 
.A1(n_1744),
.A2(n_1740),
.B1(n_1736),
.B2(n_1721),
.C1(n_1734),
.C2(n_1737),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1744),
.B(n_1755),
.C(n_1761),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1758),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1751),
.Y(n_1767)
);

OAI211xp5_ASAP7_75t_L g1768 ( 
.A1(n_1750),
.A2(n_1722),
.B(n_1741),
.C(n_1725),
.Y(n_1768)
);

OA22x2_ASAP7_75t_L g1769 ( 
.A1(n_1749),
.A2(n_1742),
.B1(n_1664),
.B2(n_1677),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1746),
.B(n_1738),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1745),
.A2(n_1516),
.B(n_1518),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1758),
.B(n_1700),
.Y(n_1772)
);

XNOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1759),
.B(n_1518),
.Y(n_1773)
);

XNOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1743),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1752),
.Y(n_1775)
);

NAND4xp25_ASAP7_75t_L g1776 ( 
.A(n_1765),
.B(n_1757),
.C(n_1754),
.D(n_1755),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1766),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1770),
.B(n_1756),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1764),
.Y(n_1779)
);

NAND4xp25_ASAP7_75t_L g1780 ( 
.A(n_1764),
.B(n_1762),
.C(n_1760),
.D(n_1753),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1773),
.B(n_1569),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1768),
.B(n_1700),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1772),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1771),
.B(n_1705),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1769),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1774),
.B(n_1540),
.Y(n_1786)
);

O2A1O1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1779),
.A2(n_1771),
.B(n_1767),
.C(n_1763),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1776),
.B(n_1775),
.C(n_1710),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1780),
.A2(n_1710),
.B1(n_1705),
.B2(n_1671),
.C(n_1661),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1782),
.A2(n_1533),
.B1(n_1535),
.B2(n_1675),
.C(n_1680),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1785),
.A2(n_1671),
.B1(n_1664),
.B2(n_1495),
.C(n_1627),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1786),
.B1(n_1781),
.B2(n_1783),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1788),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1787),
.A2(n_1778),
.B1(n_1777),
.B2(n_1784),
.C(n_1468),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1790),
.A2(n_1671),
.B1(n_1547),
.B2(n_1627),
.C(n_1617),
.Y(n_1795)
);

AOI222xp33_ASAP7_75t_L g1796 ( 
.A1(n_1789),
.A2(n_1574),
.B1(n_1562),
.B2(n_1612),
.C1(n_1615),
.C2(n_1617),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1788),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1793),
.B1(n_1794),
.B2(n_1795),
.Y(n_1798)
);

NAND4xp75_ASAP7_75t_L g1799 ( 
.A(n_1792),
.B(n_1494),
.C(n_1497),
.D(n_1512),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1796),
.B(n_1675),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1793),
.A2(n_1468),
.B1(n_1602),
.B2(n_1589),
.Y(n_1801)
);

INVx5_ASAP7_75t_L g1802 ( 
.A(n_1793),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1798),
.A2(n_1801),
.B1(n_1802),
.B2(n_1799),
.C(n_1800),
.Y(n_1803)
);

NAND3x1_ASAP7_75t_L g1804 ( 
.A(n_1801),
.B(n_1468),
.C(n_1614),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1798),
.A2(n_1499),
.B(n_1632),
.Y(n_1805)
);

NOR2x1p5_ASAP7_75t_L g1806 ( 
.A(n_1803),
.B(n_1496),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1804),
.B1(n_1805),
.B2(n_1634),
.Y(n_1807)
);

AO22x2_ASAP7_75t_SL g1808 ( 
.A1(n_1807),
.A2(n_1496),
.B1(n_1616),
.B2(n_1629),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1634),
.B1(n_1613),
.B2(n_1629),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1808),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1809),
.Y(n_1811)
);

INVxp33_ASAP7_75t_L g1812 ( 
.A(n_1811),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1810),
.B(n_1613),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1812),
.A2(n_1617),
.B(n_1616),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1813),
.B(n_1499),
.Y(n_1815)
);

AO21x2_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1617),
.B(n_1616),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1630),
.B1(n_1625),
.B2(n_1607),
.C(n_1605),
.Y(n_1817)
);

AOI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1817),
.A2(n_1494),
.B(n_1493),
.C(n_1459),
.Y(n_1818)
);


endmodule