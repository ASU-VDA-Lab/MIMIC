module fake_jpeg_13215_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_27),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_1),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_67),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_76),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_62),
.Y(n_111)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_110),
.Y(n_125)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_58),
.B(n_77),
.C(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_118),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_74),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_1),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_53),
.B1(n_60),
.B2(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_65),
.B1(n_71),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_53),
.B1(n_60),
.B2(n_72),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_31),
.B1(n_47),
.B2(n_46),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_129),
.Y(n_153)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_139),
.B1(n_32),
.B2(n_45),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_69),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_59),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_73),
.B1(n_57),
.B2(n_52),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_56),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_3),
.B(n_4),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_2),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_2),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_149),
.Y(n_174)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_158),
.Y(n_169)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_161),
.B1(n_127),
.B2(n_130),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_4),
.B(n_5),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_162),
.B(n_142),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_5),
.C(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_29),
.B1(n_43),
.B2(n_11),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_7),
.B(n_10),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_12),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_133),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_13),
.C(n_14),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_157),
.B1(n_155),
.B2(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_167),
.C(n_160),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_170),
.B1(n_174),
.B2(n_169),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.C(n_184),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_173),
.C(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_176),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_180),
.B(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_149),
.B1(n_150),
.B2(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_152),
.B1(n_17),
.B2(n_24),
.C(n_33),
.Y(n_191)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_15),
.CON(n_192),
.SN(n_192)
);


endmodule