module fake_jpeg_1574_n_210 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_76),
.Y(n_80)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_48),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_63),
.B1(n_62),
.B2(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_91),
.B1(n_78),
.B2(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_53),
.B1(n_56),
.B2(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_63),
.B1(n_62),
.B2(n_61),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_91),
.B1(n_78),
.B2(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_97),
.B1(n_106),
.B2(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_102),
.Y(n_115)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_74),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_84),
.Y(n_122)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_1),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_74),
.B1(n_68),
.B2(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_118),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_88),
.C(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_57),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_67),
.B(n_65),
.C(n_56),
.D(n_60),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_107),
.B(n_77),
.Y(n_136)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

INVxp33_ASAP7_75t_SL g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_130),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_89),
.C(n_49),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_0),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_97),
.B1(n_107),
.B2(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_143),
.B1(n_147),
.B2(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_38),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_100),
.B(n_92),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_101),
.B(n_52),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_45),
.B(n_44),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_47),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_50),
.B1(n_49),
.B2(n_52),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_50),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_128),
.B1(n_120),
.B2(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_46),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_158),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_116),
.B1(n_123),
.B2(n_112),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_159),
.B1(n_163),
.B2(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_137),
.B1(n_151),
.B2(n_136),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_119),
.B1(n_8),
.B2(n_9),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_161),
.B(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_171),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_14),
.CI(n_15),
.CON(n_167),
.SN(n_167)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_140),
.A3(n_18),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_145),
.C(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_146),
.C(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_173),
.C(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_132),
.C(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_160),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_17),
.A3(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_182),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_31),
.B(n_35),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_28),
.C(n_32),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OAI322xp33_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_189),
.A3(n_174),
.B1(n_176),
.B2(n_180),
.C1(n_184),
.C2(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_156),
.B1(n_162),
.B2(n_153),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_155),
.B1(n_164),
.B2(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_181),
.C(n_168),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_198),
.C(n_37),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_196),
.A2(n_192),
.B1(n_193),
.B2(n_188),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_167),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_34),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_202),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_201),
.A2(n_198),
.B1(n_197),
.B2(n_199),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_202),
.C(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_23),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_23),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_24),
.C(n_25),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_24),
.Y(n_210)
);


endmodule