module fake_jpeg_29283_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_47),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_63),
.B1(n_70),
.B2(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_59),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_37),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_37),
.B(n_35),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_73),
.Y(n_85)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_29),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_89),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_35),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_35),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_119),
.B1(n_116),
.B2(n_110),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_19),
.B1(n_25),
.B2(n_27),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_19),
.B(n_25),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_80),
.B(n_67),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_22),
.C(n_33),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_112),
.C(n_115),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_19),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_118),
.B1(n_64),
.B2(n_52),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_21),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_61),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_34),
.B1(n_33),
.B2(n_26),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_27),
.B1(n_25),
.B2(n_34),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_82),
.C(n_77),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_143),
.C(n_150),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_66),
.B(n_23),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_108),
.B(n_117),
.C(n_32),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_52),
.B(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_133),
.B(n_136),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_64),
.B1(n_53),
.B2(n_72),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_131),
.B1(n_144),
.B2(n_146),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_135),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_53),
.B1(n_64),
.B2(n_33),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_120),
.B1(n_87),
.B2(n_97),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_100),
.B1(n_96),
.B2(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_71),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_147),
.B1(n_95),
.B2(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_91),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_71),
.C(n_84),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_65),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_93),
.A2(n_113),
.B1(n_107),
.B2(n_106),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_6),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_71),
.C(n_84),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_164),
.B1(n_171),
.B2(n_174),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_111),
.B1(n_98),
.B2(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_92),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_97),
.B1(n_87),
.B2(n_105),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_105),
.B1(n_65),
.B2(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_181),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_71),
.B1(n_90),
.B2(n_32),
.Y(n_168)
);

CKINVDCx10_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_2),
.C(n_5),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_173),
.B(n_133),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_21),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_21),
.B1(n_7),
.B2(n_9),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_6),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_21),
.C(n_7),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_125),
.C(n_130),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_16),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_132),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_169),
.B(n_176),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_207),
.B(n_179),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_137),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_122),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_201),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_122),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_135),
.Y(n_205)
);

HB1xp67_ASAP7_75t_SL g213 ( 
.A(n_205),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_134),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_178),
.C(n_163),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_160),
.B(n_156),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_209),
.A2(n_211),
.B(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_190),
.B1(n_159),
.B2(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_176),
.C(n_172),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_159),
.C(n_136),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_136),
.B(n_162),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_136),
.C(n_153),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_226),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_136),
.B1(n_138),
.B2(n_144),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_189),
.C(n_184),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_227),
.B(n_194),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_187),
.B1(n_195),
.B2(n_192),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_233),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_211),
.B(n_216),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_217),
.B(n_208),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_194),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_239),
.Y(n_249)
);

XNOR2x2_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_188),
.Y(n_233)
);

NOR4xp25_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_207),
.C(n_192),
.D(n_196),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_203),
.C(n_193),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_225),
.C(n_215),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_257),
.C(n_183),
.Y(n_267)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_212),
.B1(n_223),
.B2(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_255),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_242),
.B(n_237),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_240),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_258),
.B1(n_231),
.B2(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_232),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_214),
.C(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_183),
.B1(n_221),
.B2(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_267),
.C(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_239),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_268),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_272),
.A2(n_275),
.B1(n_247),
.B2(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_253),
.A3(n_250),
.B1(n_262),
.B2(n_268),
.C(n_251),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_281),
.B1(n_272),
.B2(n_276),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_260),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_R g279 ( 
.A(n_274),
.B(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_265),
.Y(n_282)
);

OAI321xp33_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_254),
.A3(n_256),
.B1(n_267),
.B2(n_263),
.C(n_249),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_284),
.B(n_132),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_270),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_287),
.B(n_9),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_182),
.B1(n_141),
.B2(n_11),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_288),
.B(n_11),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_288),
.B(n_11),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_10),
.Y(n_293)
);


endmodule