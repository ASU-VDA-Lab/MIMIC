module real_jpeg_24982_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_24),
.C(n_25),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_31),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_25),
.B1(n_40),
.B2(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_4),
.A2(n_7),
.B1(n_40),
.B2(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_4),
.B(n_63),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_49),
.C(n_52),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_4),
.B(n_31),
.C(n_77),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_4),
.B(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_54),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_25),
.B1(n_34),
.B2(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_22),
.B1(n_34),
.B2(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_79)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_31),
.B1(n_35),
.B2(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_31),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_11),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_121),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_119),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_97),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_97),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.C(n_85),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_16),
.A2(n_17),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_18),
.B(n_43),
.C(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_19),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_21),
.A2(n_22),
.B1(n_24),
.B2(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_62),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_25),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_25),
.B(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_27),
.A2(n_28),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_28),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_28),
.B(n_168),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_116),
.C(n_176),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_30),
.A2(n_37),
.B1(n_69),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_30),
.B(n_32),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_31),
.A2(n_35),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_31),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_32),
.A2(n_69),
.B(n_71),
.Y(n_68)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_32),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_33),
.A2(n_72),
.B(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_38),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_56),
.B2(n_66),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_42),
.A2(n_43),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_43),
.B(n_131),
.C(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_51),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_47),
.B(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_47),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OA22x2_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_53),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_52),
.B(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_67),
.A2(n_85),
.B1(n_86),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_74),
.B2(n_84),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_73),
.A2(n_74),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_73),
.A2(n_74),
.B1(n_94),
.B2(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_95),
.C(n_183),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B(n_80),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_94),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_88),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_87),
.A2(n_88),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_118),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_116),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_116),
.B1(n_135),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_126),
.C(n_135),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_199),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_193),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_152),
.B(n_192),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_142),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_125),
.B(n_142),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_127),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_150),
.C(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_185),
.B(n_191),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_179),
.B(n_184),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_171),
.B(n_178),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_161),
.B(n_170),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_167),
.B(n_169),
.Y(n_161)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);


endmodule