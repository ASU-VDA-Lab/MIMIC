module real_aes_17424_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_660, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_660;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_0), .A2(n_28), .B1(n_115), .B2(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_1), .B(n_498), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_2), .A2(n_7), .B1(n_108), .B2(n_179), .Y(n_178) );
INVx1_ASAP7_75t_SL g650 ( .A(n_2), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_3), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_4), .A2(n_9), .B1(n_89), .B2(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_4), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_4), .Y(n_632) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_6), .Y(n_183) );
INVx1_ASAP7_75t_L g469 ( .A(n_8), .Y(n_469) );
INVx1_ASAP7_75t_L g444 ( .A(n_10), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_10), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_11), .A2(n_75), .B1(n_108), .B2(n_110), .Y(n_107) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_12), .A2(n_49), .B1(n_525), .B2(n_528), .Y(n_524) );
INVx1_ASAP7_75t_L g564 ( .A(n_12), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_13), .A2(n_25), .B1(n_140), .B2(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g437 ( .A(n_14), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_15), .B(n_109), .Y(n_137) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_16), .A2(n_38), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g465 ( .A(n_17), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_18), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_19), .A2(n_32), .B1(n_153), .B2(n_154), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_20), .A2(n_36), .B1(n_108), .B2(n_154), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_21), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_22), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_23), .Y(n_213) );
INVx1_ASAP7_75t_L g470 ( .A(n_24), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_26), .A2(n_63), .B1(n_115), .B2(n_189), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_27), .A2(n_31), .B1(n_115), .B2(n_136), .Y(n_165) );
XOR2xp5_ASAP7_75t_L g426 ( .A(n_29), .B(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_30), .A2(n_39), .B1(n_108), .B2(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g436 ( .A(n_33), .Y(n_436) );
INVx1_ASAP7_75t_L g475 ( .A(n_33), .Y(n_475) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_34), .Y(n_633) );
INVx2_ASAP7_75t_L g620 ( .A(n_35), .Y(n_620) );
INVx1_ASAP7_75t_L g479 ( .A(n_37), .Y(n_479) );
BUFx2_ASAP7_75t_L g643 ( .A(n_40), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_41), .A2(n_72), .B1(n_485), .B2(n_494), .Y(n_484) );
INVx1_ASAP7_75t_L g559 ( .A(n_41), .Y(n_559) );
OA211x2_ASAP7_75t_L g502 ( .A1(n_42), .A2(n_503), .B(n_507), .C(n_513), .Y(n_502) );
INVx1_ASAP7_75t_L g547 ( .A(n_42), .Y(n_547) );
BUFx3_ASAP7_75t_L g442 ( .A(n_43), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_44), .A2(n_56), .B1(n_114), .B2(n_153), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_45), .A2(n_57), .B1(n_115), .B2(n_136), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_46), .A2(n_74), .B1(n_108), .B2(n_164), .Y(n_210) );
AND2x4_ASAP7_75t_L g82 ( .A(n_47), .B(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_47), .Y(n_606) );
INVx1_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g555 ( .A(n_49), .Y(n_555) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_50), .Y(n_491) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
INVx1_ASAP7_75t_L g453 ( .A(n_52), .Y(n_453) );
INVx1_ASAP7_75t_L g460 ( .A(n_53), .Y(n_460) );
INVx1_ASAP7_75t_L g445 ( .A(n_54), .Y(n_445) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_55), .Y(n_490) );
INVx2_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_59), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_60), .A2(n_73), .B1(n_154), .B2(n_192), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_61), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_62), .Y(n_157) );
INVx1_ASAP7_75t_L g493 ( .A(n_64), .Y(n_493) );
BUFx3_ASAP7_75t_L g498 ( .A(n_64), .Y(n_498) );
INVx1_ASAP7_75t_SL g641 ( .A(n_65), .Y(n_641) );
INVx1_ASAP7_75t_L g514 ( .A(n_66), .Y(n_514) );
INVx1_ASAP7_75t_L g481 ( .A(n_67), .Y(n_481) );
INVx1_ASAP7_75t_L g434 ( .A(n_68), .Y(n_434) );
INVx2_ASAP7_75t_L g473 ( .A(n_68), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_69), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_70), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_71), .B(n_109), .Y(n_142) );
INVx1_ASAP7_75t_L g567 ( .A(n_72), .Y(n_567) );
INVx1_ASAP7_75t_L g517 ( .A(n_76), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_425), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_84), .Y(n_80) );
INVx2_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
AO31x2_ASAP7_75t_L g148 ( .A1(n_81), .A2(n_149), .A3(n_155), .B(n_156), .Y(n_148) );
AO31x2_ASAP7_75t_L g161 ( .A1(n_81), .A2(n_162), .A3(n_168), .B(n_170), .Y(n_161) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_81), .A2(n_174), .A3(n_181), .B(n_182), .Y(n_173) );
BUFx10_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_83), .Y(n_608) );
INVxp67_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AO21x1_ASAP7_75t_L g657 ( .A1(n_85), .A2(n_607), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_88), .Y(n_85) );
INVx6_ASAP7_75t_L g112 ( .A(n_86), .Y(n_112) );
O2A1O1Ixp5_ASAP7_75t_L g134 ( .A1(n_86), .A2(n_135), .B(n_136), .C(n_137), .Y(n_134) );
BUFx8_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
INVx1_ASAP7_75t_L g167 ( .A(n_87), .Y(n_167) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_92), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
INVx3_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
INVx1_ASAP7_75t_L g177 ( .A(n_92), .Y(n_177) );
INVx1_ASAP7_75t_L g180 ( .A(n_92), .Y(n_180) );
INVx2_ASAP7_75t_L g190 ( .A(n_92), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_92), .Y(n_192) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
OR2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_328), .Y(n_95) );
NAND4xp25_ASAP7_75t_L g96 ( .A(n_97), .B(n_252), .C(n_283), .D(n_312), .Y(n_96) );
NOR2xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_219), .Y(n_97) );
OAI322xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_158), .A3(n_184), .B1(n_197), .B2(n_205), .C1(n_214), .C2(n_216), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_100), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_128), .Y(n_100) );
AND2x2_ASAP7_75t_L g249 ( .A(n_101), .B(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g285 ( .A(n_101), .Y(n_285) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g260 ( .A(n_102), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g263 ( .A(n_102), .B(n_160), .Y(n_263) );
AND2x2_ASAP7_75t_L g280 ( .A(n_102), .B(n_173), .Y(n_280) );
AND2x2_ASAP7_75t_L g378 ( .A(n_102), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g201 ( .A(n_103), .Y(n_201) );
AND2x4_ASAP7_75t_L g384 ( .A(n_103), .B(n_379), .Y(n_384) );
AO31x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_106), .A3(n_119), .B(n_125), .Y(n_103) );
AO31x2_ASAP7_75t_L g208 ( .A1(n_104), .A2(n_168), .A3(n_209), .B(n_212), .Y(n_208) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B1(n_113), .B2(n_116), .Y(n_106) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_112), .A2(n_139), .B(n_142), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_112), .A2(n_116), .B1(n_150), .B2(n_152), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_112), .A2(n_163), .B1(n_165), .B2(n_166), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_112), .A2(n_116), .B1(n_175), .B2(n_178), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_112), .A2(n_188), .B1(n_191), .B2(n_193), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_112), .A2(n_166), .B1(n_210), .B2(n_211), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_112), .A2(n_116), .B1(n_229), .B2(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx4_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
INVx1_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_119), .A2(n_194), .A3(n_228), .B(n_231), .Y(n_227) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_121), .B(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_121), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g127 ( .A(n_122), .Y(n_127) );
INVx2_ASAP7_75t_L g169 ( .A(n_122), .Y(n_169) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_123), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_127), .B(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g389 ( .A(n_128), .B(n_290), .Y(n_389) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g218 ( .A(n_129), .Y(n_218) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_129), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_147), .Y(n_129) );
AND2x2_ASAP7_75t_L g206 ( .A(n_130), .B(n_148), .Y(n_206) );
INVx1_ASAP7_75t_L g247 ( .A(n_130), .Y(n_247) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_145), .Y(n_130) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_131), .A2(n_133), .B(n_145), .Y(n_242) );
INVx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_132), .B(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_132), .B(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_132), .B(n_213), .Y(n_212) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_138), .B(n_143), .Y(n_133) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_SL g194 ( .A(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
INVx2_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
AND2x2_ASAP7_75t_L g302 ( .A(n_147), .B(n_241), .Y(n_302) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g256 ( .A(n_148), .Y(n_256) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_148), .Y(n_309) );
OR2x2_ASAP7_75t_L g380 ( .A(n_148), .B(n_186), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_158), .B(n_259), .C(n_262), .D(n_264), .Y(n_258) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g396 ( .A(n_159), .B(n_384), .Y(n_396) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_160), .B(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g250 ( .A(n_160), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g270 ( .A(n_160), .Y(n_270) );
INVx1_ASAP7_75t_L g287 ( .A(n_160), .Y(n_287) );
INVx1_ASAP7_75t_L g295 ( .A(n_160), .Y(n_295) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_160), .Y(n_409) );
INVx4_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_161), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g327 ( .A(n_161), .B(n_227), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_161), .B(n_173), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_161), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g400 ( .A(n_161), .Y(n_400) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g204 ( .A(n_173), .Y(n_204) );
OR2x2_ASAP7_75t_L g265 ( .A(n_173), .B(n_227), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_173), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_173), .B(n_225), .Y(n_296) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_173), .Y(n_383) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_181), .A2(n_187), .A3(n_194), .B(n_195), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_184), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g207 ( .A(n_186), .B(n_208), .Y(n_207) );
BUFx2_ASAP7_75t_L g217 ( .A(n_186), .Y(n_217) );
INVx2_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
AND2x4_ASAP7_75t_L g267 ( .A(n_186), .B(n_239), .Y(n_267) );
OR2x2_ASAP7_75t_L g347 ( .A(n_186), .B(n_247), .Y(n_347) );
INVx2_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_199), .B(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g264 ( .A(n_199), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_199), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_200), .B(n_270), .Y(n_278) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
OR2x2_ASAP7_75t_L g316 ( .A(n_201), .B(n_226), .Y(n_316) );
INVx1_ASAP7_75t_L g243 ( .A(n_202), .Y(n_243) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g215 ( .A(n_203), .Y(n_215) );
INVx1_ASAP7_75t_L g251 ( .A(n_204), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
OAI322xp33_ASAP7_75t_L g219 ( .A1(n_206), .A2(n_220), .A3(n_233), .B1(n_236), .B2(n_243), .C1(n_244), .C2(n_248), .Y(n_219) );
AND2x4_ASAP7_75t_L g266 ( .A(n_206), .B(n_267), .Y(n_266) );
AOI211xp5_ASAP7_75t_SL g297 ( .A1(n_206), .A2(n_298), .B(n_299), .C(n_303), .Y(n_297) );
AND2x2_ASAP7_75t_L g317 ( .A(n_206), .B(n_207), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_206), .B(n_234), .Y(n_323) );
AND2x4_ASAP7_75t_SL g245 ( .A(n_207), .B(n_246), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_207), .B(n_263), .C(n_291), .Y(n_336) );
AND2x2_ASAP7_75t_L g367 ( .A(n_207), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g234 ( .A(n_208), .B(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g239 ( .A(n_208), .Y(n_239) );
BUFx2_ASAP7_75t_L g307 ( .A(n_208), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_217), .B(n_241), .Y(n_240) );
NAND2x1_ASAP7_75t_L g281 ( .A(n_217), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g300 ( .A(n_217), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_218), .B(n_234), .Y(n_365) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_224), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g308 ( .A(n_223), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_227), .Y(n_261) );
AND2x4_ASAP7_75t_L g271 ( .A(n_227), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g358 ( .A(n_227), .Y(n_358) );
INVx2_ASAP7_75t_L g379 ( .A(n_227), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_233), .A2(n_392), .B1(n_394), .B2(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g303 ( .A(n_234), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g257 ( .A(n_235), .B(n_241), .Y(n_257) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g276 ( .A(n_237), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x4_ASAP7_75t_L g246 ( .A(n_238), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g368 ( .A(n_238), .Y(n_368) );
INVx2_ASAP7_75t_L g254 ( .A(n_239), .Y(n_254) );
AND2x2_ASAP7_75t_L g282 ( .A(n_239), .B(n_241), .Y(n_282) );
INVx3_ASAP7_75t_L g290 ( .A(n_239), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_239), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g275 ( .A(n_240), .Y(n_275) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g291 ( .A(n_242), .Y(n_291) );
OAI222xp33_ASAP7_75t_L g414 ( .A1(n_244), .A2(n_404), .B1(n_415), .B2(n_418), .C1(n_420), .C2(n_422), .Y(n_414) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g355 ( .A(n_246), .Y(n_355) );
AND2x2_ASAP7_75t_L g419 ( .A(n_246), .B(n_289), .Y(n_419) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_249), .B(n_340), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .B1(n_266), .B2(n_268), .C(n_273), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g341 ( .A(n_254), .Y(n_341) );
INVx2_ASAP7_75t_L g403 ( .A(n_255), .Y(n_403) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g304 ( .A(n_256), .Y(n_304) );
AND2x2_ASAP7_75t_L g340 ( .A(n_256), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g306 ( .A(n_257), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g421 ( .A(n_257), .Y(n_421) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g370 ( .A(n_261), .Y(n_370) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g393 ( .A(n_263), .B(n_271), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_263), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g277 ( .A(n_265), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g412 ( .A(n_265), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_266), .A2(n_320), .B1(n_354), .B2(n_356), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_266), .A2(n_382), .B(n_385), .Y(n_381) );
INVxp67_ASAP7_75t_L g298 ( .A(n_267), .Y(n_298) );
INVx2_ASAP7_75t_SL g402 ( .A(n_267), .Y(n_402) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g315 ( .A(n_269), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g413 ( .A(n_269), .B(n_412), .Y(n_413) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g286 ( .A(n_271), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_271), .B(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g338 ( .A(n_271), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B1(n_279), .B2(n_281), .Y(n_273) );
NOR2xp33_ASAP7_75t_SL g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_275), .A2(n_349), .B1(n_362), .B2(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g371 ( .A(n_280), .B(n_372), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B(n_292), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g352 ( .A(n_285), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_285), .B(n_335), .Y(n_363) );
INVx1_ASAP7_75t_L g321 ( .A(n_287), .Y(n_321) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_289), .B(n_302), .Y(n_394) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_290), .A2(n_408), .B(n_410), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_297), .B(n_305), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
INVx1_ASAP7_75t_L g417 ( .A(n_296), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g390 ( .A(n_300), .Y(n_390) );
OR2x2_ASAP7_75t_L g401 ( .A(n_301), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .C(n_310), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_306), .A2(n_367), .B1(n_369), .B2(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_308), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_311), .B(n_315), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_311), .A2(n_374), .B1(n_377), .B2(n_380), .C(n_381), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .B(n_318), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g322 ( .A(n_316), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B1(n_324), .B2(n_660), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g405 ( .A(n_327), .B(n_383), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_329), .B(n_359), .C(n_386), .D(n_406), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_342), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_336), .B2(n_337), .C(n_339), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_332), .A2(n_389), .B1(n_411), .B2(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g385 ( .A(n_334), .Y(n_385) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g369 ( .A(n_335), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_335), .B(n_378), .Y(n_377) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_335), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_337), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_341), .B(n_345), .Y(n_344) );
OAI21xp33_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_348), .B(n_353), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_358), .A2(n_387), .B(n_391), .C(n_397), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_373), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_366), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g420 ( .A(n_368), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx3_ASAP7_75t_L g424 ( .A(n_384), .Y(n_424) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp33_ASAP7_75t_R g397 ( .A1(n_398), .A2(n_401), .B1(n_403), .B2(n_404), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g411 ( .A(n_400), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_414), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_602), .B1(n_609), .B2(n_651), .C(n_652), .Y(n_425) );
INVx1_ASAP7_75t_L g651 ( .A(n_427), .Y(n_651) );
INVxp33_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR4xp25_ASAP7_75t_L g428 ( .A(n_429), .B(n_482), .C(n_539), .D(n_576), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_438), .A3(n_454), .B1(n_466), .B2(n_471), .B3(n_477), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_432), .Y(n_575) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_432), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g538 ( .A(n_433), .Y(n_538) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g625 ( .A(n_435), .Y(n_625) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_437), .Y(n_435) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_436), .Y(n_573) );
INVx1_ASAP7_75t_L g619 ( .A(n_436), .Y(n_619) );
INVx3_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
BUFx3_ASAP7_75t_L g545 ( .A(n_437), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_445), .B1(n_446), .B2(n_453), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g478 ( .A(n_441), .Y(n_478) );
OR2x4_ASAP7_75t_L g566 ( .A(n_441), .B(n_476), .Y(n_566) );
OR2x4_ASAP7_75t_L g569 ( .A(n_441), .B(n_557), .Y(n_569) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_442), .Y(n_452) );
INVx2_ASAP7_75t_L g459 ( .A(n_442), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_442), .B(n_451), .Y(n_464) );
AND2x4_ASAP7_75t_L g551 ( .A(n_442), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g458 ( .A(n_444), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_445), .A2(n_479), .B1(n_583), .B2(n_584), .Y(n_582) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_448), .Y(n_480) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
BUFx2_ASAP7_75t_L g549 ( .A(n_450), .Y(n_549) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g552 ( .A(n_451), .Y(n_552) );
BUFx2_ASAP7_75t_L g546 ( .A(n_452), .Y(n_546) );
INVx2_ASAP7_75t_L g617 ( .A(n_452), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_453), .A2(n_481), .B1(n_589), .B2(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_460), .B1(n_461), .B2(n_465), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx8_ASAP7_75t_L g468 ( .A(n_457), .Y(n_468) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_457), .Y(n_558) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g585 ( .A1(n_460), .A2(n_469), .B1(n_586), .B2(n_589), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_461), .A2(n_467), .B1(n_469), .B2(n_470), .Y(n_466) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g562 ( .A(n_464), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_465), .A2(n_470), .B1(n_583), .B2(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
AND2x4_ASAP7_75t_L g580 ( .A(n_472), .B(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x4_ASAP7_75t_L g553 ( .A(n_476), .B(n_551), .Y(n_553) );
INVx1_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
OR2x6_ASAP7_75t_L g561 ( .A(n_476), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g618 ( .A(n_476), .B(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_480), .B2(n_481), .Y(n_477) );
AOI31xp67_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_502), .A3(n_523), .B(n_532), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_492), .Y(n_486) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_487), .Y(n_583) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g527 ( .A(n_488), .Y(n_527) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g501 ( .A(n_490), .Y(n_501) );
NAND2x1_ASAP7_75t_L g506 ( .A(n_490), .B(n_491), .Y(n_506) );
AND2x2_ASAP7_75t_L g512 ( .A(n_490), .B(n_491), .Y(n_512) );
INVx1_ASAP7_75t_L g522 ( .A(n_490), .Y(n_522) );
AND2x2_ASAP7_75t_L g530 ( .A(n_490), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g588 ( .A(n_490), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_491), .B(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g516 ( .A(n_491), .Y(n_516) );
INVx2_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
OR2x2_ASAP7_75t_L g587 ( .A(n_491), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g529 ( .A(n_492), .B(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
AND2x4_ASAP7_75t_L g515 ( .A(n_497), .B(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g510 ( .A(n_498), .Y(n_510) );
AND2x4_ASAP7_75t_L g520 ( .A(n_498), .B(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g598 ( .A(n_498), .B(n_536), .Y(n_598) );
BUFx2_ASAP7_75t_L g584 ( .A(n_499), .Y(n_584) );
INVx8_ASAP7_75t_L g601 ( .A(n_499), .Y(n_601) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx5_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_506), .Y(n_591) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_L g526 ( .A(n_510), .Y(n_526) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_514), .A2(n_517), .B1(n_543), .B2(n_547), .C1(n_548), .C2(n_550), .Y(n_542) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI31xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_554), .A3(n_563), .B(n_570), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x4_ASAP7_75t_L g548 ( .A(n_544), .B(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B1(n_559), .B2(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_567), .B2(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
CKINVDCx14_ASAP7_75t_R g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI33xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_582), .A3(n_585), .B1(n_592), .B2(n_596), .B3(n_599), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx4_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g595 ( .A(n_587), .Y(n_595) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx4_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g627 ( .A(n_606), .Y(n_627) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_608), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g658 ( .A(n_608), .B(n_627), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_628), .B1(n_644), .B2(n_649), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx12f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx4f_ASAP7_75t_SL g654 ( .A(n_612), .Y(n_654) );
BUFx8_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_620), .B(n_621), .C(n_626), .Y(n_613) );
AND2x2_ASAP7_75t_L g648 ( .A(n_614), .B(n_621), .Y(n_648) );
INVx4_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x6_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_616), .B(n_622), .C(n_625), .Y(n_621) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g647 ( .A(n_626), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_628), .A2(n_649), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_638), .B2(n_639), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_630) );
INVx1_ASAP7_75t_L g637 ( .A(n_631), .Y(n_637) );
INVx1_ASAP7_75t_L g634 ( .A(n_633), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_SL g656 ( .A(n_646), .Y(n_656) );
OR2x6_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_657), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
endmodule