module fake_jpeg_24371_n_257 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_50),
.B1(n_53),
.B2(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_21),
.B1(n_19),
.B2(n_29),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_23),
.B1(n_38),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_29),
.B1(n_20),
.B2(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_29),
.B1(n_20),
.B2(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_14),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_24),
.B1(n_20),
.B2(n_29),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_41),
.B1(n_48),
.B2(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_76),
.B1(n_49),
.B2(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_16),
.B1(n_18),
.B2(n_25),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_23),
.B(n_22),
.C(n_38),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_18),
.B1(n_15),
.B2(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_57),
.B1(n_54),
.B2(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2x1_ASAP7_75t_R g101 ( 
.A(n_74),
.B(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_36),
.B1(n_14),
.B2(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_15),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_48),
.B1(n_58),
.B2(n_43),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_88),
.B1(n_89),
.B2(n_64),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_96),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_100),
.B(n_101),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_55),
.B1(n_48),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_85),
.B1(n_80),
.B2(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_65),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_48),
.B(n_27),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_66),
.B(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_105),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_65),
.Y(n_106)
);

FAx1_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_118),
.CI(n_123),
.CON(n_125),
.SN(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_110),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_115),
.A3(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_68),
.B(n_60),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_120),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_41),
.B(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_78),
.B1(n_63),
.B2(n_77),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_61),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_87),
.B(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_86),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_23),
.B(n_56),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_91),
.B1(n_82),
.B2(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_135),
.B1(n_143),
.B2(n_122),
.Y(n_151)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_130),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_101),
.B(n_89),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_111),
.B(n_109),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_107),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_7),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_8),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_142),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_94),
.B1(n_78),
.B2(n_23),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_140),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_56),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_39),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_77),
.B1(n_73),
.B2(n_99),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_128),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_106),
.B1(n_121),
.B2(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_119),
.C(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_157),
.C(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_121),
.B1(n_103),
.B2(n_113),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_158),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_119),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_154),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_111),
.C(n_99),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_56),
.B1(n_45),
.B2(n_39),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_132),
.B1(n_144),
.B2(n_135),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_45),
.B1(n_23),
.B2(n_2),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_23),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_135),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_12),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_175),
.B1(n_135),
.B2(n_128),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_165),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_183),
.B(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_124),
.C(n_131),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_186),
.C(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_133),
.C(n_130),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_185),
.B(n_170),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_152),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_164),
.C(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_158),
.C(n_159),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_150),
.C(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_197),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_180),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_139),
.C(n_1),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_186),
.C(n_185),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_208),
.C(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_190),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_171),
.CI(n_176),
.CON(n_211),
.SN(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_216),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_179),
.B1(n_173),
.B2(n_177),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_215),
.B1(n_213),
.B2(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_181),
.C(n_175),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_214),
.C(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.C(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_139),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_0),
.C(n_1),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_0),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_9),
.B(n_12),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_11),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_210),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_220),
.B(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_235),
.C(n_233),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_248),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_9),
.B(n_13),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_239),
.B(n_240),
.C(n_9),
.D(n_13),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_3),
.C(n_4),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_3),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_247),
.B(n_250),
.C(n_4),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_5),
.Y(n_257)
);


endmodule