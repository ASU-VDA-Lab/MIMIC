module real_aes_6935_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_316;
wire n_284;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_252;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g496 ( .A1(n_0), .A2(n_160), .B(n_497), .C(n_500), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_1), .B(n_492), .Y(n_501) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g158 ( .A(n_3), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_4), .B(n_161), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_5), .A2(n_460), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_6), .A2(n_168), .B(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_7), .A2(n_35), .B1(n_148), .B2(n_196), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_8), .B(n_168), .Y(n_176) );
AND2x6_ASAP7_75t_L g163 ( .A(n_9), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_10), .A2(n_163), .B(n_465), .C(n_509), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_11), .A2(n_39), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_11), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_12), .B(n_36), .Y(n_117) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_15), .B(n_144), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_16), .B(n_161), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_17), .B(n_135), .Y(n_242) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_18), .A2(n_134), .A3(n_168), .B1(n_187), .B2(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_19), .B(n_148), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_20), .B(n_135), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_21), .A2(n_55), .B1(n_148), .B2(n_196), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g198 ( .A1(n_22), .A2(n_81), .B1(n_144), .B2(n_148), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_23), .B(n_148), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_24), .A2(n_187), .B(n_465), .C(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_25), .A2(n_187), .B(n_465), .C(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_26), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_27), .B(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_28), .A2(n_460), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_29), .B(n_189), .Y(n_230) );
INVx2_ASAP7_75t_L g146 ( .A(n_30), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_31), .A2(n_463), .B(n_467), .C(n_473), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_32), .B(n_148), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_33), .B(n_189), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_34), .B(n_207), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_37), .B(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_38), .Y(n_513) );
INVx1_ASAP7_75t_L g741 ( .A(n_39), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_40), .B(n_161), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_41), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_41), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_42), .B(n_460), .Y(n_516) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_43), .A2(n_122), .B1(n_123), .B2(n_444), .Y(n_121) );
INVx1_ASAP7_75t_L g444 ( .A(n_43), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_43), .A2(n_45), .B1(n_444), .B2(n_754), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_44), .A2(n_463), .B(n_473), .C(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_45), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_46), .B(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g498 ( .A(n_47), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_48), .A2(n_91), .B1(n_196), .B2(n_197), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_49), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_50), .B(n_148), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_51), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g529 ( .A(n_52), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_53), .B(n_460), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_54), .B(n_156), .Y(n_175) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_56), .A2(n_61), .B1(n_144), .B2(n_148), .Y(n_240) );
AOI222xp33_ASAP7_75t_L g118 ( .A1(n_57), .A2(n_119), .B1(n_738), .B2(n_739), .C1(n_742), .C2(n_745), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_58), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_59), .B(n_148), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_60), .B(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g164 ( .A(n_62), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_63), .B(n_460), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_64), .B(n_492), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_65), .A2(n_150), .B(n_156), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_66), .B(n_148), .Y(n_159) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_68), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_69), .B(n_161), .Y(n_471) );
AO32x2_ASAP7_75t_L g193 ( .A1(n_70), .A2(n_168), .A3(n_187), .B1(n_194), .B2(n_199), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_71), .B(n_162), .Y(n_510) );
INVx1_ASAP7_75t_L g183 ( .A(n_72), .Y(n_183) );
INVx1_ASAP7_75t_L g225 ( .A(n_73), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_74), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_75), .B(n_470), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_76), .A2(n_465), .B(n_473), .C(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_77), .B(n_144), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_78), .Y(n_537) );
INVx1_ASAP7_75t_L g761 ( .A(n_79), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_80), .B(n_469), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_82), .B(n_196), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g102 ( .A1(n_83), .A2(n_103), .B1(n_758), .B2(n_762), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_84), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_85), .B(n_144), .Y(n_229) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_87), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_88), .B(n_186), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_89), .B(n_144), .Y(n_172) );
OR2x2_ASAP7_75t_L g113 ( .A(n_90), .B(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g447 ( .A(n_90), .B(n_115), .Y(n_447) );
INVx2_ASAP7_75t_L g451 ( .A(n_90), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_92), .A2(n_101), .B1(n_144), .B2(n_145), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_93), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g468 ( .A(n_94), .Y(n_468) );
INVxp67_ASAP7_75t_L g540 ( .A(n_95), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_96), .B(n_144), .Y(n_181) );
INVx1_ASAP7_75t_L g506 ( .A(n_97), .Y(n_506) );
INVx1_ASAP7_75t_L g564 ( .A(n_98), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_99), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g531 ( .A(n_100), .B(n_189), .Y(n_531) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_118), .B1(n_747), .B2(n_749), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g748 ( .A(n_107), .Y(n_748) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_109), .A2(n_750), .B(n_757), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g757 ( .A(n_112), .Y(n_757) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_114), .B(n_451), .Y(n_744) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g450 ( .A(n_115), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OAI22x1_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_445), .B1(n_448), .B2(n_452), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_121), .A2(n_445), .B1(n_450), .B2(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_122), .A2(n_123), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_410), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_314), .C(n_398), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_257), .C(n_279), .D(n_295), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_190), .B1(n_216), .B2(n_235), .C(n_243), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_166), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_129), .B(n_235), .Y(n_269) );
NAND4xp25_ASAP7_75t_L g309 ( .A(n_129), .B(n_297), .C(n_310), .D(n_312), .Y(n_309) );
INVxp67_ASAP7_75t_L g426 ( .A(n_129), .Y(n_426) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g308 ( .A(n_130), .B(n_246), .Y(n_308) );
AND2x2_ASAP7_75t_L g332 ( .A(n_130), .B(n_166), .Y(n_332) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g299 ( .A(n_131), .B(n_234), .Y(n_299) );
AND2x2_ASAP7_75t_L g339 ( .A(n_131), .B(n_320), .Y(n_339) );
AND2x2_ASAP7_75t_L g356 ( .A(n_131), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_131), .B(n_167), .Y(n_380) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g233 ( .A(n_132), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g251 ( .A(n_132), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g263 ( .A(n_132), .B(n_167), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_132), .B(n_177), .Y(n_285) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_165), .Y(n_132) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_133), .A2(n_178), .B(n_188), .Y(n_177) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_134), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_136), .B(n_137), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_154), .B(n_163), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_147), .C(n_150), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_143), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_143), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx3_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_148), .Y(n_566) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g196 ( .A(n_149), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
AND2x6_ASAP7_75t_L g465 ( .A(n_149), .B(n_466), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_150), .A2(n_564), .B(n_565), .C(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_151), .A2(n_228), .B(n_229), .Y(n_227) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g470 ( .A(n_152), .Y(n_470) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx1_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
AND2x2_ASAP7_75t_L g461 ( .A(n_153), .B(n_157), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_153), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_159), .C(n_160), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_155), .A2(n_183), .B(n_184), .C(n_185), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_155), .A2(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_160), .A2(n_174), .B(n_175), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_186), .B1(n_214), .B2(n_215), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_160), .A2(n_186), .B1(n_239), .B2(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_161), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_161), .A2(n_180), .B(n_181), .Y(n_179) );
O2A1O1Ixp5_ASAP7_75t_SL g223 ( .A1(n_161), .A2(n_224), .B(n_225), .C(n_226), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_161), .B(n_540), .Y(n_539) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_162), .A2(n_186), .B1(n_195), .B2(n_198), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_163), .A2(n_170), .B(n_173), .Y(n_169) );
BUFx3_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_163), .A2(n_203), .B(n_208), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_163), .A2(n_223), .B(n_227), .Y(n_222) );
AND2x4_ASAP7_75t_L g460 ( .A(n_163), .B(n_461), .Y(n_460) );
INVx4_ASAP7_75t_SL g474 ( .A(n_163), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_163), .B(n_461), .Y(n_507) );
AND2x2_ASAP7_75t_L g266 ( .A(n_166), .B(n_267), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_166), .A2(n_316), .B1(n_319), .B2(n_321), .C(n_325), .Y(n_315) );
AND2x2_ASAP7_75t_L g374 ( .A(n_166), .B(n_339), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_166), .B(n_356), .Y(n_408) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_177), .Y(n_166) );
INVx3_ASAP7_75t_L g234 ( .A(n_167), .Y(n_234) );
AND2x2_ASAP7_75t_L g283 ( .A(n_167), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g337 ( .A(n_167), .B(n_252), .Y(n_337) );
AND2x2_ASAP7_75t_L g395 ( .A(n_167), .B(n_396), .Y(n_395) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_176), .Y(n_167) );
INVx4_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_168), .A2(n_516), .B(n_517), .Y(n_515) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_168), .Y(n_534) );
AND2x2_ASAP7_75t_L g235 ( .A(n_177), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g252 ( .A(n_177), .Y(n_252) );
INVx1_ASAP7_75t_L g307 ( .A(n_177), .Y(n_307) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_177), .Y(n_313) );
AND2x2_ASAP7_75t_L g358 ( .A(n_177), .B(n_234), .Y(n_358) );
OR2x2_ASAP7_75t_L g397 ( .A(n_177), .B(n_236), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_187), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_185), .A2(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx4_ASAP7_75t_L g499 ( .A(n_186), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_187), .B(n_237), .C(n_238), .Y(n_256) );
INVx2_ASAP7_75t_L g199 ( .A(n_189), .Y(n_199) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_189), .A2(n_202), .B(n_211), .Y(n_201) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_189), .A2(n_222), .B(n_230), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_189), .A2(n_459), .B(n_462), .Y(n_458) );
INVx1_ASAP7_75t_L g489 ( .A(n_189), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_189), .A2(n_526), .B(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_190), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
AND2x2_ASAP7_75t_L g393 ( .A(n_191), .B(n_390), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_191), .B(n_375), .Y(n_425) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g324 ( .A(n_192), .B(n_248), .Y(n_324) );
AND2x2_ASAP7_75t_L g373 ( .A(n_192), .B(n_219), .Y(n_373) );
INVx1_ASAP7_75t_L g419 ( .A(n_192), .Y(n_419) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
AND2x2_ASAP7_75t_L g274 ( .A(n_193), .B(n_248), .Y(n_274) );
INVx1_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_193), .B(n_212), .Y(n_297) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_197), .Y(n_472) );
INVx2_ASAP7_75t_L g500 ( .A(n_197), .Y(n_500) );
INVx1_ASAP7_75t_L g486 ( .A(n_199), .Y(n_486) );
AND2x2_ASAP7_75t_L g365 ( .A(n_200), .B(n_273), .Y(n_365) );
INVx2_ASAP7_75t_L g430 ( .A(n_200), .Y(n_430) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AND2x2_ASAP7_75t_L g247 ( .A(n_201), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g260 ( .A(n_201), .B(n_220), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_201), .B(n_219), .Y(n_288) );
INVx1_ASAP7_75t_L g294 ( .A(n_201), .Y(n_294) );
INVx1_ASAP7_75t_L g311 ( .A(n_201), .Y(n_311) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_201), .Y(n_323) );
INVx2_ASAP7_75t_L g391 ( .A(n_201), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g248 ( .A(n_212), .Y(n_248) );
BUFx2_ASAP7_75t_L g345 ( .A(n_212), .Y(n_345) );
AND2x2_ASAP7_75t_L g390 ( .A(n_212), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_218), .B(n_327), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_218), .A2(n_389), .B(n_403), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_218), .B(n_324), .Y(n_438) );
BUFx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g360 ( .A(n_220), .Y(n_360) );
AND2x2_ASAP7_75t_L g389 ( .A(n_220), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
INVx2_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_221), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
OR2x2_ASAP7_75t_L g259 ( .A(n_232), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g327 ( .A(n_232), .B(n_323), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_232), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g428 ( .A(n_232), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_232), .B(n_365), .Y(n_440) );
AND2x2_ASAP7_75t_L g319 ( .A(n_233), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_233), .B(n_235), .Y(n_342) );
INVx2_ASAP7_75t_L g254 ( .A(n_234), .Y(n_254) );
AND2x2_ASAP7_75t_L g282 ( .A(n_234), .B(n_255), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_234), .B(n_307), .Y(n_363) );
AND2x2_ASAP7_75t_L g277 ( .A(n_235), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g424 ( .A(n_235), .Y(n_424) );
AND2x2_ASAP7_75t_L g436 ( .A(n_235), .B(n_299), .Y(n_436) );
AND2x2_ASAP7_75t_L g262 ( .A(n_236), .B(n_252), .Y(n_262) );
INVx1_ASAP7_75t_L g357 ( .A(n_236), .Y(n_357) );
AO21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_241), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_237), .B(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g492 ( .A(n_237), .Y(n_492) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_237), .A2(n_505), .B(n_512), .Y(n_504) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_237), .A2(n_561), .B(n_568), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_237), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g255 ( .A(n_242), .B(n_256), .Y(n_255) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_246), .B(n_293), .Y(n_302) );
OR2x2_ASAP7_75t_L g434 ( .A(n_246), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g351 ( .A(n_247), .B(n_292), .Y(n_351) );
AND2x2_ASAP7_75t_L g359 ( .A(n_247), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g418 ( .A(n_247), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g442 ( .A(n_247), .B(n_289), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_248), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g429 ( .A(n_248), .B(n_292), .Y(n_429) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
AND2x2_ASAP7_75t_L g281 ( .A(n_251), .B(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g443 ( .A(n_251), .Y(n_443) );
NOR2x1_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
AND2x2_ASAP7_75t_L g329 ( .A(n_254), .B(n_262), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_254), .B(n_397), .Y(n_423) );
INVx2_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
INVx3_ASAP7_75t_L g320 ( .A(n_255), .Y(n_320) );
OR2x2_ASAP7_75t_L g348 ( .A(n_255), .B(n_349), .Y(n_348) );
AOI311xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .A3(n_263), .B(n_264), .C(n_275), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_258), .A2(n_296), .B(n_298), .C(n_300), .Y(n_295) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_SL g280 ( .A(n_260), .Y(n_280) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g298 ( .A(n_262), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_262), .B(n_278), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_262), .B(n_263), .Y(n_431) );
AND2x2_ASAP7_75t_L g353 ( .A(n_263), .B(n_267), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .B(n_270), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g411 ( .A(n_267), .B(n_299), .Y(n_411) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_268), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AND2x2_ASAP7_75t_L g296 ( .A(n_272), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g341 ( .A(n_274), .Y(n_341) );
AND2x4_ASAP7_75t_L g403 ( .A(n_274), .B(n_372), .Y(n_403) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI222xp33_ASAP7_75t_L g354 ( .A1(n_277), .A2(n_343), .B1(n_355), .B2(n_359), .C1(n_361), .C2(n_365), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_283), .C(n_286), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_324), .Y(n_347) );
INVx1_ASAP7_75t_L g369 ( .A(n_282), .Y(n_369) );
INVx1_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
OR2x2_ASAP7_75t_L g368 ( .A(n_285), .B(n_369), .Y(n_368) );
OAI21xp33_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B(n_293), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g304 ( .A(n_287), .B(n_305), .C(n_306), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_287), .A2(n_324), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_291), .Y(n_344) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_292), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g401 ( .A(n_292), .Y(n_401) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_292), .Y(n_417) );
INVx2_ASAP7_75t_L g375 ( .A(n_293), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_297), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B1(n_304), .B2(n_308), .C(n_309), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_303), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g437 ( .A(n_303), .Y(n_437) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g318 ( .A(n_310), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_310), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_310), .B(n_324), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_310), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g409 ( .A(n_310), .B(n_344), .Y(n_409) );
BUFx3_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND5xp2_ASAP7_75t_L g314 ( .A(n_315), .B(n_333), .C(n_354), .D(n_366), .E(n_381), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI32xp33_ASAP7_75t_L g406 ( .A1(n_318), .A2(n_345), .A3(n_361), .B1(n_407), .B2(n_409), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_320), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g330 ( .A(n_324), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_330), .B2(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_340), .B1(n_342), .B2(n_343), .C(n_346), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g405 ( .A(n_337), .B(n_356), .Y(n_405) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_342), .A2(n_403), .B1(n_421), .B2(n_426), .C(n_427), .Y(n_420) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_350), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g364 ( .A(n_356), .Y(n_364) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_374), .B2(n_375), .C1(n_376), .C2(n_377), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_375), .A2(n_422), .B1(n_424), .B2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_387), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B(n_394), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B(n_404), .C(n_406), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_414), .C(n_439), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g415 ( .A(n_411), .Y(n_415) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_420), .C(n_432), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_431), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g746 ( .A(n_452), .Y(n_746) );
OR3x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_652), .C(n_695), .Y(n_452) );
NAND5xp2_ASAP7_75t_L g453 ( .A(n_454), .B(n_579), .C(n_609), .D(n_626), .E(n_641), .Y(n_453) );
AOI221xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_502), .B1(n_542), .B2(n_548), .C(n_552), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_477), .Y(n_455) );
OR2x2_ASAP7_75t_L g557 ( .A(n_456), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g596 ( .A(n_456), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g614 ( .A(n_456), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_456), .B(n_550), .Y(n_631) );
OR2x2_ASAP7_75t_L g643 ( .A(n_456), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_456), .B(n_602), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_456), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_456), .B(n_580), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_456), .B(n_588), .Y(n_694) );
AND2x2_ASAP7_75t_L g726 ( .A(n_456), .B(n_490), .Y(n_726) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_456), .Y(n_734) );
INVx5_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_457), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g554 ( .A(n_457), .B(n_532), .Y(n_554) );
BUFx2_ASAP7_75t_L g576 ( .A(n_457), .Y(n_576) );
AND2x2_ASAP7_75t_L g605 ( .A(n_457), .B(n_478), .Y(n_605) );
AND2x2_ASAP7_75t_L g660 ( .A(n_457), .B(n_558), .Y(n_660) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_475), .Y(n_457) );
BUFx2_ASAP7_75t_L g481 ( .A(n_460), .Y(n_481) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_464), .A2(n_474), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_464), .A2(n_474), .B(n_537), .C(n_538), .Y(n_536) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_471), .C(n_472), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_469), .A2(n_472), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_477), .B(n_614), .Y(n_623) );
OAI32xp33_ASAP7_75t_L g637 ( .A1(n_477), .A2(n_573), .A3(n_638), .B1(n_639), .B2(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_477), .B(n_639), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_477), .B(n_557), .Y(n_680) );
INVx1_ASAP7_75t_SL g709 ( .A(n_477), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g718 ( .A(n_477), .B(n_504), .C(n_660), .D(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
INVx5_ASAP7_75t_L g551 ( .A(n_478), .Y(n_551) );
AND2x2_ASAP7_75t_L g580 ( .A(n_478), .B(n_491), .Y(n_580) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_478), .Y(n_659) );
AND2x2_ASAP7_75t_L g729 ( .A(n_478), .B(n_676), .Y(n_729) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
AOI21xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_486), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_L g602 ( .A(n_490), .B(n_551), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_490), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g636 ( .A(n_490), .B(n_558), .Y(n_636) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g550 ( .A(n_491), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g588 ( .A(n_491), .B(n_560), .Y(n_588) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_559), .Y(n_597) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_501), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_502), .A2(n_666), .B1(n_668), .B2(n_670), .C1(n_673), .C2(n_674), .Y(n_665) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_521), .Y(n_502) );
AND2x2_ASAP7_75t_L g598 ( .A(n_503), .B(n_599), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_503), .B(n_576), .C(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
INVx5_ASAP7_75t_SL g547 ( .A(n_504), .Y(n_547) );
OAI322xp33_ASAP7_75t_L g552 ( .A1(n_504), .A2(n_553), .A3(n_555), .B1(n_556), .B2(n_570), .C1(n_573), .C2(n_575), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_504), .B(n_545), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_504), .B(n_533), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g545 ( .A(n_514), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_514), .B(n_523), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_521), .B(n_583), .Y(n_638) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g617 ( .A(n_522), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
OR2x2_ASAP7_75t_L g546 ( .A(n_523), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_523), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_533), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_523), .B(n_545), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_523), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_523), .B(n_583), .Y(n_624) );
AND2x2_ASAP7_75t_L g632 ( .A(n_523), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_523), .B(n_592), .Y(n_682) );
INVx5_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g572 ( .A(n_524), .B(n_547), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_524), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_524), .B(n_533), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_524), .B(n_646), .Y(n_687) );
OR2x2_ASAP7_75t_L g703 ( .A(n_524), .B(n_647), .Y(n_703) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_524), .B(n_664), .Y(n_710) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_524), .Y(n_717) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
AND2x2_ASAP7_75t_L g571 ( .A(n_532), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g621 ( .A(n_532), .B(n_545), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_532), .B(n_547), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_532), .B(n_583), .Y(n_705) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_533), .B(n_547), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_533), .B(n_545), .Y(n_593) );
OR2x2_ASAP7_75t_L g647 ( .A(n_533), .B(n_545), .Y(n_647) );
AND2x2_ASAP7_75t_L g664 ( .A(n_533), .B(n_544), .Y(n_664) );
INVxp67_ASAP7_75t_L g686 ( .A(n_533), .Y(n_686) );
AND2x2_ASAP7_75t_L g713 ( .A(n_533), .B(n_583), .Y(n_713) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_533), .Y(n_720) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_541), .Y(n_533) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_544), .B(n_594), .Y(n_667) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g583 ( .A(n_545), .B(n_547), .Y(n_583) );
OR2x2_ASAP7_75t_L g650 ( .A(n_545), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g594 ( .A(n_546), .Y(n_594) );
OR2x2_ASAP7_75t_L g655 ( .A(n_546), .B(n_647), .Y(n_655) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g555 ( .A(n_550), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_550), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g556 ( .A(n_551), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_551), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_551), .B(n_558), .Y(n_590) );
INVx2_ASAP7_75t_L g635 ( .A(n_551), .Y(n_635) );
AND2x2_ASAP7_75t_L g648 ( .A(n_551), .B(n_588), .Y(n_648) );
AND2x2_ASAP7_75t_L g673 ( .A(n_551), .B(n_597), .Y(n_673) );
INVx1_ASAP7_75t_L g625 ( .A(n_556), .Y(n_625) );
INVx2_ASAP7_75t_SL g612 ( .A(n_557), .Y(n_612) );
INVx1_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_559), .Y(n_578) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g676 ( .A(n_560), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g645 ( .A(n_572), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g651 ( .A(n_572), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_572), .A2(n_654), .B1(n_656), .B2(n_661), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_572), .B(n_664), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_573), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g607 ( .A(n_574), .Y(n_607) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OR2x2_ASAP7_75t_L g589 ( .A(n_576), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_576), .B(n_580), .Y(n_640) );
AND2x2_ASAP7_75t_L g663 ( .A(n_576), .B(n_664), .Y(n_663) );
BUFx2_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_586), .C(n_600), .Y(n_579) );
INVx1_ASAP7_75t_L g603 ( .A(n_580), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g711 ( .A1(n_580), .A2(n_712), .B1(n_714), .B2(n_715), .C(n_718), .Y(n_711) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g730 ( .A(n_583), .Y(n_730) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g679 ( .A(n_585), .B(n_618), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_591), .C(n_595), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OAI32xp33_ASAP7_75t_L g704 ( .A1(n_593), .A2(n_594), .A3(n_657), .B1(n_694), .B2(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g736 ( .A(n_596), .B(n_635), .Y(n_736) );
AND2x2_ASAP7_75t_L g683 ( .A(n_597), .B(n_635), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_597), .B(n_605), .Y(n_701) );
AOI31xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_603), .A3(n_604), .B(n_606), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_602), .B(n_614), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_602), .B(n_612), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_602), .A2(n_632), .B1(n_722), .B2(n_725), .C(n_727), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g627 ( .A(n_607), .B(n_628), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_616), .B1(n_619), .B2(n_622), .C1(n_624), .C2(n_625), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g692 ( .A(n_611), .Y(n_692) );
INVx1_ASAP7_75t_L g714 ( .A(n_614), .Y(n_714) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_617), .A2(n_728), .B1(n_730), .B2(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g633 ( .A(n_618), .Y(n_633) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B1(n_632), .B2(n_634), .C(n_637), .Y(n_626) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g671 ( .A(n_629), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g723 ( .A(n_629), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g698 ( .A(n_634), .Y(n_698) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g662 ( .A(n_635), .Y(n_662) );
INVx1_ASAP7_75t_L g644 ( .A(n_636), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_639), .B(n_726), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_645), .B1(n_648), .B2(n_649), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g735 ( .A(n_648), .Y(n_735) );
INVxp33_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_650), .B(n_694), .Y(n_693) );
OAI32xp33_ASAP7_75t_L g684 ( .A1(n_651), .A2(n_685), .A3(n_686), .B1(n_687), .B2(n_688), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_665), .C(n_677), .D(n_689), .Y(n_652) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_660), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_674), .A2(n_690), .B1(n_707), .B2(n_710), .C(n_711), .Y(n_706) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g725 ( .A(n_676), .B(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_681), .B2(n_683), .C(n_684), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_686), .B(n_717), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_706), .C(n_721), .D(n_732), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .B(n_702), .C(n_704), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g737 ( .A(n_724), .Y(n_737) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B(n_737), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g759 ( .A(n_743), .B(n_760), .Y(n_759) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_753), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g763 ( .A(n_759), .Y(n_763) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule