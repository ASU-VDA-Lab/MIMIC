module real_jpeg_24273_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_354, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_354;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_90),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_31),
.C(n_45),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_80),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_73),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_1),
.A2(n_28),
.B1(n_170),
.B2(n_174),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_2),
.A2(n_50),
.B1(n_64),
.B2(n_67),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_2),
.A2(n_50),
.B1(n_79),
.B2(n_89),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_39),
.B1(n_64),
.B2(n_67),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_3),
.A2(n_39),
.B1(n_82),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_60),
.B1(n_64),
.B2(n_67),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_60),
.B1(n_88),
.B2(n_89),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_75),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_75),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_7),
.A2(n_75),
.B1(n_79),
.B2(n_89),
.Y(n_234)
);

INVx8_ASAP7_75t_SL g86 ( 
.A(n_8),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_9),
.A2(n_79),
.B1(n_89),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_9),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_9),
.A2(n_64),
.B1(n_67),
.B2(n_93),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_93),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_93),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_10),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_10),
.A2(n_36),
.B1(n_64),
.B2(n_67),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_10),
.A2(n_36),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_66),
.B1(n_79),
.B2(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_66),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_66),
.Y(n_163)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_347),
.C(n_352),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_345),
.B(n_350),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_344),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_295),
.A3(n_325),
.B1(n_330),
.B2(n_331),
.C(n_354),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_268),
.B(n_294),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_240),
.B(n_267),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_132),
.B(n_219),
.C(n_239),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_116),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_24),
.B(n_116),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_94),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_57),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_26),
.B(n_57),
.C(n_94),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_27),
.B(n_42),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_28),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_163),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_28),
.A2(n_37),
.B(n_152),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_28),
.A2(n_152),
.B(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_35),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_29),
.B(n_38),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_29),
.A2(n_124),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_31),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_30),
.B(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_33),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_40),
.Y(n_171)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_41),
.B(n_80),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_51),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_56),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_43),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_43),
.A2(n_53),
.B1(n_145),
.B2(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_43),
.B(n_80),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_43),
.A2(n_53),
.B(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_48),
.B1(n_70),
.B2(n_71),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_47),
.A2(n_71),
.B(n_185),
.C(n_187),
.Y(n_184)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_48),
.B(n_140),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_48),
.B(n_67),
.C(n_70),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_51),
.B(n_209),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_59),
.B(n_61),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_52),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_52),
.A2(n_143),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_52),
.A2(n_143),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_53),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_53),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_76),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_59),
.B(n_143),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_59),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_67),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_81),
.B(n_85),
.C(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_64),
.B(n_80),
.CON(n_186),
.SN(n_186)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_78),
.C(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_68),
.A2(n_73),
.B1(n_130),
.B2(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_68),
.A2(n_105),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_68),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_68),
.A2(n_73),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_68),
.A2(n_236),
.B(n_275),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_68),
.A2(n_73),
.B(n_105),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_103),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_72),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_72),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_81),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_78),
.Y(n_287)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_79),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_83),
.A2(n_90),
.B1(n_100),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_83),
.B(n_286),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_83),
.A2(n_90),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_83),
.A2(n_320),
.B(n_339),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_83),
.A2(n_90),
.B(n_257),
.Y(n_352)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_92),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_84),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_90),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_90),
.B(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_106),
.B2(n_115),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_97),
.B(n_101),
.C(n_115),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_98),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_98),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_104),
.B(n_261),
.Y(n_317)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_121),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_125),
.B(n_149),
.Y(n_225)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_218),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_213),
.B(n_217),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_197),
.B(n_212),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_180),
.B(n_196),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_159),
.B(n_179),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_166),
.B(n_178),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_165),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_172),
.B(n_177),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_191),
.C(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.C(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_230),
.C(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_242),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_266),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_251),
.B1(n_264),
.B2(n_265),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_265),
.C(n_266),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_250),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_246),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_245),
.A2(n_279),
.B(n_283),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_258),
.C(n_263),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B1(n_259),
.B2(n_263),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_256),
.B(n_301),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_270),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_278),
.B1(n_289),
.B2(n_290),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_276),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_277),
.A2(n_297),
.B1(n_309),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_289),
.C(n_293),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_288),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_285),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_311),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_311),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_309),
.C(n_310),
.Y(n_296)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_299),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_304),
.C(n_308),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_314),
.C(n_324),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_305),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_316),
.C(n_318),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_324),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_334),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_342),
.B2(n_343),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_340),
.B2(n_341),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_337),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_340),
.C(n_342),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_349),
.B(n_351),
.Y(n_350)
);


endmodule