module real_aes_7668_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_0), .A2(n_252), .B1(n_401), .B2(n_467), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_207), .B1(n_420), .B2(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_2), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_3), .A2(n_16), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_4), .A2(n_166), .B1(n_354), .B2(n_357), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_5), .A2(n_230), .B1(n_434), .B2(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_6), .Y(n_669) );
INVx1_ASAP7_75t_L g427 ( .A(n_7), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_8), .A2(n_236), .B1(n_505), .B2(n_514), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_9), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_10), .A2(n_615), .B1(n_645), .B2(n_646), .Y(n_614) );
INVx1_ASAP7_75t_L g645 ( .A(n_10), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_11), .A2(n_167), .B1(n_287), .B2(n_418), .Y(n_604) );
INVx1_ASAP7_75t_L g377 ( .A(n_12), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_13), .B(n_432), .Y(n_431) );
OA22x2_ASAP7_75t_L g282 ( .A1(n_14), .A2(n_283), .B1(n_284), .B2(n_378), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_14), .Y(n_283) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_15), .A2(n_96), .B1(n_357), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_17), .A2(n_60), .B1(n_410), .B2(n_412), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_18), .A2(n_19), .B1(n_692), .B2(n_810), .C(n_812), .Y(n_809) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_20), .B(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_21), .A2(n_197), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_22), .A2(n_87), .B1(n_699), .B2(n_740), .Y(n_739) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_23), .A2(n_77), .B1(n_292), .B2(n_297), .Y(n_300) );
INVx1_ASAP7_75t_L g784 ( .A(n_23), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_24), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_25), .A2(n_142), .B1(n_411), .B2(n_573), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_26), .A2(n_95), .B1(n_116), .B2(n_387), .C1(n_513), .C2(n_515), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_27), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_28), .A2(n_231), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g722 ( .A(n_29), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g582 ( .A1(n_30), .A2(n_84), .B1(n_248), .B2(n_374), .C1(n_426), .C2(n_583), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_31), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_32), .Y(n_590) );
INVx1_ASAP7_75t_L g371 ( .A(n_33), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_34), .A2(n_150), .B1(n_494), .B2(n_495), .Y(n_493) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_35), .A2(n_80), .B1(n_292), .B2(n_293), .Y(n_302) );
INVx1_ASAP7_75t_L g785 ( .A(n_35), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_36), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_37), .A2(n_144), .B1(n_429), .B2(n_551), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_38), .A2(n_122), .B1(n_450), .B2(n_452), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_39), .Y(n_854) );
INVx1_ASAP7_75t_L g350 ( .A(n_40), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_41), .A2(n_108), .B1(n_508), .B2(n_601), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_42), .A2(n_43), .B1(n_336), .B2(n_338), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_44), .A2(n_136), .B1(n_481), .B2(n_693), .C(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g328 ( .A(n_45), .Y(n_328) );
INVx1_ASAP7_75t_L g346 ( .A(n_46), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_47), .A2(n_258), .B1(n_513), .B2(n_515), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_48), .A2(n_135), .B1(n_410), .B2(n_412), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_49), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_50), .A2(n_133), .B1(n_529), .B2(n_636), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_51), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_52), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_53), .A2(n_232), .B1(n_488), .B2(n_489), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_54), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_55), .A2(n_109), .B1(n_452), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_56), .A2(n_196), .B1(n_412), .B2(n_695), .Y(n_743) );
INVx1_ASAP7_75t_L g813 ( .A(n_57), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_58), .A2(n_204), .B1(n_511), .B2(n_843), .Y(n_842) );
XOR2x2_ASAP7_75t_L g730 ( .A(n_59), .B(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_61), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_62), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_63), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_64), .A2(n_257), .B1(n_374), .B2(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_65), .B(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_66), .A2(n_83), .B1(n_484), .B2(n_640), .Y(n_639) );
OA22x2_ASAP7_75t_L g749 ( .A1(n_67), .A2(n_750), .B1(n_751), .B2(n_767), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_67), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_68), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_69), .B(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_70), .A2(n_156), .B1(n_407), .B2(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_71), .A2(n_178), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_72), .A2(n_143), .B1(n_402), .B2(n_464), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_73), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_74), .A2(n_152), .B1(n_763), .B2(n_838), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_75), .A2(n_107), .B1(n_305), .B2(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_76), .A2(n_259), .B1(n_395), .B2(n_471), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_78), .A2(n_79), .B1(n_352), .B2(n_357), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_81), .A2(n_255), .B1(n_305), .B2(n_443), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_82), .A2(n_211), .B1(n_411), .B2(n_447), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_85), .A2(n_224), .B1(n_583), .B2(n_699), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_86), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_88), .A2(n_788), .B1(n_816), .B2(n_817), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_88), .Y(n_816) );
AND2x2_ASAP7_75t_L g277 ( .A(n_89), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_90), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_91), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_92), .A2(n_180), .B1(n_580), .B2(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_93), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g274 ( .A(n_94), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_97), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_98), .A2(n_137), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_99), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_100), .A2(n_188), .B1(n_335), .B2(n_407), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_101), .A2(n_165), .B1(n_287), .B2(n_325), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_102), .A2(n_111), .B1(n_418), .B2(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g725 ( .A(n_103), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_104), .B(n_390), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_105), .Y(n_806) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_106), .A2(n_120), .B1(n_217), .B2(n_475), .C1(n_681), .C2(n_683), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_110), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_112), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_113), .A2(n_219), .B1(n_511), .B2(n_526), .Y(n_761) );
INVx1_ASAP7_75t_L g718 ( .A(n_114), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_115), .A2(n_172), .B1(n_310), .B2(n_318), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_117), .A2(n_208), .B1(n_538), .B2(n_540), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_118), .Y(n_801) );
AO22x2_ASAP7_75t_L g652 ( .A1(n_119), .A2(n_653), .B1(n_684), .B2(n_685), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_119), .Y(n_684) );
INVx1_ASAP7_75t_L g303 ( .A(n_121), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_123), .A2(n_125), .B1(n_692), .B2(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g720 ( .A(n_124), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_126), .A2(n_170), .B1(n_489), .B2(n_695), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g727 ( .A1(n_127), .A2(n_176), .B1(n_184), .B2(n_370), .C1(n_390), .C2(n_514), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_128), .A2(n_269), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_129), .A2(n_246), .B1(n_401), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_130), .A2(n_194), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_131), .A2(n_171), .B1(n_210), .B2(n_370), .C1(n_373), .C2(n_429), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_132), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_134), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_138), .A2(n_179), .B1(n_330), .B2(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g278 ( .A(n_139), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_140), .A2(n_268), .B1(n_335), .B2(n_338), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_141), .A2(n_237), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_145), .A2(n_153), .B1(n_480), .B2(n_637), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_146), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_147), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_148), .A2(n_250), .B1(n_497), .B2(n_498), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_149), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_151), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_154), .A2(n_238), .B1(n_402), .B2(n_699), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_155), .A2(n_220), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_157), .A2(n_264), .B1(n_318), .B2(n_763), .Y(n_762) );
AND2x6_ASAP7_75t_L g273 ( .A(n_158), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_158), .Y(n_778) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_159), .A2(n_227), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_160), .A2(n_256), .B1(n_485), .B2(n_489), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_161), .A2(n_201), .B1(n_362), .B2(n_390), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_162), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_163), .B(n_471), .Y(n_503) );
INVx1_ASAP7_75t_L g607 ( .A(n_164), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_168), .A2(n_267), .B1(n_415), .B2(n_416), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_169), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_173), .A2(n_271), .B(n_279), .C(n_786), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_174), .A2(n_262), .B1(n_439), .B2(n_495), .Y(n_701) );
INVx1_ASAP7_75t_L g712 ( .A(n_175), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_177), .Y(n_517) );
INVx1_ASAP7_75t_L g728 ( .A(n_181), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_182), .A2(n_223), .B1(n_526), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_183), .A2(n_222), .B1(n_443), .B2(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_185), .B(n_432), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_186), .B(n_373), .Y(n_798) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_187), .A2(n_239), .B1(n_292), .B2(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_189), .A2(n_244), .B1(n_439), .B2(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_190), .B(n_393), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_191), .Y(n_630) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_192), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g827 ( .A(n_193), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_193), .A2(n_827), .B1(n_831), .B2(n_857), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_195), .A2(n_200), .B1(n_442), .B2(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g815 ( .A(n_198), .Y(n_815) );
INVx1_ASAP7_75t_L g368 ( .A(n_199), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_202), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_203), .A2(n_247), .B1(n_583), .B2(n_699), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_205), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_206), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_209), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_212), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_213), .B(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_214), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_215), .A2(n_265), .B1(n_354), .B2(n_429), .Y(n_596) );
INVx1_ASAP7_75t_L g308 ( .A(n_216), .Y(n_308) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_218), .A2(n_261), .B1(n_573), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_221), .Y(n_667) );
XOR2x2_ASAP7_75t_L g382 ( .A(n_225), .B(n_383), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_226), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_227), .B(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_228), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_229), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_233), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_234), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_235), .A2(n_242), .B1(n_484), .B2(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g781 ( .A(n_239), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_240), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_241), .A2(n_266), .B1(n_393), .B2(n_674), .Y(n_697) );
INVx1_ASAP7_75t_L g388 ( .A(n_243), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_245), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_249), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_251), .B(n_471), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_253), .Y(n_618) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
INVx1_ASAP7_75t_L g333 ( .A(n_260), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_263), .A2(n_521), .B1(n_563), .B2(n_564), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_263), .Y(n_563) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_274), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_275), .A2(n_776), .B(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_611), .B1(n_771), .B2(n_772), .C(n_773), .Y(n_279) );
INVx1_ASAP7_75t_L g771 ( .A(n_280), .Y(n_771) );
AOI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_567), .B1(n_609), .B2(n_610), .Y(n_280) );
INVx1_ASAP7_75t_L g609 ( .A(n_281), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_379), .B1(n_565), .B2(n_566), .Y(n_281) );
INVx1_ASAP7_75t_L g565 ( .A(n_282), .Y(n_565) );
INVx1_ASAP7_75t_L g378 ( .A(n_284), .Y(n_378) );
OR4x1_ASAP7_75t_L g284 ( .A(n_285), .B(n_323), .C(n_341), .D(n_360), .Y(n_284) );
OAI221xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_303), .B1(n_304), .B2(n_308), .C(n_309), .Y(n_285) );
OAI221xp5_ASAP7_75t_SL g523 ( .A1(n_286), .A2(n_524), .B1(n_525), .B2(n_527), .C(n_528), .Y(n_523) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_287), .Y(n_415) );
BUFx3_ASAP7_75t_L g643 ( .A(n_287), .Y(n_643) );
BUFx3_ASAP7_75t_L g843 ( .A(n_287), .Y(n_843) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g451 ( .A(n_288), .Y(n_451) );
BUFx2_ASAP7_75t_SL g508 ( .A(n_288), .Y(n_508) );
BUFx2_ASAP7_75t_SL g692 ( .A(n_288), .Y(n_692) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_298), .Y(n_288) );
AND2x6_ASAP7_75t_L g325 ( .A(n_289), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g332 ( .A(n_289), .B(n_317), .Y(n_332) );
AND2x6_ASAP7_75t_L g370 ( .A(n_289), .B(n_359), .Y(n_370) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_290), .B(n_296), .Y(n_307) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g315 ( .A(n_291), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_296), .Y(n_322) );
AND2x2_ASAP7_75t_L g356 ( .A(n_291), .B(n_300), .Y(n_356) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
AND2x4_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g337 ( .A(n_298), .B(n_315), .Y(n_337) );
AND2x4_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_298), .B(n_315), .Y(n_535) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_299), .B(n_302), .Y(n_317) );
OR2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_302), .Y(n_327) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g359 ( .A(n_300), .B(n_302), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_301), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g444 ( .A(n_301), .Y(n_444) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g321 ( .A(n_302), .Y(n_321) );
INVx4_ASAP7_75t_L g693 ( .A(n_304), .Y(n_693) );
INVx3_ASAP7_75t_L g709 ( .A(n_304), .Y(n_709) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g452 ( .A(n_306), .Y(n_452) );
BUFx3_ASAP7_75t_L g488 ( .A(n_306), .Y(n_488) );
BUFx3_ASAP7_75t_L g509 ( .A(n_306), .Y(n_509) );
INVx2_ASAP7_75t_L g602 ( .A(n_306), .Y(n_602) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_307), .B(n_317), .Y(n_349) );
AND2x6_ASAP7_75t_L g395 ( .A(n_307), .B(n_317), .Y(n_395) );
AND2x4_ASAP7_75t_L g399 ( .A(n_307), .B(n_326), .Y(n_399) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx5_ASAP7_75t_L g411 ( .A(n_313), .Y(n_411) );
INVx2_ASAP7_75t_L g442 ( .A(n_313), .Y(n_442) );
BUFx3_ASAP7_75t_L g486 ( .A(n_313), .Y(n_486) );
INVx3_ASAP7_75t_L g497 ( .A(n_313), .Y(n_497) );
INVx1_ASAP7_75t_L g539 ( .A(n_313), .Y(n_539) );
INVx8_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_315), .B(n_317), .Y(n_661) );
INVx1_ASAP7_75t_L g358 ( .A(n_316), .Y(n_358) );
INVxp67_ASAP7_75t_L g663 ( .A(n_318), .Y(n_663) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g412 ( .A(n_319), .Y(n_412) );
BUFx2_ASAP7_75t_L g489 ( .A(n_319), .Y(n_489) );
BUFx2_ASAP7_75t_L g498 ( .A(n_319), .Y(n_498) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_319), .Y(n_808) );
INVx6_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g540 ( .A(n_320), .Y(n_540) );
INVx1_ASAP7_75t_SL g838 ( .A(n_320), .Y(n_838) );
OR2x6_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g355 ( .A(n_321), .Y(n_355) );
INVx1_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_329), .B2(n_333), .C(n_334), .Y(n_323) );
INVx4_ASAP7_75t_L g447 ( .A(n_324), .Y(n_447) );
INVx4_ASAP7_75t_L g529 ( .A(n_324), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_324), .A2(n_531), .B1(n_666), .B2(n_667), .Y(n_665) );
INVx3_ASAP7_75t_L g724 ( .A(n_324), .Y(n_724) );
INVx2_ASAP7_75t_SL g747 ( .A(n_324), .Y(n_747) );
INVx11_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx11_ASAP7_75t_L g408 ( .A(n_325), .Y(n_408) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g344 ( .A(n_327), .B(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_329), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_812) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g448 ( .A(n_331), .Y(n_448) );
INVx2_ASAP7_75t_L g484 ( .A(n_331), .Y(n_484) );
INVx6_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g511 ( .A(n_332), .Y(n_511) );
BUFx3_ASAP7_75t_L g573 ( .A(n_332), .Y(n_573) );
BUFx3_ASAP7_75t_L g606 ( .A(n_332), .Y(n_606) );
BUFx4f_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g418 ( .A(n_337), .Y(n_418) );
BUFx3_ASAP7_75t_L g439 ( .A(n_337), .Y(n_439) );
BUFx3_ASAP7_75t_L g494 ( .A(n_337), .Y(n_494) );
BUFx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_SL g420 ( .A(n_339), .Y(n_420) );
BUFx2_ASAP7_75t_L g440 ( .A(n_339), .Y(n_440) );
BUFx3_ASAP7_75t_L g481 ( .A(n_339), .Y(n_481) );
BUFx3_ASAP7_75t_L g495 ( .A(n_339), .Y(n_495) );
BUFx3_ASAP7_75t_L g580 ( .A(n_339), .Y(n_580) );
BUFx3_ASAP7_75t_L g638 ( .A(n_339), .Y(n_638) );
AND2x2_ASAP7_75t_L g443 ( .A(n_340), .B(n_444), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .B1(n_347), .B2(n_350), .C(n_351), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g544 ( .A(n_343), .Y(n_544) );
INVx1_ASAP7_75t_SL g792 ( .A(n_343), .Y(n_792) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_344), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_347), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g621 ( .A(n_348), .Y(n_621) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g502 ( .A(n_349), .Y(n_502) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g699 ( .A(n_353), .Y(n_699) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
BUFx3_ASAP7_75t_L g505 ( .A(n_354), .Y(n_505) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x4_ASAP7_75t_L g365 ( .A(n_356), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g375 ( .A(n_356), .B(n_376), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_356), .B(n_444), .Y(n_556) );
BUFx2_ASAP7_75t_SL g402 ( .A(n_357), .Y(n_402) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_357), .Y(n_467) );
BUFx3_ASAP7_75t_L g583 ( .A(n_357), .Y(n_583) );
BUFx2_ASAP7_75t_SL g740 ( .A(n_357), .Y(n_740) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g562 ( .A(n_358), .Y(n_562) );
INVx1_ASAP7_75t_L g561 ( .A(n_359), .Y(n_561) );
OAI222xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_368), .B1(n_369), .B2(n_371), .C1(n_372), .C2(n_377), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx4f_ASAP7_75t_SL g429 ( .A(n_365), .Y(n_429) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_365), .Y(n_475) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_365), .Y(n_514) );
INVx1_ASAP7_75t_L g376 ( .A(n_367), .Y(n_376) );
INVx4_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
BUFx2_ASAP7_75t_L g682 ( .A(n_369), .Y(n_682) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g426 ( .A(n_370), .Y(n_426) );
INVx2_ASAP7_75t_SL g461 ( .A(n_370), .Y(n_461) );
INVx2_ASAP7_75t_L g589 ( .A(n_370), .Y(n_589) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_370), .Y(n_624) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx4f_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g516 ( .A(n_374), .Y(n_516) );
BUFx12f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_375), .Y(n_390) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_375), .Y(n_464) );
INVx1_ASAP7_75t_L g566 ( .A(n_379), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_454), .B2(n_455), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
XNOR2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_421), .Y(n_381) );
NAND3x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_403), .C(n_413), .Y(n_383) );
NOR2x1_ASAP7_75t_SL g384 ( .A(n_385), .B(n_391), .Y(n_384) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_389), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .C(n_400), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g759 ( .A(n_394), .Y(n_759) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
BUFx4f_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
BUFx2_ASAP7_75t_L g473 ( .A(n_395), .Y(n_473) );
BUFx2_ASAP7_75t_L g675 ( .A(n_395), .Y(n_675) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx5_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
INVx2_ASAP7_75t_L g594 ( .A(n_398), .Y(n_594) );
INVx4_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g640 ( .A(n_408), .Y(n_640) );
INVx1_ASAP7_75t_L g703 ( .A(n_408), .Y(n_703) );
INVx2_ASAP7_75t_L g841 ( .A(n_408), .Y(n_841) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_411), .Y(n_695) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g835 ( .A(n_420), .Y(n_835) );
OAI22xp5_ASAP7_75t_SL g612 ( .A1(n_421), .A2(n_613), .B1(n_614), .B2(n_647), .Y(n_612) );
INVx3_ASAP7_75t_SL g613 ( .A(n_421), .Y(n_613) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_453), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_423), .B(n_436), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_430), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_427), .B(n_428), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g753 ( .A1(n_425), .A2(n_754), .B(n_755), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g794 ( .A1(n_425), .A2(n_795), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_794) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g548 ( .A(n_429), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .C(n_435), .Y(n_430) );
BUFx2_ASAP7_75t_L g714 ( .A(n_434), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_445), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g811 ( .A(n_439), .Y(n_811) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_442), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g726 ( .A(n_448), .Y(n_726) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g480 ( .A(n_451), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_451), .A2(n_525), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_520), .Y(n_455) );
AO22x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_490), .B1(n_518), .B2(n_519), .Y(n_456) );
INVx2_ASAP7_75t_L g518 ( .A(n_457), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_459), .B(n_476), .Y(n_458) );
NOR2xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_468), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_462), .B(n_463), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_461), .A2(n_547), .B1(n_548), .B2(n_549), .C(n_550), .Y(n_546) );
BUFx2_ASAP7_75t_L g551 ( .A(n_464), .Y(n_551) );
BUFx3_ASAP7_75t_L g683 ( .A(n_464), .Y(n_683) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_472), .C(n_474), .Y(n_468) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_471), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_475), .Y(n_852) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_482), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_SL g519 ( .A(n_490), .Y(n_519) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_517), .Y(n_490) );
NAND4xp75_ASAP7_75t_L g491 ( .A(n_492), .B(n_499), .C(n_506), .D(n_512), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
BUFx3_ASAP7_75t_L g636 ( .A(n_494), .Y(n_636) );
INVxp67_ASAP7_75t_L g719 ( .A(n_495), .Y(n_719) );
OA211x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_503), .C(n_504), .Y(n_499) );
OA211x2_ASAP7_75t_L g711 ( .A1(n_501), .A2(n_712), .B(n_713), .C(n_715), .Y(n_711) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g848 ( .A(n_502), .Y(n_848) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_510), .Y(n_506) );
BUFx2_ASAP7_75t_L g526 ( .A(n_509), .Y(n_526) );
INVx1_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
INVx2_ASAP7_75t_SL g626 ( .A(n_513), .Y(n_626) );
INVx2_ASAP7_75t_SL g796 ( .A(n_513), .Y(n_796) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g564 ( .A(n_521), .Y(n_564) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_522), .B(n_541), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_530), .Y(n_522) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g814 ( .A(n_529), .Y(n_814) );
OAI221xp5_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_532), .B1(n_533), .B2(n_536), .C(n_537), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_533), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g670 ( .A(n_534), .Y(n_670) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .C(n_552), .Y(n_541) );
INVxp67_ASAP7_75t_L g855 ( .A(n_551), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_557), .B2(n_558), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_554), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_799) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_556), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
BUFx3_ASAP7_75t_L g678 ( .A(n_556), .Y(n_678) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g802 ( .A(n_559), .Y(n_802) );
CKINVDCx16_ASAP7_75t_R g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g632 ( .A(n_560), .Y(n_632) );
OR2x6_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
AO22x2_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_585), .B2(n_608), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_584), .Y(n_569) );
NAND4xp75_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .C(n_578), .D(n_582), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g608 ( .A(n_585), .Y(n_608) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_607), .Y(n_585) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_597), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_590), .B(n_591), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .C(n_596), .Y(n_592) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g772 ( .A(n_611), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_648), .Y(n_611) );
INVx1_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
INVx1_ASAP7_75t_L g646 ( .A(n_615), .Y(n_646) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_633), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_622), .C(n_629), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g845 ( .A1(n_619), .A2(n_846), .B1(n_847), .B2(n_849), .C(n_850), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_621), .A2(n_791), .B1(n_792), .B2(n_793), .Y(n_790) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_623), .A2(n_734), .B(n_735), .Y(n_733) );
OAI222xp33_ASAP7_75t_L g851 ( .A1(n_623), .A2(n_852), .B1(n_853), .B2(n_854), .C1(n_855), .C2(n_856), .Y(n_851) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_632), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_641), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g672 ( .A(n_637), .Y(n_672) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_729), .B1(n_769), .B2(n_770), .Y(n_648) );
INVx1_ASAP7_75t_L g769 ( .A(n_649), .Y(n_769) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_686), .B2(n_687), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g685 ( .A(n_653), .Y(n_685) );
AND4x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_664), .C(n_673), .D(n_680), .Y(n_653) );
NOR2xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_658), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_662), .B2(n_663), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_660), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_804) );
BUFx2_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_SL g664 ( .A(n_665), .B(n_668), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_668) );
OAI221xp5_ASAP7_75t_SL g833 ( .A1(n_670), .A2(n_834), .B1(n_835), .B2(n_836), .C(n_837), .Y(n_833) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_705), .Y(n_687) );
NAND4xp75_ASAP7_75t_L g689 ( .A(n_690), .B(n_696), .C(n_700), .D(n_704), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
XOR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_728), .Y(n_705) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_707), .B(n_711), .C(n_716), .D(n_727), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_725), .B2(n_726), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g770 ( .A(n_729), .Y(n_770) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_748), .B1(n_749), .B2(n_768), .Y(n_729) );
INVx1_ASAP7_75t_L g768 ( .A(n_730), .Y(n_768) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_741), .C(n_744), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .C(n_739), .Y(n_736) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g767 ( .A(n_751), .Y(n_767) );
NAND3x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_760), .C(n_764), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
OR2x2_ASAP7_75t_SL g860 ( .A(n_775), .B(n_780), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_778), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_776), .Y(n_819) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_777), .B(n_823), .Y(n_826) );
CKINVDCx16_ASAP7_75t_R g823 ( .A(n_778), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
OAI322xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_818), .A3(n_820), .B1(n_824), .B2(n_827), .C1(n_828), .C2(n_858), .Y(n_786) );
INVx1_ASAP7_75t_L g817 ( .A(n_788), .Y(n_817) );
AND3x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_803), .C(n_809), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_794), .C(n_799), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
BUFx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx16_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g857 ( .A(n_831), .Y(n_857) );
AND2x2_ASAP7_75t_SL g831 ( .A(n_832), .B(n_844), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_839), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .Y(n_839) );
NOR2xp33_ASAP7_75t_SL g844 ( .A(n_845), .B(n_851), .Y(n_844) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
endmodule