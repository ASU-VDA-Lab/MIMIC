module real_aes_7108_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_1), .A2(n_138), .B(n_142), .C(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_2), .A2(n_174), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g470 ( .A(n_3), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_4), .A2(n_457), .B1(n_737), .B2(n_740), .C1(n_743), .C2(n_744), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_5), .B(n_214), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_6), .A2(n_174), .B(n_498), .Y(n_497) );
AND2x6_ASAP7_75t_L g138 ( .A(n_7), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g197 ( .A(n_8), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_9), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_9), .B(n_40), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_10), .A2(n_173), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_11), .B(n_150), .Y(n_241) );
INVx1_ASAP7_75t_L g502 ( .A(n_12), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_13), .B(n_208), .Y(n_525) );
INVx1_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
INVx1_ASAP7_75t_L g547 ( .A(n_15), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_16), .A2(n_148), .B(n_222), .C(n_224), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_17), .B(n_214), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_18), .B(n_481), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_19), .B(n_174), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_20), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_21), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_22), .B(n_214), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_23), .B(n_150), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_24), .A2(n_182), .B(n_224), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_25), .B(n_150), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_26), .Y(n_254) );
INVx1_ASAP7_75t_L g146 ( .A(n_27), .Y(n_146) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_28), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_29), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_30), .B(n_150), .Y(n_471) );
INVx1_ASAP7_75t_L g180 ( .A(n_31), .Y(n_180) );
INVx1_ASAP7_75t_L g492 ( .A(n_32), .Y(n_492) );
INVx2_ASAP7_75t_L g136 ( .A(n_33), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_34), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_35), .A2(n_208), .B(n_267), .C(n_269), .Y(n_266) );
INVxp67_ASAP7_75t_L g181 ( .A(n_36), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_37), .A2(n_142), .B(n_145), .C(n_153), .Y(n_141) );
CKINVDCx14_ASAP7_75t_R g265 ( .A(n_38), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_39), .A2(n_138), .B(n_142), .C(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g491 ( .A(n_41), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_42), .A2(n_195), .B(n_196), .C(n_198), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_43), .B(n_150), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_44), .A2(n_47), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_44), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_45), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_46), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_47), .Y(n_124) );
INVx1_ASAP7_75t_L g206 ( .A(n_48), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_49), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_50), .B(n_174), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_51), .A2(n_142), .B1(n_211), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_52), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_53), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g193 ( .A(n_54), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_55), .A2(n_195), .B(n_269), .C(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_56), .Y(n_540) );
INVx1_ASAP7_75t_L g499 ( .A(n_57), .Y(n_499) );
INVx1_ASAP7_75t_L g139 ( .A(n_58), .Y(n_139) );
INVx1_ASAP7_75t_L g157 ( .A(n_59), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_60), .A2(n_90), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_60), .Y(n_738) );
INVx1_ASAP7_75t_SL g268 ( .A(n_61), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_62), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_63), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_64), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g257 ( .A(n_65), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_SL g480 ( .A1(n_66), .A2(n_269), .B(n_481), .C(n_482), .Y(n_480) );
INVxp67_ASAP7_75t_L g483 ( .A(n_67), .Y(n_483) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_69), .A2(n_174), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_70), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_71), .A2(n_174), .B(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_72), .Y(n_495) );
INVx1_ASAP7_75t_L g534 ( .A(n_73), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_74), .A2(n_173), .B(n_175), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_75), .Y(n_140) );
INVx1_ASAP7_75t_L g220 ( .A(n_76), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_77), .A2(n_138), .B(n_142), .C(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_78), .A2(n_102), .B1(n_115), .B2(n_747), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_79), .A2(n_174), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g223 ( .A(n_80), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_81), .B(n_147), .Y(n_516) );
INVx2_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
INVx1_ASAP7_75t_L g238 ( .A(n_83), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_84), .B(n_481), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_85), .A2(n_138), .B(n_142), .C(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OR2x2_ASAP7_75t_L g447 ( .A(n_86), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g736 ( .A(n_86), .B(n_449), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_87), .A2(n_142), .B(n_256), .C(n_259), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_88), .B(n_154), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_89), .Y(n_474) );
CKINVDCx14_ASAP7_75t_R g739 ( .A(n_90), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_91), .A2(n_138), .B(n_142), .C(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_92), .Y(n_529) );
INVx1_ASAP7_75t_L g479 ( .A(n_93), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_94), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_95), .B(n_147), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_96), .B(n_162), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_97), .B(n_162), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g210 ( .A(n_99), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_100), .A2(n_174), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g747 ( .A(n_104), .Y(n_747) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g449 ( .A(n_110), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g734 ( .A(n_111), .B(n_449), .Y(n_734) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_111), .B(n_448), .Y(n_744) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_455), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g746 ( .A(n_119), .Y(n_746) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_444), .B(n_451), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_SL g735 ( .A(n_126), .Y(n_735) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_126), .A2(n_459), .B1(n_732), .B2(n_741), .Y(n_740) );
OR5x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_338), .C(n_402), .D(n_418), .E(n_433), .Y(n_126) );
NAND4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_272), .C(n_299), .D(n_322), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_215), .B(n_226), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx3_ASAP7_75t_SL g249 ( .A(n_131), .Y(n_249) );
AND2x4_ASAP7_75t_L g285 ( .A(n_131), .B(n_274), .Y(n_285) );
OR2x2_ASAP7_75t_L g295 ( .A(n_131), .B(n_251), .Y(n_295) );
OR2x2_ASAP7_75t_L g341 ( .A(n_131), .B(n_167), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_131), .B(n_250), .Y(n_355) );
AND2x2_ASAP7_75t_L g398 ( .A(n_131), .B(n_288), .Y(n_398) );
AND2x2_ASAP7_75t_L g405 ( .A(n_131), .B(n_262), .Y(n_405) );
AND2x2_ASAP7_75t_L g424 ( .A(n_131), .B(n_314), .Y(n_424) );
AND2x2_ASAP7_75t_L g442 ( .A(n_131), .B(n_284), .Y(n_442) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_159), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_141), .C(n_154), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_133), .A2(n_235), .B(n_236), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_133), .A2(n_254), .B(n_255), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_133), .A2(n_467), .B(n_468), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_133), .A2(n_184), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_133), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
AND2x4_ASAP7_75t_L g174 ( .A(n_134), .B(n_138), .Y(n_174) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
INVx1_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx3_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx1_ASAP7_75t_L g481 ( .A(n_137), .Y(n_481) );
BUFx3_ASAP7_75t_L g153 ( .A(n_138), .Y(n_153) );
INVx4_ASAP7_75t_SL g184 ( .A(n_138), .Y(n_184) );
INVx5_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_143), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_149), .C(n_151), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_147), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_147), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_148), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_148), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_148), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx4_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_152), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_154), .A2(n_191), .B(n_200), .Y(n_190) );
INVx1_ASAP7_75t_L g233 ( .A(n_154), .Y(n_233) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_154), .A2(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_L g163 ( .A(n_155), .B(n_156), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_161), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_161), .A2(n_253), .B(n_260), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_161), .B(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_162), .A2(n_477), .B(n_484), .Y(n_476) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
INVx1_ASAP7_75t_L g407 ( .A(n_164), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_189), .Y(n_164) );
AND2x2_ASAP7_75t_L g317 ( .A(n_165), .B(n_250), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_165), .B(n_337), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g350 ( .A1(n_165), .A2(n_351), .A3(n_354), .B1(n_356), .B2(n_360), .Y(n_350) );
AND2x2_ASAP7_75t_L g420 ( .A(n_165), .B(n_314), .Y(n_420) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g284 ( .A(n_167), .B(n_251), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_167), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g326 ( .A(n_167), .B(n_273), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_167), .B(n_405), .Y(n_404) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_185), .Y(n_167) );
INVx1_ASAP7_75t_L g289 ( .A(n_168), .Y(n_289) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_168), .A2(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g512 ( .A1(n_169), .A2(n_513), .B(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_170), .A2(n_466), .B(n_473), .Y(n_465) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_170), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_170), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_172), .A2(n_186), .B(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_184), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_177), .A2(n_184), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_SL g205 ( .A1(n_177), .A2(n_184), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g219 ( .A1(n_177), .A2(n_184), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_177), .A2(n_184), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_177), .A2(n_184), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_177), .A2(n_184), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_177), .A2(n_184), .B(n_544), .C(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_182), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_182), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_182), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_183), .A2(n_240), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_188), .B(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_188), .A2(n_521), .B(n_528), .Y(n_520) );
AND2x2_ASAP7_75t_L g291 ( .A(n_189), .B(n_230), .Y(n_291) );
AND2x2_ASAP7_75t_L g367 ( .A(n_189), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g439 ( .A(n_189), .Y(n_439) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_201), .Y(n_189) );
OR2x2_ASAP7_75t_L g229 ( .A(n_190), .B(n_202), .Y(n_229) );
AND2x2_ASAP7_75t_L g246 ( .A(n_190), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_190), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
AND2x2_ASAP7_75t_L g325 ( .A(n_190), .B(n_202), .Y(n_325) );
BUFx3_ASAP7_75t_L g328 ( .A(n_190), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_190), .B(n_303), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_190), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g224 ( .A(n_199), .Y(n_224) );
INVx2_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_201), .B(n_277), .Y(n_297) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g308 ( .A(n_202), .B(n_217), .Y(n_308) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_202), .Y(n_321) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_213), .Y(n_202) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_203), .A2(n_218), .B(n_225), .Y(n_217) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_203), .A2(n_263), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_208), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g472 ( .A(n_211), .Y(n_472) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_214), .A2(n_497), .B(n_503), .Y(n_496) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_328), .Y(n_378) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_SL g247 ( .A(n_217), .Y(n_247) );
NAND3xp33_ASAP7_75t_L g296 ( .A(n_217), .B(n_297), .C(n_298), .Y(n_296) );
OR2x2_ASAP7_75t_L g304 ( .A(n_217), .B(n_277), .Y(n_304) );
AND2x2_ASAP7_75t_L g324 ( .A(n_217), .B(n_277), .Y(n_324) );
AND2x2_ASAP7_75t_L g368 ( .A(n_217), .B(n_232), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_245), .B(n_248), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g443 ( .A(n_228), .B(n_368), .Y(n_443) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_229), .A2(n_341), .B1(n_383), .B2(n_385), .Y(n_382) );
OR2x2_ASAP7_75t_L g389 ( .A(n_229), .B(n_304), .Y(n_389) );
OR2x2_ASAP7_75t_L g413 ( .A(n_229), .B(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_229), .B(n_333), .Y(n_426) );
AND2x2_ASAP7_75t_L g319 ( .A(n_230), .B(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_230), .A2(n_392), .B(n_407), .Y(n_406) );
AOI32xp33_ASAP7_75t_L g427 ( .A1(n_230), .A2(n_317), .A3(n_428), .B1(n_430), .B2(n_431), .Y(n_427) );
OR2x2_ASAP7_75t_L g438 ( .A(n_230), .B(n_439), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g306 ( .A(n_231), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_231), .B(n_320), .Y(n_385) );
BUFx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g277 ( .A(n_232), .Y(n_277) );
AND2x2_ASAP7_75t_L g343 ( .A(n_232), .B(n_308), .Y(n_343) );
AND3x2_ASAP7_75t_L g352 ( .A(n_232), .B(n_246), .C(n_353), .Y(n_352) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_243), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_233), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_233), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_233), .B(n_540), .Y(n_539) );
O2A1O1Ixp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_241), .C(n_242), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_239), .A2(n_242), .B(n_257), .C(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_242), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_242), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g278 ( .A(n_247), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_247), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_247), .B(n_277), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x2_ASAP7_75t_L g273 ( .A(n_249), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g313 ( .A(n_249), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_249), .B(n_262), .Y(n_331) );
AND2x2_ASAP7_75t_L g349 ( .A(n_249), .B(n_251), .Y(n_349) );
OR2x2_ASAP7_75t_L g363 ( .A(n_249), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g409 ( .A(n_249), .B(n_337), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_250), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_262), .Y(n_250) );
AND2x2_ASAP7_75t_L g310 ( .A(n_251), .B(n_288), .Y(n_310) );
OR2x2_ASAP7_75t_L g364 ( .A(n_251), .B(n_288), .Y(n_364) );
AND2x2_ASAP7_75t_L g417 ( .A(n_251), .B(n_274), .Y(n_417) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g315 ( .A(n_252), .Y(n_315) );
AND2x2_ASAP7_75t_L g337 ( .A(n_252), .B(n_262), .Y(n_337) );
INVx2_ASAP7_75t_L g274 ( .A(n_262), .Y(n_274) );
INVx1_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_270), .Y(n_526) );
AOI211xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_280), .C(n_292), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_273), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g436 ( .A(n_273), .Y(n_436) );
AND2x2_ASAP7_75t_L g314 ( .A(n_274), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_277), .B(n_278), .Y(n_286) );
INVx1_ASAP7_75t_L g371 ( .A(n_277), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_277), .B(n_298), .Y(n_395) );
AND2x2_ASAP7_75t_L g411 ( .A(n_277), .B(n_325), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_278), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_286), .B1(n_287), .B2(n_290), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_283), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_284), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_SL g374 ( .A1(n_285), .A2(n_327), .B1(n_375), .B2(n_380), .C(n_382), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_285), .B(n_348), .Y(n_381) );
INVx1_ASAP7_75t_L g441 ( .A(n_287), .Y(n_441) );
BUFx3_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g357 ( .A(n_294), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_294), .B(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_295), .B(n_348), .Y(n_359) );
INVxp67_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g320 ( .A(n_298), .B(n_321), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_305), .B(n_309), .C(n_311), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_SL g334 ( .A(n_302), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_303), .B(n_334), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_303), .B(n_325), .Y(n_376) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_306), .A2(n_312), .B1(n_316), .B2(n_318), .Y(n_311) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g327 ( .A(n_308), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g372 ( .A(n_308), .B(n_373), .Y(n_372) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_310), .A2(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_314), .A2(n_323), .B1(n_326), .B2(n_327), .C(n_329), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_314), .B(n_348), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_314), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g430 ( .A(n_320), .Y(n_430) );
INVxp67_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
INVx1_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g399 ( .A(n_324), .B(n_328), .Y(n_399) );
INVx1_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_328), .B(n_343), .Y(n_403) );
OAI32xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .A3(n_334), .B1(n_335), .B2(n_336), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_SL g342 ( .A(n_337), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_337), .B(n_369), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_337), .B(n_398), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_337), .B(n_348), .Y(n_437) );
NAND5xp2_ASAP7_75t_L g338 ( .A(n_339), .B(n_361), .C(n_374), .D(n_386), .E(n_387), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .B1(n_344), .B2(n_346), .C(n_350), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp33_ASAP7_75t_SL g365 ( .A(n_345), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_348), .B(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_349), .A2(n_362), .B1(n_365), .B2(n_369), .Y(n_361) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OAI211xp5_ASAP7_75t_SL g356 ( .A1(n_352), .A2(n_357), .B(n_358), .C(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g384 ( .A(n_364), .Y(n_384) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_373), .B(n_422), .Y(n_432) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_392), .B2(n_396), .C1(n_399), .C2(n_400), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_402) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_415), .Y(n_410) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g422 ( .A(n_414), .Y(n_422) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B(n_438), .C(n_440), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_451), .B(n_456), .C(n_745), .Y(n_455) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_732), .B1(n_735), .B2(n_736), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR4x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_621), .C(n_681), .D(n_708), .Y(n_459) );
NAND4xp25_ASAP7_75t_SL g460 ( .A(n_461), .B(n_569), .C(n_600), .D(n_617), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_504), .B(n_506), .C(n_549), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_485), .Y(n_462) );
INVx1_ASAP7_75t_L g611 ( .A(n_463), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_463), .A2(n_652), .B1(n_700), .B2(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_464), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g562 ( .A(n_464), .B(n_487), .Y(n_562) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_464), .B(n_505), .Y(n_616) );
INVx1_ASAP7_75t_L g656 ( .A(n_464), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_464), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g584 ( .A(n_465), .B(n_487), .Y(n_584) );
INVx3_ASAP7_75t_L g588 ( .A(n_465), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_465), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g675 ( .A(n_475), .B(n_496), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_475), .B(n_588), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_475), .B(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g505 ( .A(n_476), .B(n_487), .Y(n_505) );
INVx1_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
BUFx2_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g605 ( .A(n_476), .B(n_486), .Y(n_605) );
OR2x2_ASAP7_75t_L g644 ( .A(n_476), .B(n_486), .Y(n_644) );
AND2x2_ASAP7_75t_L g669 ( .A(n_476), .B(n_496), .Y(n_669) );
AND2x2_ASAP7_75t_L g728 ( .A(n_476), .B(n_558), .Y(n_728) );
INVx1_ASAP7_75t_L g703 ( .A(n_485), .Y(n_703) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_486), .B(n_496), .Y(n_589) );
AND2x2_ASAP7_75t_L g599 ( .A(n_486), .B(n_588), .Y(n_599) );
BUFx2_ASAP7_75t_L g610 ( .A(n_486), .Y(n_610) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g632 ( .A(n_487), .B(n_496), .Y(n_632) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_487), .Y(n_687) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_496), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g558 ( .A(n_496), .Y(n_558) );
BUFx2_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
INVx2_ASAP7_75t_L g602 ( .A(n_496), .Y(n_602) );
AND2x2_ASAP7_75t_L g664 ( .A(n_496), .B(n_588), .Y(n_664) );
AOI321xp33_ASAP7_75t_L g683 ( .A1(n_504), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_505), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_505), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g677 ( .A(n_505), .B(n_656), .Y(n_677) );
AND2x2_ASAP7_75t_L g710 ( .A(n_505), .B(n_602), .Y(n_710) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_530), .Y(n_507) );
OR2x2_ASAP7_75t_L g612 ( .A(n_508), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_511), .B(n_532), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_511), .B(n_554), .Y(n_579) );
INVx1_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_511), .B(n_577), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_511), .B(n_553), .Y(n_620) );
OR2x2_ASAP7_75t_L g652 ( .A(n_511), .B(n_641), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_511), .B(n_565), .Y(n_691) );
AND2x2_ASAP7_75t_L g725 ( .A(n_511), .B(n_551), .Y(n_725) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_L g552 ( .A(n_520), .Y(n_552) );
INVx2_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_520), .B(n_578), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_520), .B(n_554), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g713 ( .A(n_531), .B(n_564), .Y(n_713) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
INVx2_ASAP7_75t_L g554 ( .A(n_532), .Y(n_554) );
AND2x2_ASAP7_75t_L g707 ( .A(n_532), .B(n_567), .Y(n_707) );
AND2x2_ASAP7_75t_L g553 ( .A(n_541), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g568 ( .A(n_541), .Y(n_568) );
INVx1_ASAP7_75t_L g578 ( .A(n_541), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_555), .B1(n_559), .B2(n_563), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_550), .A2(n_668), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_554), .B(n_567), .Y(n_641) );
INVx1_ASAP7_75t_L g657 ( .A(n_554), .Y(n_657) );
AND2x2_ASAP7_75t_L g598 ( .A(n_556), .B(n_599), .Y(n_598) );
INVx3_ASAP7_75t_SL g637 ( .A(n_556), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_556), .B(n_562), .Y(n_714) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g723 ( .A(n_559), .Y(n_723) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_560), .B(n_656), .Y(n_698) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_SL g603 ( .A(n_562), .Y(n_603) );
NAND2x1_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g624 ( .A(n_564), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_568), .Y(n_631) );
AND2x2_ASAP7_75t_L g636 ( .A(n_564), .B(n_577), .Y(n_636) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_564), .Y(n_685) );
OAI311xp33_ASAP7_75t_L g708 ( .A1(n_565), .A2(n_709), .A3(n_711), .B1(n_712), .C1(n_722), .Y(n_708) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g721 ( .A(n_566), .B(n_594), .Y(n_721) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g577 ( .A(n_567), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g625 ( .A(n_567), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g680 ( .A(n_567), .Y(n_680) );
INVx1_ASAP7_75t_L g573 ( .A(n_568), .Y(n_573) );
INVx1_ASAP7_75t_L g593 ( .A(n_568), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_568), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g626 ( .A(n_568), .Y(n_626) );
AOI221xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_572), .B1(n_580), .B2(n_585), .C(n_590), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx4_ASAP7_75t_L g594 ( .A(n_574), .Y(n_594) );
AND2x2_ASAP7_75t_L g688 ( .A(n_574), .B(n_607), .Y(n_688) );
AND2x2_ASAP7_75t_L g695 ( .A(n_574), .B(n_577), .Y(n_695) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_577), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g606 ( .A(n_579), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_582), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g731 ( .A(n_584), .B(n_675), .Y(n_731) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g716 ( .A(n_588), .B(n_644), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_589), .A2(n_682), .B(n_683), .C(n_696), .Y(n_681) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_595), .B(n_597), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g660 ( .A(n_594), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_595), .A2(n_690), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_689) );
AND2x2_ASAP7_75t_L g666 ( .A(n_596), .B(n_607), .Y(n_666) );
AND2x2_ASAP7_75t_L g719 ( .A(n_596), .B(n_614), .Y(n_719) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_599), .B(n_637), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B(n_606), .C(n_608), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g647 ( .A(n_602), .B(n_605), .Y(n_647) );
OR2x2_ASAP7_75t_L g690 ( .A(n_602), .B(n_644), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_603), .B(n_669), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_603), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g634 ( .A(n_604), .Y(n_634) );
INVx1_ASAP7_75t_L g700 ( .A(n_607), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_615), .B2(n_616), .Y(n_608) );
INVx1_ASAP7_75t_L g623 ( .A(n_609), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_610), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g686 ( .A(n_611), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g672 ( .A(n_613), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_614), .B(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_615), .A2(n_674), .B1(n_676), .B2(n_678), .Y(n_673) );
INVx1_ASAP7_75t_L g682 ( .A(n_618), .Y(n_682) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g724 ( .A(n_619), .B(n_719), .Y(n_724) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_620), .A2(n_654), .B1(n_657), .B2(n_658), .C1(n_661), .C2(n_662), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_622), .B(n_642), .C(n_653), .D(n_665), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_627), .B2(n_632), .C(n_633), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_625), .B(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_627), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_704), .Y(n_696) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g639 ( .A(n_631), .B(n_640), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_632), .A2(n_694), .B(n_695), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_648), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g684 ( .A(n_655), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_656), .B(n_675), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_656), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_660), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g692 ( .A(n_664), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_670), .B2(n_672), .C(n_673), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_675), .A2(n_713), .B1(n_714), .B2(n_715), .C1(n_717), .C2(n_720), .Y(n_712) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_679), .B(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g711 ( .A(n_685), .Y(n_711) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp33_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g742 ( .A(n_736), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_737), .Y(n_743) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule