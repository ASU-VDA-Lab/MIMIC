module fake_jpeg_12897_n_660 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_660);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_660;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_16),
.A2(n_14),
.B(n_6),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_67),
.Y(n_192)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_87),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_48),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_84),
.B(n_130),
.Y(n_145)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_18),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_90),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_27),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_97),
.Y(n_167)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_92),
.Y(n_204)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_93),
.Y(n_132)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_94),
.Y(n_216)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_96),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_31),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_110),
.Y(n_217)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_15),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_24),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_126),
.Y(n_189)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g153 ( 
.A(n_120),
.Y(n_153)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_32),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_40),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_129),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_40),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_87),
.A2(n_62),
.B1(n_28),
.B2(n_41),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_146),
.A2(n_160),
.B1(n_185),
.B2(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_154),
.B(n_159),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_92),
.B(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_157),
.B(n_170),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_42),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_62),
.B1(n_42),
.B2(n_60),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_176),
.B(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_180),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_94),
.B(n_39),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_184),
.B(n_198),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_101),
.A2(n_60),
.B1(n_45),
.B2(n_57),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_64),
.A2(n_29),
.B1(n_39),
.B2(n_56),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_186),
.A2(n_54),
.B1(n_26),
.B2(n_24),
.Y(n_287)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_187),
.Y(n_283)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_194),
.B(n_199),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_65),
.A2(n_29),
.B1(n_56),
.B2(n_43),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_52),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_57),
.C(n_51),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_73),
.A2(n_52),
.B1(n_43),
.B2(n_45),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_203),
.A2(n_214),
.B1(n_54),
.B2(n_26),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_51),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_130),
.B(n_58),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_86),
.A2(n_90),
.B1(n_81),
.B2(n_102),
.Y(n_214)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_145),
.A2(n_36),
.B1(n_76),
.B2(n_71),
.Y(n_218)
);

AO21x2_ASAP7_75t_SL g327 ( 
.A1(n_218),
.A2(n_222),
.B(n_153),
.Y(n_327)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_143),
.A2(n_67),
.A3(n_128),
.B1(n_125),
.B2(n_119),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_220),
.B(n_226),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_134),
.A2(n_83),
.B1(n_66),
.B2(n_103),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_58),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_232),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_224),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_227),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_228),
.B(n_231),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_71),
.B1(n_33),
.B2(n_50),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_20),
.B1(n_55),
.B2(n_53),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_76),
.B(n_50),
.C(n_20),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_167),
.B(n_33),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_236),
.B(n_292),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_133),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_237),
.B(n_244),
.Y(n_354)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_238),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_186),
.A2(n_129),
.B1(n_118),
.B2(n_79),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_239),
.A2(n_287),
.B1(n_290),
.B2(n_177),
.Y(n_318)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_135),
.Y(n_240)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_137),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_246),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_247),
.Y(n_328)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g305 ( 
.A(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_161),
.A2(n_88),
.B1(n_53),
.B2(n_55),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_250),
.A2(n_253),
.B1(n_192),
.B2(n_196),
.Y(n_304)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_151),
.A2(n_79),
.B1(n_108),
.B2(n_120),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_262),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_263),
.Y(n_350)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_265),
.Y(n_323)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_164),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_166),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_277),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_132),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_268),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_139),
.A2(n_120),
.B1(n_108),
.B2(n_24),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_271),
.A2(n_279),
.B(n_218),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_171),
.A2(n_163),
.A3(n_156),
.B1(n_202),
.B2(n_192),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_282),
.Y(n_329)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_275),
.B1(n_286),
.B2(n_289),
.Y(n_296)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_175),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_171),
.B(n_24),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_294),
.Y(n_307)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_279),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_134),
.A2(n_24),
.B1(n_26),
.B2(n_54),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_211),
.B1(n_207),
.B2(n_162),
.Y(n_322)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_282),
.Y(n_334)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_284),
.B(n_285),
.Y(n_353)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_288),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_179),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_149),
.A2(n_54),
.B1(n_26),
.B2(n_2),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_227),
.B1(n_262),
.B2(n_234),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_144),
.B(n_0),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_196),
.B(n_14),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_12),
.Y(n_308)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_138),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_239),
.A2(n_162),
.B1(n_195),
.B2(n_165),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_297),
.A2(n_306),
.B1(n_326),
.B2(n_327),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_223),
.B(n_236),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_300),
.B(n_12),
.C(n_11),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_270),
.A2(n_195),
.B1(n_182),
.B2(n_174),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_302),
.A2(n_321),
.B1(n_329),
.B2(n_346),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_270),
.A2(n_220),
.B1(n_266),
.B2(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_221),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_225),
.B(n_155),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_312),
.B(n_257),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_322),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_225),
.A2(n_278),
.B1(n_256),
.B2(n_269),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_282),
.A2(n_165),
.B1(n_182),
.B2(n_174),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_243),
.A2(n_173),
.B1(n_213),
.B2(n_152),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_333),
.A2(n_344),
.B(n_304),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_337),
.A2(n_238),
.B1(n_261),
.B2(n_259),
.Y(n_359)
);

AO22x1_ASAP7_75t_SL g342 ( 
.A1(n_272),
.A2(n_152),
.B1(n_54),
.B2(n_26),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_219),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_292),
.A2(n_173),
.B1(n_150),
.B2(n_168),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_218),
.A2(n_210),
.B1(n_168),
.B2(n_2),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_224),
.B1(n_294),
.B2(n_286),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_290),
.A2(n_222),
.B1(n_240),
.B2(n_232),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_355),
.B1(n_283),
.B2(n_246),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_222),
.A2(n_210),
.B1(n_12),
.B2(n_11),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_340),
.A2(n_271),
.B1(n_222),
.B2(n_291),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_362),
.B1(n_370),
.B2(n_391),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_359),
.A2(n_368),
.B1(n_385),
.B2(n_311),
.Y(n_429)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_276),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_374),
.C(n_390),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

OAI21xp33_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_373),
.B(n_386),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_295),
.A2(n_242),
.B1(n_267),
.B2(n_283),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_366),
.A2(n_380),
.B(n_381),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_384),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_273),
.B1(n_288),
.B2(n_284),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_372),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_SL g373 ( 
.A(n_310),
.B(n_255),
.C(n_241),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_258),
.Y(n_374)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_378),
.A2(n_311),
.B1(n_328),
.B2(n_347),
.Y(n_436)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_344),
.A2(n_295),
.B(n_339),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_248),
.B(n_264),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_382),
.Y(n_435)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

OAI32xp33_ASAP7_75t_L g387 ( 
.A1(n_310),
.A2(n_254),
.A3(n_245),
.B1(n_249),
.B2(n_251),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_393),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_322),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_300),
.B(n_281),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_252),
.B1(n_275),
.B2(n_274),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_348),
.A2(n_260),
.B1(n_265),
.B2(n_277),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_399),
.B(n_296),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_235),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_327),
.A2(n_318),
.B1(n_307),
.B2(n_342),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_394),
.A2(n_396),
.B1(n_327),
.B2(n_353),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_395),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_327),
.A2(n_233),
.B1(n_1),
.B2(n_3),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_314),
.B(n_0),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_402),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_314),
.B(n_12),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_398),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_307),
.A2(n_233),
.B(n_3),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_323),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_400),
.Y(n_426)
);

INVx13_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_401),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_308),
.B(n_1),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_404),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_307),
.B(n_3),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_376),
.B1(n_378),
.B2(n_362),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_413),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_321),
.C(n_352),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_414),
.B(n_421),
.C(n_423),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_334),
.C(n_312),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_380),
.A2(n_399),
.B(n_388),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_445),
.B(n_398),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_334),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_357),
.A2(n_353),
.B1(n_342),
.B2(n_327),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_424),
.A2(n_442),
.B1(n_400),
.B2(n_364),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_334),
.C(n_330),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_431),
.C(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_360),
.A2(n_342),
.B1(n_355),
.B2(n_333),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_436),
.B1(n_440),
.B2(n_389),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_353),
.C(n_346),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_360),
.B(n_331),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_437),
.A2(n_373),
.B(n_361),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_389),
.A2(n_376),
.B1(n_396),
.B2(n_358),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_438),
.A2(n_391),
.B1(n_404),
.B2(n_397),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_370),
.A2(n_336),
.B1(n_349),
.B2(n_343),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_331),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_387),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_357),
.A2(n_336),
.B1(n_315),
.B2(n_338),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_399),
.A2(n_331),
.B(n_349),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_446),
.A2(n_448),
.B1(n_450),
.B2(n_465),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_451),
.B1(n_464),
.B2(n_479),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_389),
.B1(n_381),
.B2(n_366),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_395),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_452),
.Y(n_489)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_405),
.B(n_402),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_470),
.C(n_481),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_406),
.B(n_367),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_455),
.B(n_458),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_457),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_365),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_461),
.B(n_421),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_433),
.B1(n_441),
.B2(n_444),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_424),
.A2(n_369),
.B1(n_372),
.B2(n_382),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_443),
.A2(n_384),
.B1(n_371),
.B2(n_377),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_467),
.A2(n_426),
.B(n_428),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_409),
.A2(n_403),
.B1(n_401),
.B2(n_383),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_468),
.A2(n_469),
.B1(n_472),
.B2(n_475),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_409),
.A2(n_401),
.B1(n_385),
.B2(n_375),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_405),
.B(n_323),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_410),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_474),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_444),
.A2(n_437),
.B1(n_442),
.B2(n_413),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_418),
.B(n_379),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_375),
.B1(n_385),
.B2(n_341),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_478),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_445),
.A2(n_341),
.B1(n_347),
.B2(n_350),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_477),
.A2(n_420),
.B1(n_439),
.B2(n_430),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_319),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_324),
.B1(n_335),
.B2(n_350),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_319),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_423),
.B(n_325),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_416),
.A2(n_332),
.B1(n_325),
.B2(n_324),
.Y(n_482)
);

OA22x2_ASAP7_75t_L g513 ( 
.A1(n_482),
.A2(n_436),
.B1(n_435),
.B2(n_415),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_483),
.B(n_490),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_447),
.A2(n_432),
.B1(n_410),
.B2(n_414),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_486),
.A2(n_449),
.B1(n_471),
.B2(n_467),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_458),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_487),
.B(n_496),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_462),
.B(n_425),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_493),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_452),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g498 ( 
.A1(n_456),
.A2(n_472),
.B1(n_448),
.B2(n_451),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_475),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_474),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_508),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_419),
.C(n_434),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_506),
.C(n_507),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_455),
.B(n_434),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_503),
.B(n_516),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_419),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_509),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_431),
.C(n_432),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_462),
.B(n_428),
.C(n_417),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_478),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_417),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_415),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_511),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_435),
.Y(n_511)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_513),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_461),
.B(n_332),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_477),
.C(n_480),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_443),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_517),
.A2(n_453),
.B1(n_420),
.B2(n_439),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_522),
.B(n_505),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_515),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_524),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_495),
.A2(n_450),
.B1(n_469),
.B2(n_471),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_525),
.A2(n_505),
.B1(n_491),
.B2(n_486),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_488),
.A2(n_446),
.B1(n_465),
.B2(n_461),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_526),
.A2(n_536),
.B1(n_542),
.B2(n_491),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_543),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_468),
.C(n_463),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_529),
.B(n_534),
.C(n_544),
.Y(n_569)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_494),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_533),
.Y(n_560)
);

FAx1_ASAP7_75t_SL g533 ( 
.A(n_506),
.B(n_479),
.CI(n_476),
.CON(n_533),
.SN(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_459),
.C(n_457),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_535),
.A2(n_484),
.B1(n_512),
.B2(n_513),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_489),
.A2(n_473),
.B1(n_430),
.B2(n_335),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_500),
.B(n_317),
.Y(n_537)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_317),
.Y(n_539)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_539),
.Y(n_557)
);

AOI22x1_ASAP7_75t_SL g540 ( 
.A1(n_498),
.A2(n_305),
.B1(n_313),
.B2(n_316),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_540),
.A2(n_517),
.B(n_513),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_497),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_541),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_499),
.A2(n_316),
.B1(n_313),
.B2(n_303),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_483),
.B(n_305),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_298),
.C(n_303),
.Y(n_544)
);

AOI22x1_ASAP7_75t_L g545 ( 
.A1(n_485),
.A2(n_305),
.B1(n_298),
.B2(n_11),
.Y(n_545)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_545),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_514),
.B(n_10),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_509),
.Y(n_566)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_497),
.Y(n_548)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_494),
.B(n_4),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_549),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_526),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_510),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_555),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_554),
.A2(n_558),
.B1(n_518),
.B2(n_531),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_502),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_556),
.A2(n_535),
.B1(n_533),
.B2(n_549),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_530),
.A2(n_485),
.B1(n_499),
.B2(n_498),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_559),
.A2(n_558),
.B(n_560),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_562),
.A2(n_565),
.B1(n_532),
.B2(n_518),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_531),
.A2(n_498),
.B1(n_513),
.B2(n_484),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_566),
.B(n_573),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_492),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_575),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_536),
.A2(n_512),
.B1(n_493),
.B2(n_490),
.Y(n_570)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_570),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_4),
.C(n_5),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_519),
.B(n_6),
.C(n_7),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_574),
.B(n_546),
.C(n_544),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_519),
.B(n_6),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_577),
.B(n_590),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_560),
.Y(n_578)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_578),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_585),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_580),
.A2(n_592),
.B1(n_594),
.B2(n_597),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_527),
.C(n_538),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_589),
.C(n_568),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_561),
.A2(n_547),
.B1(n_523),
.B2(n_548),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_582),
.A2(n_584),
.B1(n_588),
.B2(n_556),
.Y(n_605)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_586),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_557),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_587),
.B(n_588),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_563),
.A2(n_528),
.B1(n_537),
.B2(n_521),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_527),
.C(n_538),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_564),
.B(n_555),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_559),
.A2(n_540),
.B(n_533),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_591),
.A2(n_562),
.B1(n_567),
.B2(n_572),
.Y(n_602)
);

A2O1A1Ixp33_ASAP7_75t_SL g594 ( 
.A1(n_563),
.A2(n_545),
.B(n_543),
.C(n_542),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_594),
.A2(n_8),
.B(n_580),
.Y(n_613)
);

OAI21x1_ASAP7_75t_SL g595 ( 
.A1(n_565),
.A2(n_545),
.B(n_7),
.Y(n_595)
);

INVx11_ASAP7_75t_L g598 ( 
.A(n_595),
.Y(n_598)
);

FAx1_ASAP7_75t_SL g596 ( 
.A(n_571),
.B(n_6),
.CI(n_7),
.CON(n_596),
.SN(n_596)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_596),
.A2(n_573),
.B(n_567),
.C(n_574),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_600),
.B(n_602),
.Y(n_620)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_605),
.A2(n_598),
.B1(n_616),
.B2(n_603),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_583),
.A2(n_551),
.B1(n_550),
.B2(n_566),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_607),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_550),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_576),
.B(n_552),
.C(n_575),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_608),
.B(n_609),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_576),
.B(n_9),
.C(n_7),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_7),
.C(n_8),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_612),
.C(n_577),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_8),
.C(n_589),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_613),
.A2(n_596),
.B(n_598),
.Y(n_626)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_614),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_578),
.B(n_584),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_605),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_616),
.A2(n_613),
.B1(n_599),
.B2(n_603),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_617),
.B(n_629),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_599),
.A2(n_579),
.B(n_594),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_619),
.A2(n_629),
.B(n_626),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_615),
.A2(n_594),
.B(n_581),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_627),
.Y(n_641)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_601),
.Y(n_623)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_623),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_611),
.A2(n_596),
.B(n_615),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_624),
.A2(n_631),
.B(n_604),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_626),
.Y(n_636)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_628),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_601),
.B(n_614),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_620),
.B(n_612),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_642),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_618),
.B(n_600),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_633),
.B(n_640),
.Y(n_650)
);

AO21x1_ASAP7_75t_L g644 ( 
.A1(n_637),
.A2(n_631),
.B(n_622),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_621),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_630),
.B(n_608),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_607),
.Y(n_642)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_643),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_644),
.A2(n_647),
.B(n_649),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_634),
.A2(n_625),
.B(n_619),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_645),
.B(n_646),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_641),
.A2(n_625),
.B(n_617),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_639),
.B(n_609),
.C(n_610),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_637),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g653 ( 
.A1(n_648),
.A2(n_641),
.B(n_636),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_653),
.B(n_650),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_650),
.C(n_636),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_655),
.B(n_656),
.Y(n_657)
);

BUFx24_ASAP7_75t_SL g658 ( 
.A(n_657),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_658),
.A2(n_651),
.B(n_652),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_635),
.Y(n_660)
);


endmodule