module fake_jpeg_2186_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_50),
.Y(n_126)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_2),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_65),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_5),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_38),
.B1(n_34),
.B2(n_26),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_29),
.B(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_69),
.B(n_75),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_28),
.B1(n_11),
.B2(n_13),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_16),
.Y(n_77)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_35),
.C(n_31),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_87),
.C(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_102),
.B1(n_116),
.B2(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_31),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_41),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_30),
.B1(n_41),
.B2(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_41),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_54),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_28),
.B1(n_22),
.B2(n_12),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_94),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_22),
.B1(n_11),
.B2(n_13),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_71),
.B1(n_80),
.B2(n_22),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_129),
.B(n_132),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_140),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_67),
.B(n_74),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_66),
.B1(n_76),
.B2(n_56),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_140),
.B1(n_167),
.B2(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_60),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_152),
.B1(n_154),
.B2(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_22),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_126),
.B(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_158),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_85),
.B1(n_122),
.B2(n_95),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_159),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_125),
.B1(n_101),
.B2(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_127),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_162),
.Y(n_177)
);

OR2x2_ASAP7_75t_SL g161 ( 
.A(n_86),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_93),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g163 ( 
.A(n_101),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_93),
.A2(n_111),
.B1(n_105),
.B2(n_107),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_107),
.B1(n_115),
.B2(n_117),
.Y(n_170)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_159),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_117),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_195),
.C(n_173),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_179),
.B1(n_194),
.B2(n_155),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_115),
.B1(n_131),
.B2(n_153),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_SL g214 ( 
.A(n_174),
.B(n_173),
.C(n_176),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_141),
.A3(n_148),
.B1(n_150),
.B2(n_147),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_134),
.B(n_135),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_148),
.B1(n_161),
.B2(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_142),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_198),
.B(n_202),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_145),
.B1(n_143),
.B2(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_204),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_175),
.B(n_184),
.C(n_183),
.D(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_151),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_165),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_176),
.B1(n_170),
.B2(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_136),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_210),
.C(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_181),
.C(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_228),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_200),
.B1(n_199),
.B2(n_215),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_181),
.CI(n_189),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_188),
.B(n_182),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_208),
.B1(n_202),
.B2(n_203),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_247)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_221),
.B1(n_232),
.B2(n_230),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_199),
.B1(n_204),
.B2(n_200),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_225),
.C(n_197),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_248),
.C(n_235),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_201),
.A3(n_222),
.B1(n_225),
.B2(n_228),
.C1(n_218),
.C2(n_223),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_229),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_211),
.B1(n_212),
.B2(n_188),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_242),
.B(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_238),
.B(n_239),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_247),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_248),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_245),
.C(n_220),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_261),
.B(n_241),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_239),
.B(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_251),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_260),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_228),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_262),
.C(n_217),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);


endmodule