module fake_jpeg_21997_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_0),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_22),
.B1(n_24),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_38),
.B1(n_36),
.B2(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_36),
.B1(n_18),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_70),
.B1(n_73),
.B2(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_2),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_20),
.B1(n_29),
.B2(n_34),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_29),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_77),
.C(n_23),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_20),
.B1(n_35),
.B2(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_1),
.Y(n_77)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_81),
.Y(n_119)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_37),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_42),
.C(n_43),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_91),
.C(n_109),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_94),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_43),
.B(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_58),
.B1(n_94),
.B2(n_100),
.Y(n_122)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_97),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_62),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_43),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_54),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_71),
.B(n_23),
.C(n_5),
.Y(n_134)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_118),
.B1(n_19),
.B2(n_33),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_31),
.B1(n_25),
.B2(n_19),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_52),
.B1(n_77),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_77),
.B1(n_83),
.B2(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_60),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_76),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_108),
.B(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_53),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_53),
.B1(n_63),
.B2(n_66),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_110),
.B(n_115),
.C(n_96),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_89),
.A2(n_71),
.B1(n_23),
.B2(n_6),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_152),
.B1(n_156),
.B2(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_157),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_23),
.B1(n_4),
.B2(n_7),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_167),
.B1(n_177),
.B2(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_172),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_85),
.B1(n_86),
.B2(n_107),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_106),
.B(n_105),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_146),
.B1(n_145),
.B2(n_142),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_121),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_186),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_188),
.B(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_101),
.B1(n_102),
.B2(n_114),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_3),
.B(n_4),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_9),
.B(n_11),
.Y(n_216)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_102),
.B1(n_116),
.B2(n_10),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_149),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_8),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_132),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_16),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_135),
.B(n_133),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_202),
.B(n_220),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_135),
.B(n_146),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_151),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_169),
.B1(n_178),
.B2(n_172),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_221),
.B1(n_13),
.B2(n_14),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_215),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_154),
.C(n_136),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.C(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_144),
.C(n_132),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_149),
.B(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_181),
.C(n_165),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_233),
.C(n_246),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_169),
.B1(n_179),
.B2(n_177),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_243),
.B1(n_221),
.B2(n_195),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_230),
.B(n_236),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_162),
.B1(n_188),
.B2(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_240),
.B1(n_202),
.B2(n_220),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_191),
.C(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_237),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g240 ( 
.A1(n_196),
.A2(n_189),
.B1(n_161),
.B2(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_184),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_15),
.C(n_16),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_260),
.B(n_263),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_235),
.B1(n_228),
.B2(n_246),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_212),
.C(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_265),
.C(n_242),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_216),
.B(n_206),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_262),
.A2(n_245),
.B1(n_194),
.B2(n_203),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_207),
.B(n_203),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_199),
.C(n_192),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_215),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_239),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_213),
.B1(n_218),
.B2(n_192),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_234),
.B1(n_231),
.B2(n_241),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_276),
.B1(n_284),
.B2(n_256),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_255),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_264),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_235),
.B1(n_236),
.B2(n_228),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_279),
.B1(n_270),
.B2(n_278),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.C(n_281),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_224),
.C(n_199),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_210),
.C(n_213),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_201),
.C(n_15),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_280),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_285),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_15),
.B1(n_248),
.B2(n_254),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_280),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_250),
.A3(n_263),
.B1(n_260),
.B2(n_265),
.C1(n_257),
.C2(n_253),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_256),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_294),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_272),
.C(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_275),
.C(n_281),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_304),
.C(n_308),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_268),
.B1(n_277),
.B2(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_288),
.C(n_307),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_316),
.B(n_312),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_302),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_318),
.A2(n_302),
.B(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_300),
.C(n_317),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_319),
.B(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_320),
.B(n_326),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);


endmodule