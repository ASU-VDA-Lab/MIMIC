module real_aes_7331_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_88), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g516 ( .A(n_1), .Y(n_516) );
INVx1_ASAP7_75t_L g157 ( .A(n_2), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_3), .A2(n_741), .B1(n_744), .B2(n_745), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_3), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_4), .A2(n_128), .B1(n_129), .B2(n_452), .Y(n_127) );
INVx1_ASAP7_75t_L g452 ( .A(n_4), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_5), .A2(n_41), .B1(n_182), .B2(n_472), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g201 ( .A1(n_6), .A2(n_173), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_7), .B(n_171), .Y(n_527) );
AND2x6_ASAP7_75t_L g150 ( .A(n_8), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_9), .A2(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_10), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_10), .B(n_42), .Y(n_126) );
INVx1_ASAP7_75t_L g207 ( .A(n_11), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_12), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_14), .B(n_163), .Y(n_480) );
INVx1_ASAP7_75t_L g261 ( .A(n_15), .Y(n_261) );
INVx1_ASAP7_75t_L g510 ( .A(n_16), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_17), .B(n_138), .Y(n_532) );
AO32x2_ASAP7_75t_L g499 ( .A1(n_18), .A2(n_137), .A3(n_171), .B1(n_474), .B2(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_19), .B(n_182), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_20), .B(n_178), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_21), .B(n_138), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g448 ( .A1(n_22), .A2(n_34), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_22), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_23), .A2(n_53), .B1(n_182), .B2(n_472), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_24), .B(n_173), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_25), .A2(n_104), .B1(n_112), .B2(n_753), .Y(n_103) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_26), .A2(n_79), .B1(n_163), .B2(n_182), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_27), .B(n_182), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_28), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_29), .A2(n_259), .B(n_260), .C(n_262), .Y(n_258) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_30), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_31), .B(n_168), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_32), .B(n_161), .Y(n_160) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_33), .A2(n_458), .B1(n_740), .B2(n_746), .C1(n_749), .C2(n_750), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_34), .Y(n_450) );
INVx1_ASAP7_75t_L g196 ( .A(n_35), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_36), .B(n_168), .Y(n_497) );
INVx2_ASAP7_75t_L g148 ( .A(n_37), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_38), .B(n_182), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_39), .B(n_168), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_40), .A2(n_150), .B(n_153), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g194 ( .A(n_43), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_44), .B(n_161), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_45), .B(n_182), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_46), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_47), .A2(n_89), .B1(n_225), .B2(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_48), .B(n_182), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_49), .B(n_182), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_50), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_51), .B(n_515), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_52), .B(n_173), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_54), .A2(n_63), .B1(n_163), .B2(n_182), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_55), .A2(n_153), .B1(n_163), .B2(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_56), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_57), .B(n_182), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_58), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_59), .B(n_182), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_60), .A2(n_181), .B(n_205), .C(n_206), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_61), .Y(n_252) );
INVx1_ASAP7_75t_L g203 ( .A(n_62), .Y(n_203) );
INVx1_ASAP7_75t_L g151 ( .A(n_64), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_65), .B(n_182), .Y(n_517) );
INVx1_ASAP7_75t_L g141 ( .A(n_66), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_67), .Y(n_117) );
AO32x2_ASAP7_75t_L g469 ( .A1(n_68), .A2(n_171), .A3(n_230), .B1(n_470), .B2(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g549 ( .A(n_69), .Y(n_549) );
INVx1_ASAP7_75t_L g492 ( .A(n_70), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_71), .A2(n_78), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_71), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_72), .A2(n_178), .B(n_179), .C(n_181), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_73), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_74), .B(n_163), .Y(n_493) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_76), .Y(n_199) );
INVx1_ASAP7_75t_L g245 ( .A(n_77), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_78), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_80), .A2(n_150), .B(n_153), .C(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_81), .B(n_472), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_82), .B(n_163), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_83), .B(n_158), .Y(n_221) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_85), .B(n_178), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_86), .B(n_163), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_87), .A2(n_150), .B(n_153), .C(n_156), .Y(n_152) );
OR2x2_ASAP7_75t_L g122 ( .A(n_88), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g461 ( .A(n_88), .B(n_124), .Y(n_461) );
INVx2_ASAP7_75t_L g739 ( .A(n_88), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_90), .A2(n_102), .B1(n_163), .B2(n_164), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_91), .B(n_168), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_92), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_93), .A2(n_150), .B(n_153), .C(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_94), .Y(n_240) );
INVx1_ASAP7_75t_L g176 ( .A(n_95), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_96), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_97), .B(n_158), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_98), .B(n_163), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_99), .B(n_171), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_100), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_101), .A2(n_173), .B(n_174), .Y(n_172) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g754 ( .A(n_105), .Y(n_754) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_456), .Y(n_112) );
BUFx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_114), .B(n_453), .C(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B(n_453), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_122), .Y(n_455) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_123), .B(n_739), .Y(n_752) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g738 ( .A(n_124), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_447), .B1(n_448), .B2(n_451), .Y(n_129) );
INVx2_ASAP7_75t_L g451 ( .A(n_130), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_130), .A2(n_459), .B1(n_462), .B2(n_736), .Y(n_458) );
OR4x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_336), .C(n_396), .D(n_423), .Y(n_130) );
NAND4xp25_ASAP7_75t_SL g131 ( .A(n_132), .B(n_284), .C(n_315), .D(n_332), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_209), .B(n_211), .C(n_264), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_187), .Y(n_133) );
INVx1_ASAP7_75t_L g326 ( .A(n_134), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_134), .A2(n_367), .B1(n_415), .B2(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_135), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g277 ( .A(n_135), .B(n_189), .Y(n_277) );
AND2x2_ASAP7_75t_L g319 ( .A(n_135), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_135), .B(n_210), .Y(n_331) );
INVx1_ASAP7_75t_L g371 ( .A(n_135), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_135), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g299 ( .A(n_136), .B(n_189), .Y(n_299) );
INVx3_ASAP7_75t_L g303 ( .A(n_136), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_136), .B(n_361), .Y(n_360) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_165), .Y(n_136) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_137), .A2(n_190), .B(n_198), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_137), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_139), .B(n_140), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_152), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_145), .A2(n_183), .B1(n_191), .B2(n_197), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_145), .A2(n_245), .B(n_246), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
AND2x4_ASAP7_75t_L g173 ( .A(n_146), .B(n_150), .Y(n_173) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g515 ( .A(n_147), .Y(n_515) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx3_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
INVx4_ASAP7_75t_SL g183 ( .A(n_150), .Y(n_183) );
BUFx3_ASAP7_75t_L g474 ( .A(n_150), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_150), .A2(n_478), .B(n_482), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_150), .A2(n_491), .B(n_494), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_150), .A2(n_509), .B(n_513), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_150), .A2(n_521), .B(n_524), .Y(n_520) );
INVx5_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
BUFx3_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
INVx1_ASAP7_75t_L g472 ( .A(n_154), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_160), .C(n_162), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_SL g491 ( .A1(n_158), .A2(n_181), .B(n_492), .C(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g502 ( .A(n_158), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_158), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_158), .A2(n_546), .B(n_547), .Y(n_545) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_159), .B(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_159), .B(n_207), .Y(n_206) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_159), .A2(n_161), .B1(n_471), .B2(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
INVx4_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_161), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_161), .A2(n_502), .B1(n_535), .B2(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_162), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_167), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_167), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g230 ( .A(n_168), .Y(n_230) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_168), .A2(n_254), .B(n_263), .Y(n_253) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_168), .A2(n_477), .B(n_485), .Y(n_476) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_168), .A2(n_490), .B(n_497), .Y(n_489) );
AND2x2_ASAP7_75t_L g390 ( .A(n_169), .B(n_200), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_169), .B(n_303), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_169), .B(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g210 ( .A(n_170), .B(n_189), .Y(n_210) );
INVx1_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
BUFx2_ASAP7_75t_L g276 ( .A(n_170), .Y(n_276) );
AND2x2_ASAP7_75t_L g320 ( .A(n_170), .B(n_188), .Y(n_320) );
OR2x2_ASAP7_75t_L g359 ( .A(n_170), .B(n_188), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_170), .B(n_200), .Y(n_384) );
AND2x2_ASAP7_75t_L g443 ( .A(n_170), .B(n_273), .Y(n_443) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_184), .Y(n_170) );
INVx4_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_171), .A2(n_520), .B(n_527), .Y(n_519) );
BUFx2_ASAP7_75t_L g255 ( .A(n_173), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_175), .A2(n_183), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_175), .A2(n_183), .B(n_257), .C(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g481 ( .A(n_178), .Y(n_481) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_182), .Y(n_237) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_185), .A2(n_201), .B(n_208), .Y(n_200) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_SL g227 ( .A(n_186), .B(n_228), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_186), .B(n_474), .C(n_534), .Y(n_533) );
AO21x1_ASAP7_75t_L g580 ( .A1(n_186), .A2(n_534), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g418 ( .A(n_187), .Y(n_418) );
OR2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_200), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_188), .B(n_200), .Y(n_304) );
AND2x2_ASAP7_75t_L g314 ( .A(n_188), .B(n_303), .Y(n_314) );
BUFx2_ASAP7_75t_L g325 ( .A(n_188), .Y(n_325) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g347 ( .A(n_189), .B(n_200), .Y(n_347) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_189), .Y(n_402) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g195 ( .A(n_193), .Y(n_195) );
INVx4_ASAP7_75t_L g259 ( .A(n_193), .Y(n_259) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_200), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_SL g273 ( .A(n_200), .Y(n_273) );
BUFx2_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
INVx2_ASAP7_75t_L g317 ( .A(n_200), .Y(n_317) );
AND2x2_ASAP7_75t_L g379 ( .A(n_200), .B(n_303), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_205), .A2(n_483), .B(n_484), .Y(n_482) );
O2A1O1Ixp5_ASAP7_75t_L g548 ( .A1(n_205), .A2(n_514), .B(n_549), .C(n_550), .Y(n_548) );
AOI321xp33_ASAP7_75t_L g398 ( .A1(n_209), .A2(n_399), .A3(n_400), .B1(n_401), .B2(n_403), .C(n_404), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_210), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_210), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_210), .B(n_371), .Y(n_392) );
AND2x2_ASAP7_75t_L g425 ( .A(n_210), .B(n_317), .Y(n_425) );
INVx1_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_241), .Y(n_212) );
OR2x2_ASAP7_75t_L g327 ( .A(n_213), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_229), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g279 ( .A(n_216), .Y(n_279) );
AND2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_243), .Y(n_289) );
AND2x2_ASAP7_75t_L g294 ( .A(n_216), .B(n_269), .Y(n_294) );
INVx1_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_216), .B(n_292), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_216), .B(n_268), .Y(n_335) );
OR2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_356), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_216), .B(n_280), .Y(n_406) );
AND2x2_ASAP7_75t_L g440 ( .A(n_216), .B(n_266), .Y(n_440) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
AOI21xp5_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_219), .B(n_226), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_223), .A2(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
INVx1_ASAP7_75t_L g250 ( .A(n_226), .Y(n_250) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_226), .A2(n_508), .B(n_518), .Y(n_507) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_226), .A2(n_544), .B(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
INVx2_ASAP7_75t_L g282 ( .A(n_229), .Y(n_282) );
AND2x2_ASAP7_75t_L g322 ( .A(n_229), .B(n_293), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_229), .B(n_269), .Y(n_344) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g428 ( .A(n_242), .B(n_279), .Y(n_428) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_253), .Y(n_242) );
INVx2_ASAP7_75t_L g269 ( .A(n_243), .Y(n_269) );
AND2x2_ASAP7_75t_L g422 ( .A(n_243), .B(n_282), .Y(n_422) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_250), .B(n_251), .Y(n_243) );
AND2x2_ASAP7_75t_L g268 ( .A(n_253), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g283 ( .A(n_253), .Y(n_283) );
INVx1_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_259), .B(n_261), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_259), .A2(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g512 ( .A(n_259), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_270), .B1(n_274), .B2(n_278), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_265), .A2(n_383), .B1(n_420), .B2(n_421), .Y(n_419) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g334 ( .A(n_267), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_268), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_269), .B(n_282), .Y(n_356) );
INVx1_ASAP7_75t_L g372 ( .A(n_269), .Y(n_372) );
AND2x2_ASAP7_75t_L g313 ( .A(n_271), .B(n_314), .Y(n_313) );
INVx3_ASAP7_75t_SL g352 ( .A(n_271), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_271), .B(n_277), .Y(n_429) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g438 ( .A(n_274), .Y(n_438) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_275), .B(n_371), .Y(n_413) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_SL g318 ( .A(n_277), .Y(n_318) );
NAND2x1_ASAP7_75t_SL g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g339 ( .A(n_279), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g346 ( .A(n_279), .B(n_283), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_279), .B(n_292), .Y(n_351) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_279), .Y(n_400) );
OAI311xp33_ASAP7_75t_L g423 ( .A1(n_280), .A2(n_424), .A3(n_426), .B1(n_427), .C1(n_437), .Y(n_423) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g436 ( .A(n_281), .B(n_309), .Y(n_436) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g292 ( .A(n_282), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g340 ( .A(n_282), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g395 ( .A(n_282), .Y(n_395) );
INVx1_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_283), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g341 ( .A(n_283), .Y(n_341) );
AOI221xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_287), .B1(n_295), .B2(n_300), .C(n_305), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx4_ASAP7_75t_L g309 ( .A(n_289), .Y(n_309) );
AND2x2_ASAP7_75t_L g403 ( .A(n_289), .B(n_322), .Y(n_403) );
AND2x2_ASAP7_75t_L g410 ( .A(n_289), .B(n_292), .Y(n_410) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_292), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g321 ( .A(n_294), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_297), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g446 ( .A(n_299), .B(n_390), .Y(n_446) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g431 ( .A(n_303), .B(n_359), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_304), .A2(n_397), .B(n_398), .C(n_411), .Y(n_396) );
AOI21xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_310), .B(n_312), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_310), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_408), .Y(n_404) );
AND2x2_ASAP7_75t_L g381 ( .A(n_311), .B(n_322), .Y(n_381) );
AND2x2_ASAP7_75t_L g434 ( .A(n_311), .B(n_329), .Y(n_434) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_314), .B(n_352), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_321), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g362 ( .A(n_317), .B(n_320), .Y(n_362) );
OR2x2_ASAP7_75t_L g405 ( .A(n_317), .B(n_359), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_318), .B(n_384), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_318), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g349 ( .A(n_319), .Y(n_349) );
INVx1_ASAP7_75t_L g415 ( .A(n_322), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_330), .B2(n_331), .Y(n_323) );
INVx1_ASAP7_75t_L g338 ( .A(n_324), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_325), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g401 ( .A(n_326), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g387 ( .A(n_328), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_329), .B(n_415), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_330), .A2(n_389), .B1(n_391), .B2(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g439 ( .A(n_334), .B(n_434), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_335), .A2(n_369), .B1(n_372), .B2(n_373), .C1(n_376), .C2(n_377), .Y(n_368) );
NAND4xp25_ASAP7_75t_SL g336 ( .A(n_337), .B(n_357), .C(n_368), .D(n_380), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B1(n_342), .B2(n_347), .C(n_348), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_340), .B(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_342), .A2(n_412), .B1(n_414), .B2(n_416), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g354 ( .A(n_346), .B(n_355), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_347), .A2(n_409), .B(n_410), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_352), .B2(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B(n_363), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_371), .B(n_390), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_371), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_375), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g407 ( .A(n_379), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_385), .B2(n_387), .C(n_388), .Y(n_380) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_390), .A2(n_428), .B1(n_429), .B2(n_430), .C1(n_432), .C2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_394), .B(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g426 ( .A(n_400), .Y(n_426) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp33_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_440), .B2(n_441), .C(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_451), .A2(n_459), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g748 ( .A(n_462), .Y(n_748) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_656), .C(n_704), .Y(n_463) );
NOR4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_584), .C(n_629), .D(n_643), .Y(n_464) );
OAI311xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_504), .A3(n_528), .B1(n_537), .C1(n_552), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_467), .A2(n_538), .B(n_540), .Y(n_537) );
AND2x2_ASAP7_75t_L g645 ( .A(n_467), .B(n_572), .Y(n_645) );
AND2x2_ASAP7_75t_L g702 ( .A(n_467), .B(n_588), .Y(n_702) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g595 ( .A(n_468), .B(n_498), .Y(n_595) );
AND2x2_ASAP7_75t_L g652 ( .A(n_468), .B(n_600), .Y(n_652) );
INVx1_ASAP7_75t_L g693 ( .A(n_468), .Y(n_693) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_469), .Y(n_561) );
AND2x2_ASAP7_75t_L g602 ( .A(n_469), .B(n_498), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_469), .B(n_499), .Y(n_606) );
INVx1_ASAP7_75t_L g618 ( .A(n_469), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_474), .A2(n_545), .B(n_548), .Y(n_544) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g539 ( .A(n_476), .B(n_498), .Y(n_539) );
INVx2_ASAP7_75t_L g573 ( .A(n_476), .Y(n_573) );
AND2x2_ASAP7_75t_L g588 ( .A(n_476), .B(n_499), .Y(n_588) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_476), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_476), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g608 ( .A(n_476), .B(n_571), .Y(n_608) );
INVx1_ASAP7_75t_L g620 ( .A(n_476), .Y(n_620) );
INVx1_ASAP7_75t_L g661 ( .A(n_476), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_476), .B(n_561), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_481), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g538 ( .A(n_488), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_488), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g623 ( .A(n_488), .B(n_498), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_488), .B(n_618), .Y(n_681) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
OR2x2_ASAP7_75t_L g660 ( .A(n_489), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g567 ( .A(n_499), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_499), .B(n_573), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_502), .A2(n_514), .B(n_516), .C(n_517), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_502), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_504), .B(n_555), .Y(n_718) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g688 ( .A(n_505), .B(n_530), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_519), .Y(n_505) );
AND2x2_ASAP7_75t_L g564 ( .A(n_506), .B(n_555), .Y(n_564) );
INVx2_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
AND2x2_ASAP7_75t_L g610 ( .A(n_506), .B(n_558), .Y(n_610) );
AND2x2_ASAP7_75t_L g677 ( .A(n_506), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_507), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g557 ( .A(n_507), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g597 ( .A(n_507), .B(n_519), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_507), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g540 ( .A(n_519), .B(n_541), .Y(n_540) );
INVx3_ASAP7_75t_L g558 ( .A(n_519), .Y(n_558) );
AND2x2_ASAP7_75t_L g563 ( .A(n_519), .B(n_543), .Y(n_563) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_615), .Y(n_636) );
AND2x2_ASAP7_75t_L g701 ( .A(n_519), .B(n_691), .Y(n_701) );
OAI311xp33_ASAP7_75t_L g584 ( .A1(n_528), .A2(n_585), .A3(n_589), .B1(n_591), .C1(n_611), .Y(n_584) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g596 ( .A(n_529), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g655 ( .A(n_529), .B(n_563), .Y(n_655) );
AND2x2_ASAP7_75t_L g729 ( .A(n_529), .B(n_610), .Y(n_729) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_530), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g664 ( .A(n_530), .Y(n_664) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g555 ( .A(n_531), .Y(n_555) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_531), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g684 ( .A(n_531), .B(n_558), .Y(n_684) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g581 ( .A(n_532), .Y(n_581) );
AND2x2_ASAP7_75t_L g559 ( .A(n_539), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g612 ( .A(n_539), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g692 ( .A(n_539), .B(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_540), .A2(n_572), .B1(n_592), .B2(n_596), .C(n_598), .Y(n_591) );
INVx1_ASAP7_75t_L g716 ( .A(n_541), .Y(n_716) );
OR2x2_ASAP7_75t_L g682 ( .A(n_542), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g577 ( .A(n_543), .B(n_558), .Y(n_577) );
OR2x2_ASAP7_75t_L g579 ( .A(n_543), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g604 ( .A(n_543), .Y(n_604) );
INVx2_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
AND2x2_ASAP7_75t_L g642 ( .A(n_543), .B(n_580), .Y(n_642) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_543), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_559), .B1(n_562), .B2(n_565), .C(n_568), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g653 ( .A(n_555), .B(n_563), .Y(n_653) );
AND2x2_ASAP7_75t_L g703 ( .A(n_555), .B(n_557), .Y(n_703) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g590 ( .A(n_557), .B(n_561), .Y(n_590) );
AND2x2_ASAP7_75t_L g669 ( .A(n_557), .B(n_642), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_558), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g628 ( .A(n_558), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_559), .A2(n_639), .B(n_641), .Y(n_638) );
OR2x2_ASAP7_75t_L g582 ( .A(n_560), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g648 ( .A(n_560), .B(n_608), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_560), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g625 ( .A(n_561), .B(n_594), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_561), .B(n_708), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_562), .B(n_588), .Y(n_698) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_576), .Y(n_621) );
INVx1_ASAP7_75t_L g637 ( .A(n_564), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_574), .B1(n_578), .B2(n_582), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g600 ( .A(n_571), .Y(n_600) );
INVx1_ASAP7_75t_L g613 ( .A(n_571), .Y(n_613) );
INVx1_ASAP7_75t_L g583 ( .A(n_572), .Y(n_583) );
AND2x2_ASAP7_75t_L g654 ( .A(n_572), .B(n_600), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_572), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
OR2x2_ASAP7_75t_L g578 ( .A(n_575), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_575), .B(n_691), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_575), .B(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g725 ( .A(n_577), .B(n_677), .Y(n_725) );
INVx1_ASAP7_75t_SL g691 ( .A(n_579), .Y(n_691) );
AND2x2_ASAP7_75t_L g631 ( .A(n_580), .B(n_615), .Y(n_631) );
INVx1_ASAP7_75t_L g678 ( .A(n_580), .Y(n_678) );
OAI222xp33_ASAP7_75t_L g719 ( .A1(n_585), .A2(n_675), .B1(n_720), .B2(n_721), .C1(n_724), .C2(n_726), .Y(n_719) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g640 ( .A(n_587), .Y(n_640) );
AND2x2_ASAP7_75t_L g651 ( .A(n_588), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_588), .B(n_693), .Y(n_720) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_590), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g695 ( .A(n_592), .Y(n_695) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g633 ( .A(n_595), .Y(n_633) );
AND2x2_ASAP7_75t_L g712 ( .A(n_595), .B(n_673), .Y(n_712) );
AND2x2_ASAP7_75t_L g735 ( .A(n_595), .B(n_619), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_597), .B(n_631), .Y(n_630) );
OAI32xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .A3(n_603), .B1(n_605), .B2(n_609), .Y(n_598) );
BUFx2_ASAP7_75t_L g673 ( .A(n_600), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_601), .B(n_619), .Y(n_700) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g639 ( .A(n_602), .B(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g707 ( .A(n_602), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g696 ( .A(n_603), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g667 ( .A(n_606), .B(n_640), .Y(n_667) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g629 ( .A1(n_608), .A2(n_630), .B1(n_632), .B2(n_634), .C(n_638), .Y(n_629) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g641 ( .A(n_610), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_631), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B1(n_616), .B2(n_621), .C(n_622), .Y(n_611) );
INVx1_ASAP7_75t_L g730 ( .A(n_612), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_613), .B(n_707), .Y(n_706) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_614), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_619), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g685 ( .A(n_619), .Y(n_685) );
BUFx3_ASAP7_75t_L g708 ( .A(n_620), .Y(n_708) );
INVx1_ASAP7_75t_SL g649 ( .A(n_621), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_621), .B(n_663), .Y(n_662) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B(n_626), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_623), .A2(n_724), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_727) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g670 ( .A(n_628), .B(n_631), .Y(n_670) );
INVx1_ASAP7_75t_L g734 ( .A(n_628), .Y(n_734) );
INVx2_ASAP7_75t_L g723 ( .A(n_631), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_631), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g676 ( .A(n_636), .B(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_646), .B1(n_648), .B2(n_649), .C(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_652), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_655), .A2(n_732), .B(n_735), .Y(n_731) );
NOR4xp25_ASAP7_75t_SL g656 ( .A(n_657), .B(n_665), .C(n_674), .D(n_694), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B1(n_671), .B2(n_672), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B1(n_682), .B2(n_685), .C(n_686), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g697 ( .A(n_677), .Y(n_697) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_689), .B(n_692), .Y(n_686) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .C(n_699), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_699) );
CKINVDCx14_ASAP7_75t_R g709 ( .A(n_703), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_719), .C(n_727), .Y(n_704) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B1(n_710), .B2(n_711), .C(n_713), .Y(n_705) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g747 ( .A(n_737), .Y(n_747) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_740), .Y(n_749) );
INVx1_ASAP7_75t_L g744 ( .A(n_741), .Y(n_744) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
endmodule