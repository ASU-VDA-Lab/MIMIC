module fake_jpeg_24842_n_140 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_39),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_19),
.A2(n_1),
.B(n_2),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_17),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_32),
.B(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_54),
.B1(n_28),
.B2(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_20),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_15),
.B1(n_23),
.B2(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_61),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.C(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_48),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_35),
.B(n_26),
.C(n_23),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_14),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_15),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_47),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_85),
.B(n_88),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_44),
.B1(n_41),
.B2(n_37),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_68),
.B1(n_44),
.B2(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_46),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_64),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_85),
.C(n_78),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_61),
.B(n_22),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_97),
.B(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_61),
.B1(n_63),
.B2(n_69),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_57),
.B(n_25),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_75),
.C(n_78),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_110),
.C(n_111),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_82),
.C(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_95),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_117),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_97),
.B(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_93),
.B1(n_97),
.B2(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_120),
.B1(n_106),
.B2(n_111),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_66),
.B1(n_73),
.B2(n_86),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_86),
.B(n_14),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_127),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_109),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_6),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_14),
.C(n_16),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.C(n_116),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_114),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_132),
.B(n_125),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_8),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_9),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_136),
.B(n_9),
.Y(n_138)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_138),
.A3(n_11),
.B1(n_12),
.B2(n_134),
.C(n_85),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_11),
.Y(n_140)
);


endmodule