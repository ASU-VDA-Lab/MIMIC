module real_jpeg_268_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_12),
.C(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_1),
.A2(n_20),
.B1(n_44),
.B2(n_50),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_3),
.A2(n_12),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_18),
.B1(n_44),
.B2(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_4),
.A2(n_12),
.B1(n_19),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_12),
.B1(n_19),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_33),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_23),
.B(n_32),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_16),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_14),
.Y(n_11)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_22),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_16)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_27),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_49),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_31),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_54),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_41),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);


endmodule