module fake_jpeg_712_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_12),
.B1(n_15),
.B2(n_23),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_35),
.B1(n_26),
.B2(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_43),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_20),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_48),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_28),
.B(n_29),
.C(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_13),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_44),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_39),
.B1(n_31),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_64),
.C(n_67),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_54),
.C(n_47),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_49),
.B1(n_11),
.B2(n_28),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_66),
.B1(n_58),
.B2(n_62),
.C(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_71),
.B(n_76),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_82),
.B(n_1),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_60),
.B1(n_73),
.B2(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_89),
.B1(n_0),
.B2(n_1),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_82),
.B(n_81),
.C(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_2),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_6),
.C(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_95),
.C(n_10),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.C(n_10),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_2),
.Y(n_101)
);


endmodule