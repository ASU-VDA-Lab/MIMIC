module fake_ariane_2886_n_23 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_23);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_23;

wire n_22;
wire n_13;
wire n_20;
wire n_17;
wire n_18;
wire n_11;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_10;

INVx4_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

OAI21xp33_ASAP7_75t_L g11 ( 
.A1(n_7),
.A2(n_3),
.B(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_2),
.B(n_4),
.Y(n_12)
);

OAI22xp33_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_3),
.B1(n_8),
.B2(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

OAI21x1_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_11),
.B(n_10),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_14),
.B(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_14),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_16),
.B1(n_17),
.B2(n_13),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_0),
.C(n_2),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_17),
.C(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_21),
.Y(n_23)
);


endmodule