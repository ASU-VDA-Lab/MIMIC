module fake_jpeg_18851_n_292 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_292);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_20),
.Y(n_38)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_51),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_32),
.C(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_30),
.B(n_29),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_61),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_28),
.B(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_28),
.B1(n_27),
.B2(n_35),
.Y(n_71)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_65),
.B1(n_41),
.B2(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_66),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_46),
.B1(n_40),
.B2(n_47),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_78),
.B1(n_57),
.B2(n_54),
.Y(n_91)
);

AO22x2_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_28),
.B1(n_47),
.B2(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_71),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_47),
.B1(n_28),
.B2(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_54),
.B1(n_50),
.B2(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_34),
.B1(n_41),
.B2(n_15),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_17),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_42),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_69),
.B1(n_73),
.B2(n_80),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_71),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_69),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_53),
.B1(n_57),
.B2(n_48),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_67),
.B1(n_69),
.B2(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_73),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_65),
.B1(n_62),
.B2(n_16),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_16),
.B1(n_15),
.B2(n_24),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_43),
.B1(n_84),
.B2(n_15),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_42),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_83),
.B1(n_81),
.B2(n_74),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_120),
.B1(n_121),
.B2(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_68),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_85),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_116),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_117),
.B(n_126),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_69),
.B(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_125),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_42),
.C(n_80),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_112),
.C(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_73),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_13),
.B1(n_52),
.B2(n_25),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_141),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_89),
.B(n_92),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_140),
.B(n_114),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_91),
.B1(n_99),
.B2(n_104),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_120),
.B1(n_133),
.B2(n_153),
.Y(n_168)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_94),
.B(n_25),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_94),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_153),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_76),
.A3(n_97),
.B1(n_43),
.B2(n_31),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_124),
.B(n_127),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_31),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_97),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_76),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_52),
.C(n_32),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_123),
.C(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_52),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_126),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_115),
.C(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_170),
.C(n_175),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_182),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_114),
.C(n_109),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_52),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_52),
.C(n_32),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_180),
.C(n_181),
.Y(n_194)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_146),
.B1(n_136),
.B2(n_144),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_64),
.C(n_39),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_23),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_23),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_11),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_170),
.B1(n_173),
.B2(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_174),
.A2(n_138),
.B1(n_155),
.B2(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_205),
.B1(n_181),
.B2(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_23),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_142),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_171),
.A2(n_136),
.B1(n_142),
.B2(n_13),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_163),
.C(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_198),
.C(n_194),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_213),
.B1(n_205),
.B2(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_158),
.B1(n_13),
.B2(n_17),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_25),
.B1(n_21),
.B2(n_18),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_49),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_21),
.B(n_18),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_213),
.B(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_49),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_186),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_188),
.B(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_198),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_192),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_64),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_195),
.C(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_202),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_215),
.B(n_217),
.C(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_208),
.B1(n_215),
.B2(n_217),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_249),
.C(n_19),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_219),
.A3(n_220),
.B1(n_206),
.B2(n_191),
.C1(n_221),
.C2(n_214),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_19),
.C(n_33),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_64),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_33),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_237),
.C(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_262),
.C(n_249),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_228),
.B(n_1),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_64),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_0),
.B(n_2),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_19),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_263),
.B1(n_252),
.B2(n_4),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_19),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_2),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_245),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_3),
.B(n_4),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_270),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_272),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_7),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_274),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_7),
.B(n_8),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_274),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_268),
.C(n_269),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_285),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_265),
.C(n_279),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_10),
.C(n_7),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_290),
.B(n_9),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_9),
.C(n_10),
.Y(n_292)
);


endmodule