module fake_jpeg_5573_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_1),
.Y(n_6)
);

BUFx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_16),
.B1(n_8),
.B2(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

OR2x2_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_9),
.B1(n_11),
.B2(n_8),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_19),
.B1(n_14),
.B2(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_6),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_17),
.B1(n_12),
.B2(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_28),
.B1(n_10),
.B2(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_13),
.B1(n_8),
.B2(n_6),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_10),
.C(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_27),
.C(n_30),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_33),
.Y(n_37)
);

AOI221xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.C(n_3),
.Y(n_36)
);

NAND5xp2_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_29),
.C(n_1),
.D(n_2),
.E(n_3),
.Y(n_38)
);

OAI31xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_0),
.A3(n_2),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_3),
.Y(n_40)
);


endmodule