module fake_jpeg_25837_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_50),
.B1(n_30),
.B2(n_29),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_29),
.B1(n_27),
.B2(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_28),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_51),
.B(n_59),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_44),
.B(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_78)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_71),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_17),
.B1(n_31),
.B2(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_87),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_58),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_94),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_45),
.B(n_58),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_86),
.B(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_53),
.B1(n_55),
.B2(n_46),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_91),
.B1(n_92),
.B2(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_75),
.B1(n_63),
.B2(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_53),
.B1(n_48),
.B2(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_63),
.C(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_11),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_94),
.B(n_78),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_66),
.B1(n_53),
.B2(n_48),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_93),
.B1(n_87),
.B2(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_81),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_105),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_100),
.C(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.C(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_100),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_103),
.C(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_135),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_82),
.C(n_89),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_113),
.C(n_1),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_10),
.CI(n_9),
.CON(n_135),
.SN(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_115),
.B1(n_123),
.B2(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_144),
.B(n_145),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_121),
.A3(n_118),
.B1(n_114),
.B2(n_116),
.C1(n_113),
.C2(n_117),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_127),
.B(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_119),
.B1(n_134),
.B2(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_133),
.C(n_132),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_126),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_135),
.B(n_2),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_138),
.B1(n_146),
.B2(n_3),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_10),
.C(n_8),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_3),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_0),
.C(n_2),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_7),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_155),
.B(n_4),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_149),
.B1(n_152),
.B2(n_5),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_7),
.B(n_156),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_160),
.C(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_164),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_167),
.Y(n_169)
);


endmodule