module fake_jpeg_25407_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_23),
.Y(n_48)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_27),
.B1(n_34),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_16),
.B1(n_28),
.B2(n_29),
.Y(n_76)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx11_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_86),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_41),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_73),
.B1(n_16),
.B2(n_28),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_27),
.B1(n_23),
.B2(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_78),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_87),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_84)
);

CKINVDCx6p67_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_20),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_50),
.B1(n_67),
.B2(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_92),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_33),
.B1(n_18),
.B2(n_34),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_18),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_43),
.A3(n_39),
.B1(n_31),
.B2(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_108),
.B1(n_117),
.B2(n_95),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_47),
.C(n_62),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_104),
.C(n_71),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_120),
.B1(n_90),
.B2(n_88),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_109),
.Y(n_133)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_66),
.B1(n_95),
.B2(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_47),
.C(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_50),
.B1(n_47),
.B2(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_29),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_65),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_81),
.B1(n_73),
.B2(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_121),
.B1(n_79),
.B2(n_92),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_54),
.B1(n_49),
.B2(n_21),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_49),
.B1(n_21),
.B2(n_19),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_132),
.B1(n_151),
.B2(n_107),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_149),
.B1(n_59),
.B2(n_2),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_139),
.C(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_130),
.B(n_131),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_87),
.B1(n_71),
.B2(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_80),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_89),
.B1(n_66),
.B2(n_33),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_80),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_145),
.B(n_152),
.Y(n_155)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_150),
.Y(n_177)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_85),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_77),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_94),
.B1(n_19),
.B2(n_49),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_49),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_0),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_59),
.C(n_8),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_8),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_106),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_164),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_107),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_163),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_161),
.B(n_165),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_107),
.B(n_123),
.C(n_117),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_168),
.Y(n_193)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_135),
.B1(n_127),
.B2(n_129),
.Y(n_189)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_179),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_107),
.B1(n_100),
.B2(n_116),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_181),
.B1(n_9),
.B2(n_14),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_123),
.B1(n_99),
.B2(n_115),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_99),
.B(n_1),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_0),
.B(n_2),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_153),
.B1(n_133),
.B2(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_187),
.Y(n_209)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_7),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_176),
.B1(n_171),
.B2(n_187),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_152),
.B1(n_132),
.B2(n_126),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_202),
.B1(n_208),
.B2(n_165),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_139),
.C(n_152),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_204),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_201),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_186),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_180),
.B1(n_184),
.B2(n_157),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_11),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_213),
.B(n_161),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_158),
.A2(n_3),
.B(n_4),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_182),
.B(n_210),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_229),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_218),
.A2(n_231),
.B(n_233),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_155),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_234),
.B1(n_237),
.B2(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_159),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_202),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_160),
.B1(n_158),
.B2(n_168),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_177),
.B(n_157),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_239),
.B(n_207),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_177),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_213),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_203),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_215),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_195),
.C(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_256),
.C(n_218),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_208),
.Y(n_249)
);

OA21x2_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_216),
.B(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_228),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_206),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_230),
.C(n_238),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_239),
.B1(n_234),
.B2(n_231),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_211),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_236),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_245),
.B(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_273),
.B1(n_259),
.B2(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_223),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_195),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_167),
.C(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_167),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_214),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_214),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_198),
.B1(n_203),
.B2(n_163),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_258),
.B1(n_253),
.B2(n_256),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_286),
.B1(n_4),
.B2(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_243),
.CI(n_249),
.CON(n_278),
.SN(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_261),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_252),
.B(n_244),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_285),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_198),
.B(n_241),
.Y(n_284)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_15),
.C(n_287),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_166),
.B(n_242),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_166),
.B1(n_172),
.B2(n_170),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_267),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_297),
.B(n_285),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_261),
.C(n_11),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_281),
.C(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_277),
.B(n_15),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_277),
.B(n_4),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_286),
.A3(n_282),
.B1(n_275),
.B2(n_278),
.C1(n_279),
.C2(n_287),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_295),
.B(n_291),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_R g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_308),
.B(n_311),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_292),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_309),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_312),
.B(n_300),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_304),
.B(n_278),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_302),
.Y(n_317)
);


endmodule