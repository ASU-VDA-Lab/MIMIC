module real_aes_8602_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_668;
wire n_237;
wire n_429;
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_0), .A2(n_192), .B1(n_569), .B2(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_1), .B(n_278), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_2), .A2(n_15), .B1(n_455), .B2(n_636), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_3), .A2(n_112), .B1(n_488), .B2(n_489), .C(n_491), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_4), .A2(n_127), .B1(n_453), .B2(n_578), .Y(n_616) );
XOR2x2_ASAP7_75t_L g530 ( .A(n_5), .B(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_6), .A2(n_18), .B1(n_418), .B2(n_420), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_7), .A2(n_140), .B1(n_313), .B2(n_376), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_8), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_9), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_10), .A2(n_95), .B1(n_122), .B2(n_344), .C1(n_449), .C2(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_11), .A2(n_104), .B1(n_251), .B2(n_422), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_12), .A2(n_108), .B1(n_364), .B2(n_557), .Y(n_556) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_13), .A2(n_392), .B1(n_393), .B2(n_431), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_13), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_14), .A2(n_147), .B1(n_293), .B2(n_422), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_16), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_17), .A2(n_179), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_19), .A2(n_198), .B1(n_262), .B2(n_267), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_20), .Y(n_515) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_21), .A2(n_62), .B1(n_230), .B2(n_235), .Y(n_239) );
INVx1_ASAP7_75t_L g656 ( .A(n_21), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_22), .A2(n_182), .B1(n_313), .B2(n_315), .C(n_317), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_23), .A2(n_26), .B1(n_345), .B2(n_369), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_24), .A2(n_44), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_25), .A2(n_79), .B1(n_120), .B2(n_341), .C1(n_342), .C2(n_344), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_27), .Y(n_309) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_28), .A2(n_97), .B1(n_153), .B2(n_554), .C1(n_638), .C2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_29), .A2(n_199), .B1(n_282), .B2(n_449), .Y(n_448) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_30), .A2(n_64), .B1(n_230), .B2(n_231), .Y(n_237) );
INVx1_ASAP7_75t_L g657 ( .A(n_30), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_31), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_32), .A2(n_91), .B1(n_419), .B2(n_453), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_33), .A2(n_149), .B1(n_477), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_34), .A2(n_77), .B1(n_420), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_35), .A2(n_206), .B1(n_311), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_36), .A2(n_57), .B1(n_563), .B2(n_565), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_37), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_38), .A2(n_184), .B1(n_519), .B2(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_39), .A2(n_549), .B1(n_550), .B2(n_581), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_39), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_40), .A2(n_103), .B1(n_267), .B2(n_282), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_41), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_42), .A2(n_187), .B1(n_428), .B2(n_525), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_43), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_45), .A2(n_99), .B1(n_385), .B2(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_46), .A2(n_148), .B1(n_291), .B2(n_293), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_47), .A2(n_107), .B1(n_299), .B2(n_301), .C(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_48), .B(n_272), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_49), .A2(n_88), .B1(n_419), .B2(n_521), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_50), .A2(n_109), .B1(n_327), .B2(n_329), .C(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g545 ( .A(n_51), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_52), .A2(n_173), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_53), .A2(n_119), .B1(n_246), .B2(n_251), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_54), .A2(n_195), .B1(n_263), .B2(n_343), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_55), .A2(n_461), .B1(n_496), .B2(n_497), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_55), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_56), .A2(n_297), .B1(n_346), .B2(n_347), .Y(n_296) );
INVx1_ASAP7_75t_L g346 ( .A(n_56), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_58), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_59), .A2(n_163), .B1(n_268), .B2(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_60), .A2(n_96), .B1(n_311), .B2(n_388), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_61), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_63), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_65), .A2(n_165), .B1(n_293), .B2(n_383), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_66), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_67), .A2(n_138), .B1(n_299), .B2(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g214 ( .A(n_68), .B(n_215), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_69), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_70), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_71), .A2(n_146), .B1(n_246), .B2(n_251), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_72), .A2(n_170), .B1(n_361), .B2(n_404), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_73), .A2(n_106), .B1(n_345), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g211 ( .A(n_74), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_75), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_76), .A2(n_87), .B1(n_624), .B2(n_625), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_78), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_80), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_81), .A2(n_126), .B1(n_272), .B2(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_82), .A2(n_102), .B1(n_368), .B2(n_369), .Y(n_367) );
OA22x2_ASAP7_75t_L g499 ( .A1(n_83), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_83), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_84), .A2(n_85), .B1(n_572), .B2(n_574), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_86), .A2(n_101), .B1(n_282), .B2(n_343), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_89), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_90), .A2(n_123), .B1(n_422), .B2(n_627), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_92), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_93), .A2(n_169), .B1(n_226), .B2(n_240), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_94), .A2(n_137), .B1(n_385), .B2(n_387), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_98), .A2(n_171), .B1(n_374), .B2(n_375), .Y(n_373) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_100), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g215 ( .A(n_105), .Y(n_215) );
INVx1_ASAP7_75t_L g688 ( .A(n_110), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_111), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_113), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_114), .B(n_328), .Y(n_446) );
AND2x6_ASAP7_75t_L g210 ( .A(n_115), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_115), .Y(n_650) );
AO22x2_ASAP7_75t_L g229 ( .A1(n_116), .A2(n_175), .B1(n_230), .B2(n_231), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_117), .A2(n_161), .B1(n_313), .B2(n_422), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_118), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_121), .A2(n_193), .B1(n_262), .B2(n_267), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_124), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_125), .A2(n_183), .B1(n_303), .B2(n_311), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_128), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_129), .A2(n_168), .B1(n_280), .B2(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_130), .B(n_488), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_131), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_132), .B(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_133), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_134), .A2(n_143), .B1(n_374), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_135), .A2(n_205), .B1(n_328), .B2(n_329), .Y(n_540) );
AO22x2_ASAP7_75t_L g234 ( .A1(n_136), .A2(n_186), .B1(n_230), .B2(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_139), .A2(n_203), .B1(n_291), .B2(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_141), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_142), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_144), .A2(n_194), .B1(n_521), .B2(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_145), .B(n_371), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_150), .A2(n_174), .B1(n_291), .B2(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_151), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_152), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_154), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_155), .A2(n_159), .B1(n_378), .B2(n_380), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_156), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_157), .A2(n_201), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_158), .A2(n_160), .B1(n_525), .B2(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_162), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_164), .B(n_278), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_166), .Y(n_478) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_167), .A2(n_208), .B(n_216), .C(n_658), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_172), .A2(n_660), .B1(n_661), .B2(n_679), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_172), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_175), .B(n_655), .Y(n_654) );
OA22x2_ASAP7_75t_L g353 ( .A1(n_176), .A2(n_354), .B1(n_355), .B2(n_389), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_176), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_177), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_178), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_180), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_181), .A2(n_204), .B1(n_287), .B2(n_288), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_185), .Y(n_257) );
INVx1_ASAP7_75t_L g653 ( .A(n_186), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_188), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_189), .B(n_511), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_190), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_191), .B(n_488), .Y(n_630) );
INVx1_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_197), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_200), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_202), .Y(n_359) );
INVx1_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_211), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_212), .A2(n_648), .B(n_687), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_528), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_216) );
INVxp67_ASAP7_75t_L g643 ( .A(n_217), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B1(n_433), .B2(n_527), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AOI22xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B1(n_350), .B2(n_432), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_296), .B1(n_348), .B2(n_349), .Y(n_221) );
INVx3_ASAP7_75t_L g348 ( .A(n_222), .Y(n_348) );
XOR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_295), .Y(n_222) );
NAND3x1_ASAP7_75t_SL g223 ( .A(n_224), .B(n_255), .C(n_285), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_245), .Y(n_224) );
INVx6_ASAP7_75t_L g314 ( .A(n_226), .Y(n_314) );
BUFx3_ASAP7_75t_L g374 ( .A(n_226), .Y(n_374) );
BUFx3_ASAP7_75t_L g453 ( .A(n_226), .Y(n_453) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
AND2x6_ASAP7_75t_L g259 ( .A(n_227), .B(n_260), .Y(n_259) );
AND2x6_ASAP7_75t_L g287 ( .A(n_227), .B(n_275), .Y(n_287) );
AND2x2_ASAP7_75t_L g292 ( .A(n_227), .B(n_248), .Y(n_292) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_233), .Y(n_227) );
AND2x2_ASAP7_75t_L g250 ( .A(n_228), .B(n_234), .Y(n_250) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g243 ( .A(n_229), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_229), .B(n_234), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_229), .B(n_239), .Y(n_266) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g235 ( .A(n_232), .Y(n_235) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g244 ( .A(n_234), .Y(n_244) );
INVx1_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
AND2x2_ASAP7_75t_L g242 ( .A(n_236), .B(n_243), .Y(n_242) );
AND2x6_ASAP7_75t_L g278 ( .A(n_236), .B(n_250), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_236), .B(n_243), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_236), .B(n_250), .Y(n_415) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g249 ( .A(n_237), .Y(n_249) );
AND2x2_ASAP7_75t_L g260 ( .A(n_237), .B(n_239), .Y(n_260) );
OR2x2_ASAP7_75t_L g276 ( .A(n_237), .B(n_238), .Y(n_276) );
INVx1_ASAP7_75t_L g284 ( .A(n_237), .Y(n_284) );
AND2x2_ASAP7_75t_L g248 ( .A(n_238), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_240), .Y(n_612) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g379 ( .A(n_241), .Y(n_379) );
INVx5_ASAP7_75t_L g419 ( .A(n_241), .Y(n_419) );
INVx3_ASAP7_75t_L g455 ( .A(n_241), .Y(n_455) );
INVx2_ASAP7_75t_L g535 ( .A(n_241), .Y(n_535) );
BUFx3_ASAP7_75t_L g573 ( .A(n_241), .Y(n_573) );
INVx8_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g289 ( .A(n_243), .B(n_248), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_243), .B(n_248), .Y(n_486) );
INVx1_ASAP7_75t_L g269 ( .A(n_244), .Y(n_269) );
INVx4_ASAP7_75t_L g316 ( .A(n_246), .Y(n_316) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx3_ASAP7_75t_L g388 ( .A(n_247), .Y(n_388) );
INVx2_ASAP7_75t_L g430 ( .A(n_247), .Y(n_430) );
BUFx3_ASAP7_75t_L g440 ( .A(n_247), .Y(n_440) );
BUFx3_ASAP7_75t_L g519 ( .A(n_247), .Y(n_519) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND2x4_ASAP7_75t_L g294 ( .A(n_248), .B(n_253), .Y(n_294) );
INVx1_ASAP7_75t_L g252 ( .A(n_249), .Y(n_252) );
AND2x2_ASAP7_75t_L g281 ( .A(n_249), .B(n_265), .Y(n_281) );
AND2x4_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g411 ( .A(n_250), .Y(n_411) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_252), .B(n_266), .Y(n_334) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x6_ASAP7_75t_L g325 ( .A(n_254), .B(n_284), .Y(n_325) );
NOR2x1_ASAP7_75t_L g255 ( .A(n_256), .B(n_270), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_261), .Y(n_256) );
INVx4_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
BUFx2_ASAP7_75t_L g358 ( .A(n_258), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_258), .A2(n_443), .B(n_444), .Y(n_442) );
INVx4_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g402 ( .A(n_259), .Y(n_402) );
BUFx3_ASAP7_75t_L g513 ( .A(n_259), .Y(n_513) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_259), .Y(n_554) );
AND2x4_ASAP7_75t_L g268 ( .A(n_260), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
BUFx4f_ASAP7_75t_L g364 ( .A(n_262), .Y(n_364) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx12f_ASAP7_75t_L g345 ( .A(n_263), .Y(n_345) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_263), .Y(n_406) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g280 ( .A(n_266), .B(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g282 ( .A(n_266), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g566 ( .A(n_267), .Y(n_566) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g369 ( .A(n_268), .Y(n_369) );
INVx1_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .C(n_279), .Y(n_270) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_272), .Y(n_488) );
INVx5_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g328 ( .A(n_273), .Y(n_328) );
INVx2_ASAP7_75t_L g668 ( .A(n_273), .Y(n_668) );
INVx4_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g410 ( .A(n_276), .B(n_411), .Y(n_410) );
BUFx4f_ASAP7_75t_L g329 ( .A(n_278), .Y(n_329) );
BUFx2_ASAP7_75t_L g371 ( .A(n_278), .Y(n_371) );
INVx1_ASAP7_75t_SL g490 ( .A(n_278), .Y(n_490) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_280), .Y(n_361) );
BUFx4f_ASAP7_75t_SL g449 ( .A(n_280), .Y(n_449) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_280), .Y(n_511) );
BUFx2_ASAP7_75t_L g368 ( .A(n_282), .Y(n_368) );
BUFx3_ASAP7_75t_L g542 ( .A(n_282), .Y(n_542) );
INVx1_ASAP7_75t_L g564 ( .A(n_282), .Y(n_564) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
INVx11_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
INVx11_ASAP7_75t_L g425 ( .A(n_287), .Y(n_425) );
BUFx4f_ASAP7_75t_SL g578 ( .A(n_288), .Y(n_578) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
BUFx3_ASAP7_75t_L g376 ( .A(n_289), .Y(n_376) );
BUFx3_ASAP7_75t_L g422 ( .A(n_289), .Y(n_422) );
INVx3_ASAP7_75t_L g300 ( .A(n_291), .Y(n_300) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_291), .Y(n_577) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g386 ( .A(n_292), .Y(n_386) );
BUFx2_ASAP7_75t_SL g428 ( .A(n_292), .Y(n_428) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
BUFx2_ASAP7_75t_SL g426 ( .A(n_294), .Y(n_426) );
BUFx3_ASAP7_75t_L g468 ( .A(n_294), .Y(n_468) );
BUFx2_ASAP7_75t_L g570 ( .A(n_294), .Y(n_570) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_294), .Y(n_610) );
BUFx3_ASAP7_75t_L g625 ( .A(n_294), .Y(n_625) );
INVx1_ASAP7_75t_L g349 ( .A(n_296), .Y(n_349) );
INVx1_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
AND4x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_312), .C(n_326), .D(n_340), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_309), .B2(n_310), .Y(n_304) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
INVx2_ASAP7_75t_SL g452 ( .A(n_308), .Y(n_452) );
INVx2_ASAP7_75t_L g624 ( .A(n_308), .Y(n_624) );
INVx5_ASAP7_75t_SL g675 ( .A(n_308), .Y(n_675) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g479 ( .A(n_313), .Y(n_479) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g580 ( .A(n_314), .Y(n_580) );
INVx3_ASAP7_75t_L g634 ( .A(n_314), .Y(n_634) );
INVx4_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g569 ( .A(n_316), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_322), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_319), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_469) );
BUFx2_ASAP7_75t_R g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx2_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
BUFx2_ASAP7_75t_L g521 ( .A(n_324), .Y(n_521) );
BUFx2_ASAP7_75t_L g636 ( .A(n_324), .Y(n_636) );
INVx6_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g420 ( .A(n_325), .Y(n_420) );
INVx1_ASAP7_75t_SL g574 ( .A(n_325), .Y(n_574) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_335), .B2(n_336), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_332), .A2(n_336), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_334), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_334), .A2(n_337), .B1(n_515), .B2(n_516), .Y(n_514) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_334), .Y(n_604) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_337), .Y(n_399) );
OR2x6_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx4f_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g640 ( .A(n_345), .Y(n_640) );
INVx1_ASAP7_75t_L g432 ( .A(n_350), .Y(n_432) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_390), .B2(n_391), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_372), .C(n_381), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_366), .Y(n_356) );
OAI222xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_360), .B2(n_362), .C1(n_363), .C2(n_365), .Y(n_357) );
INVx1_ASAP7_75t_L g495 ( .A(n_358), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g472 ( .A(n_380), .Y(n_472) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g627 ( .A(n_386), .Y(n_627) );
INVx1_ASAP7_75t_L g465 ( .A(n_387), .Y(n_465) );
BUFx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_416), .Y(n_393) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_395), .B(n_400), .C(n_407), .Y(n_394) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g606 ( .A(n_399), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_403), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_402), .A2(n_597), .B1(n_598), .B2(n_600), .C(n_601), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_402), .A2(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g599 ( .A(n_406), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_412), .B2(n_413), .Y(n_407) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g506 ( .A(n_410), .Y(n_506) );
INVx2_ASAP7_75t_L g592 ( .A(n_410), .Y(n_592) );
OA211x2_ASAP7_75t_L g628 ( .A1(n_413), .A2(n_629), .B(n_630), .C(n_631), .Y(n_628) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g508 ( .A(n_415), .Y(n_508) );
AND4x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_421), .C(n_423), .D(n_427), .Y(n_416) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx4_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_SL g477 ( .A(n_425), .Y(n_477) );
INVx4_ASAP7_75t_L g525 ( .A(n_425), .Y(n_525) );
INVx1_ASAP7_75t_L g482 ( .A(n_428), .Y(n_482) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_457), .B1(n_458), .B2(n_526), .Y(n_433) );
INVx1_ASAP7_75t_L g526 ( .A(n_434), .Y(n_526) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
XOR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_456), .Y(n_435) );
NAND3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .C(n_450), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
BUFx2_ASAP7_75t_L g615 ( .A(n_440), .Y(n_615) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .C(n_448), .Y(n_445) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_498), .B2(n_499), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g497 ( .A(n_461), .Y(n_497) );
AND4x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .C(n_487), .D(n_494), .Y(n_461) );
NOR2xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_469), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_463) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_480), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_478), .B2(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND3x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_517), .C(n_522), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .C(n_514), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_504) );
INVx2_ASAP7_75t_L g595 ( .A(n_508), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
INVx4_ASAP7_75t_L g558 ( .A(n_511), .Y(n_558) );
BUFx2_ASAP7_75t_L g638 ( .A(n_511), .Y(n_638) );
INVx3_ASAP7_75t_L g544 ( .A(n_513), .Y(n_544) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_528), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_583), .B1(n_584), .B2(n_642), .Y(n_528) );
INVx1_ASAP7_75t_L g642 ( .A(n_529), .Y(n_642) );
AO22x1_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_547), .B1(n_548), .B2(n_582), .Y(n_529) );
INVx1_ASAP7_75t_SL g582 ( .A(n_530), .Y(n_582) );
NOR4xp75_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .C(n_539), .D(n_543), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
NAND3x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_567), .C(n_575), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_559), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_555), .B(n_556), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .C(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B1(n_617), .B2(n_618), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_607), .Y(n_587) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_596), .C(n_602), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_594), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_613), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_641), .Y(n_620) );
NAND4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_628), .C(n_632), .D(n_637), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
OR2x2_ASAP7_75t_SL g692 ( .A(n_647), .B(n_652), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_648), .Y(n_681) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_649), .B(n_684), .Y(n_687) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_650), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OAI322xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_680), .A3(n_682), .B1(n_685), .B2(n_688), .C1(n_689), .C2(n_692), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
XOR2x2_ASAP7_75t_L g691 ( .A(n_661), .B(n_688), .Y(n_691) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_662), .B(n_671), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .C(n_670), .Y(n_666) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g685 ( .A(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
endmodule