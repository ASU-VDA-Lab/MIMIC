module fake_jpeg_9561_n_46 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_10),
.B1(n_1),
.B2(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_36),
.B1(n_30),
.B2(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_11),
.CI(n_15),
.CON(n_37),
.SN(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI31xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_41),
.A3(n_28),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_17),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_18),
.C(n_22),
.Y(n_46)
);


endmodule