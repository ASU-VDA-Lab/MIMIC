module fake_jpeg_13760_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_0),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_55),
.B1(n_49),
.B2(n_59),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_55),
.B1(n_59),
.B2(n_54),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_95),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_46),
.B(n_80),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_53),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_60),
.B1(n_50),
.B2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_2),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_122),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_80),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_121),
.B1(n_16),
.B2(n_17),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_14),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_124),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_31),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_8),
.B(n_12),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_131),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_18),
.B(n_19),
.C(n_21),
.D(n_22),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_26),
.C(n_27),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_29),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_128),
.C(n_106),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_129),
.B1(n_133),
.B2(n_114),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_144),
.A2(n_145),
.B1(n_140),
.B2(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_146),
.A2(n_147),
.B(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_118),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_118),
.B(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_138),
.C(n_39),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_37),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_113),
.B(n_107),
.Y(n_154)
);


endmodule