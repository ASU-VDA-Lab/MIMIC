module real_jpeg_22273_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_0),
.B(n_75),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_0),
.A2(n_14),
.B(n_34),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_0),
.A2(n_59),
.B1(n_121),
.B2(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_0),
.B(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_0),
.B(n_46),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_0),
.A2(n_46),
.B(n_230),
.Y(n_234)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_73),
.B1(n_78),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_129),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_5),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_29),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_7),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_73),
.B1(n_78),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_8),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_96),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_96),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_9),
.A2(n_73),
.B1(n_78),
.B2(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_151),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_151),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_151),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_12),
.A2(n_38),
.B1(n_73),
.B2(n_78),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_103)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_30),
.B(n_32),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_105),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_104),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_54),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_25),
.A2(n_40),
.B(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_26),
.Y(n_142)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_27),
.A2(n_35),
.B(n_149),
.C(n_197),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_27),
.B(n_44),
.Y(n_231)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_30),
.A2(n_45),
.A3(n_47),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_31),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_32),
.A2(n_40),
.B1(n_65),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_32),
.A2(n_36),
.B(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_32),
.A2(n_40),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_32),
.B(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_32),
.A2(n_40),
.B1(n_201),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_32),
.A2(n_40),
.B1(n_221),
.B2(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_33),
.B(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_40),
.A2(n_66),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_42)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_43),
.A2(n_49),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_43),
.A2(n_49),
.B1(n_179),
.B2(n_234),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_46),
.B(n_72),
.Y(n_155)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_47),
.A2(n_74),
.B1(n_148),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_50),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_49),
.B(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_49),
.B(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_49),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_69),
.B1(n_81),
.B2(n_82),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_64),
.B1(n_82),
.B2(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_59),
.A2(n_118),
.B1(n_121),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_59),
.A2(n_61),
.B1(n_191),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_59),
.A2(n_89),
.B(n_193),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_60),
.A2(n_90),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_60),
.A2(n_63),
.B(n_120),
.Y(n_228)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_76),
.B(n_79),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_95),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_70),
.A2(n_128),
.B1(n_130),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_71),
.A2(n_75),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_73),
.B(n_149),
.CON(n_148),
.SN(n_148)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_75),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.C(n_98),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_85),
.B(n_91),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

OAI21x1_ASAP7_75t_SL g175 ( 
.A1(n_86),
.A2(n_121),
.B(n_157),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_101),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_111),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_109),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_111),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.C(n_126),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_112),
.A2(n_113),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_121),
.B(n_149),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_122),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_275),
.B(n_280),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_182),
.B(n_260),
.C(n_274),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_167),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_135),
.B(n_167),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_152),
.B2(n_166),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_138),
.B(n_139),
.C(n_166),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_153),
.B(n_159),
.C(n_163),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_156),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_168),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_177),
.B(n_247),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_259),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_254),
.B(n_258),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_242),
.B(n_253),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_224),
.B(n_241),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_213),
.B(n_223),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_202),
.B(n_212),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_194),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_207),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_222),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_232),
.B1(n_239),
.B2(n_240),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_251),
.C(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_262),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_268),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);


endmodule