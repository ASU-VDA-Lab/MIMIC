module real_jpeg_19465_n_11 (n_5, n_4, n_8, n_0, n_251, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_251;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_2),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_6),
.B1(n_16),
.B2(n_23),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_5),
.B1(n_16),
.B2(n_46),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_4),
.B1(n_16),
.B2(n_40),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_2),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_6),
.B1(n_23),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_4),
.B1(n_25),
.B2(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_1),
.A2(n_5),
.B1(n_25),
.B2(n_46),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_10),
.B1(n_17),
.B2(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_2),
.A2(n_20),
.B(n_33),
.C(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_7),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_9),
.B1(n_40),
.B2(n_47),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_10),
.B1(n_33),
.B2(n_40),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_4),
.A2(n_33),
.B(n_47),
.C(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_9),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_5),
.B(n_81),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_10),
.B1(n_33),
.B2(n_46),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_9),
.B(n_10),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_7),
.B1(n_23),
.B2(n_38),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_10),
.B1(n_23),
.B2(n_33),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_10),
.B(n_94),
.Y(n_93)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.C(n_139),
.Y(n_138)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_10),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_10),
.B(n_39),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_58),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_56),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_18),
.B1(n_26),
.B2(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_51),
.C(n_52),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_28),
.A2(n_29),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_42),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_30),
.A2(n_70),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_72),
.B(n_90),
.C(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_30),
.A2(n_70),
.B1(n_190),
.B2(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_30),
.A2(n_70),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_30),
.A2(n_191),
.B(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_30),
.A2(n_70),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_30),
.A2(n_70),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_33),
.B(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_33),
.B(n_84),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_33),
.A2(n_38),
.B(n_40),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_34),
.A2(n_42),
.B1(n_220),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_34),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_42),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_42),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_45),
.A2(n_48),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OA22x2_ASAP7_75t_SL g206 ( 
.A1(n_45),
.A2(n_48),
.B1(n_50),
.B2(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_46),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_51),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_243),
.B(n_249),
.Y(n_58)
);

OAI321xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_215),
.A3(n_235),
.B1(n_241),
.B2(n_242),
.C(n_251),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_200),
.B(n_214),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_182),
.B(n_199),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_109),
.B(n_164),
.C(n_181),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_98),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_64),
.B(n_98),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_87),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_66),
.B(n_78),
.C(n_87),
.Y(n_165)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI211xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_70),
.B(n_71),
.C(n_76),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_75),
.B1(n_79),
.B2(n_86),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_68),
.A2(n_75),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_75),
.B1(n_116),
.B2(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_95),
.C(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_68),
.A2(n_75),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_147),
.C(n_153),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_68),
.A2(n_75),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_68),
.B(n_79),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_171),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_70),
.B(n_73),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_70),
.B(n_220),
.C(n_222),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_70),
.B(n_229),
.C(n_234),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_71),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_75),
.B(n_141),
.C(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_72),
.A2(n_73),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_72),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_72),
.B(n_206),
.Y(n_207)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_95),
.C(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_74),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_97),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_88),
.A2(n_89),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_88),
.A2(n_89),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_105),
.B1(n_119),
.B2(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_95),
.A2(n_105),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_95),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g154 ( 
.A(n_95),
.B(n_138),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_106),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_100),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_102),
.B1(n_137),
.B2(n_141),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_163),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_156),
.B(n_162),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_143),
.B(n_155),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_134),
.B(n_142),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_123),
.B(n_133),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_118),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_180),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_177),
.C(n_180),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_174),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_179),
.B(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_187),
.B(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_201),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.CI(n_197),
.CON(n_185),
.SN(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_196),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_212),
.B2(n_213),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_209),
.C(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_217),
.B1(n_224),
.B2(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_212),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_227),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_227),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.C(n_225),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_226),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);


endmodule