module fake_jpeg_32100_n_385 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_385);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_385;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_11),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_9),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_40),
.B1(n_41),
.B2(n_17),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_63),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_62),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_72),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_16),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_41),
.B1(n_35),
.B2(n_17),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_40),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_34),
.B1(n_22),
.B2(n_38),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_82),
.A2(n_88),
.B1(n_96),
.B2(n_108),
.Y(n_145)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_89),
.A2(n_66),
.B1(n_54),
.B2(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_90),
.B(n_100),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_93),
.B(n_99),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_45),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_18),
.C(n_30),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_28),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_18),
.B1(n_30),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_112),
.B1(n_121),
.B2(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_43),
.B1(n_18),
.B2(n_27),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_111),
.B1(n_54),
.B2(n_57),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_43),
.B1(n_61),
.B2(n_67),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_47),
.A2(n_56),
.B1(n_43),
.B2(n_66),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_2),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_125),
.A2(n_130),
.B1(n_132),
.B2(n_143),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_51),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_133),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_106),
.B1(n_99),
.B2(n_121),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_69),
.B1(n_65),
.B2(n_68),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_135),
.B(n_136),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx2_ASAP7_75t_SL g137 ( 
.A(n_87),
.Y(n_137)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_62),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_59),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_144),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_77),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_27),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

BUFx2_ASAP7_75t_SL g149 ( 
.A(n_86),
.Y(n_149)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_150),
.A2(n_117),
.B1(n_20),
.B2(n_103),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_100),
.B(n_35),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_158),
.Y(n_186)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_53),
.B1(n_73),
.B2(n_70),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_81),
.A2(n_78),
.B1(n_28),
.B2(n_19),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_161),
.Y(n_182)
);

NOR4xp25_ASAP7_75t_SL g157 ( 
.A(n_89),
.B(n_11),
.C(n_9),
.D(n_8),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_83),
.A3(n_118),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_20),
.B(n_28),
.C(n_3),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_1),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g162 ( 
.A(n_92),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_20),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_92),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_20),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_20),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_116),
.B1(n_102),
.B2(n_95),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_196),
.B1(n_128),
.B2(n_139),
.Y(n_209)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_95),
.B1(n_116),
.B2(n_102),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_198),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_97),
.B1(n_118),
.B2(n_107),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_179),
.A2(n_131),
.B1(n_4),
.B2(n_7),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_103),
.B1(n_105),
.B2(n_92),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_94),
.C(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_117),
.C(n_114),
.Y(n_189)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_134),
.B1(n_147),
.B2(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_98),
.B1(n_97),
.B2(n_7),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_126),
.B(n_2),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_160),
.B(n_164),
.C(n_4),
.D(n_7),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_98),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_2),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_151),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_165),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_152),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_215),
.B1(n_184),
.B2(n_198),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_175),
.B(n_142),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_210),
.B(n_229),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_144),
.B(n_126),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_220),
.B(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_138),
.B(n_144),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_221),
.B(n_231),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_132),
.B1(n_140),
.B2(n_135),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_236),
.B1(n_196),
.B2(n_169),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_158),
.B(n_136),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_187),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_147),
.B1(n_131),
.B2(n_127),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_159),
.B(n_134),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_159),
.B(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_175),
.B(n_159),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_176),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_4),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_200),
.Y(n_252)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_173),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_174),
.C(n_181),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_249),
.C(n_251),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_174),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_261),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_257),
.B1(n_264),
.B2(n_232),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_206),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_169),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_211),
.B1(n_207),
.B2(n_234),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_169),
.Y(n_251)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_182),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_217),
.A2(n_190),
.B1(n_192),
.B2(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_172),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_217),
.A2(n_184),
.B1(n_188),
.B2(n_178),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_182),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_172),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_220),
.A2(n_189),
.B(n_178),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_243),
.B(n_241),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_271),
.B(n_283),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_278),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_275),
.B1(n_281),
.B2(n_286),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_210),
.Y(n_274)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_209),
.B1(n_218),
.B2(n_211),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_197),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_270),
.B1(n_263),
.B2(n_255),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_215),
.B1(n_231),
.B2(n_178),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_282),
.B(n_295),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_221),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_221),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_289),
.C(n_248),
.Y(n_296)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_230),
.B1(n_216),
.B2(n_222),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_244),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_219),
.Y(n_288)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_226),
.B1(n_228),
.B2(n_223),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_237),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_241),
.A2(n_250),
.B(n_243),
.C(n_249),
.D(n_269),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_297),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_270),
.B(n_259),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_176),
.B(n_173),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_288),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_277),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_302),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_310),
.B1(n_312),
.B2(n_314),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_173),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_279),
.A2(n_267),
.B1(n_246),
.B2(n_256),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_281),
.A2(n_236),
.B1(n_256),
.B2(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_258),
.B1(n_224),
.B2(n_227),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_258),
.B1(n_224),
.B2(n_235),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_271),
.C(n_292),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_318),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_280),
.C(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_324),
.C(n_326),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_292),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_280),
.C(n_276),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_276),
.C(n_283),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_309),
.A2(n_295),
.B(n_291),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_331),
.B(n_312),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_294),
.C(n_284),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_330),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_278),
.B1(n_252),
.B2(n_201),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_333),
.B1(n_316),
.B2(n_308),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_342),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_304),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_338),
.Y(n_358)
);

AOI31xp67_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_302),
.A3(n_316),
.B(n_304),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_323),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_310),
.B(n_314),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_340),
.A2(n_325),
.B(n_332),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_313),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_311),
.B(n_183),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_339),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_355),
.B(n_343),
.Y(n_361)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_320),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_353),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_330),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_324),
.C(n_325),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_353),
.C(n_352),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_321),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_356),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_331),
.C(n_323),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_347),
.Y(n_369)
);

OA21x2_ASAP7_75t_SL g359 ( 
.A1(n_344),
.A2(n_348),
.B(n_342),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_329),
.Y(n_360)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_360),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_183),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_343),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_369),
.C(n_240),
.Y(n_373)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_364),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_358),
.A2(n_347),
.B1(n_341),
.B2(n_346),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_366),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_366),
.A2(n_354),
.B(n_351),
.Y(n_372)
);

AOI322xp5_ASAP7_75t_L g377 ( 
.A1(n_372),
.A2(n_364),
.A3(n_367),
.B1(n_363),
.B2(n_368),
.C1(n_362),
.C2(n_365),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_374),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_201),
.C(n_183),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_R g380 ( 
.A(n_375),
.B(n_168),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_380),
.B(n_379),
.Y(n_382)
);

AOI322xp5_ASAP7_75t_L g378 ( 
.A1(n_370),
.A2(n_4),
.A3(n_168),
.B1(n_361),
.B2(n_371),
.C1(n_376),
.C2(n_374),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_378),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_168),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_383),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_381),
.Y(n_385)
);


endmodule