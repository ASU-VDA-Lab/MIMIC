module real_aes_7698_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g540 ( .A1(n_0), .A2(n_187), .B(n_541), .C(n_544), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_1), .B(n_529), .Y(n_545) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_91), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g432 ( .A(n_2), .Y(n_432) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_3), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_3), .Y(n_755) );
INVx1_ASAP7_75t_L g205 ( .A(n_4), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_5), .B(n_176), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_6), .A2(n_444), .B(n_523), .Y(n_522) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_7), .A2(n_152), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_8), .A2(n_37), .B1(n_132), .B2(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_9), .B(n_152), .Y(n_216) );
AND2x6_ASAP7_75t_L g150 ( .A(n_10), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_11), .A2(n_150), .B(n_447), .C(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_12), .B(n_38), .Y(n_433) );
INVx1_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_14), .B(n_139), .Y(n_159) );
INVx1_ASAP7_75t_L g197 ( .A(n_15), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_16), .B(n_176), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_17), .B(n_153), .Y(n_221) );
AO32x2_ASAP7_75t_L g184 ( .A1(n_18), .A2(n_149), .A3(n_152), .B1(n_185), .B2(n_189), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_19), .B(n_141), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_20), .B(n_153), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_21), .A2(n_53), .B1(n_132), .B2(n_141), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g138 ( .A1(n_22), .A2(n_82), .B1(n_139), .B2(n_141), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_23), .B(n_141), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_24), .A2(n_149), .B(n_447), .C(n_449), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_25), .A2(n_149), .B(n_447), .C(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_27), .B(n_144), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_28), .A2(n_444), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_29), .A2(n_103), .B1(n_114), .B2(n_762), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_30), .B(n_144), .Y(n_182) );
INVx2_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_32), .A2(n_468), .B(n_477), .C(n_479), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_33), .B(n_141), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_34), .B(n_144), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_35), .A2(n_74), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_35), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_36), .B(n_161), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_38), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_39), .B(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_40), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_41), .B(n_176), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_42), .B(n_444), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_43), .A2(n_468), .B(n_477), .C(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_44), .A2(n_122), .B1(n_426), .B2(n_427), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_44), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_44), .A2(n_80), .B1(n_426), .B2(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_45), .B(n_141), .Y(n_211) );
INVx1_ASAP7_75t_L g542 ( .A(n_46), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_47), .A2(n_90), .B1(n_132), .B2(n_135), .Y(n_131) );
INVx1_ASAP7_75t_L g515 ( .A(n_48), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_49), .B(n_141), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_141), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_51), .B(n_444), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_203), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_54), .A2(n_59), .B1(n_139), .B2(n_141), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_55), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_56), .B(n_141), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_57), .B(n_141), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_58), .Y(n_759) );
INVx1_ASAP7_75t_L g151 ( .A(n_60), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_61), .B(n_444), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_62), .B(n_529), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_63), .A2(n_200), .B(n_203), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_64), .B(n_141), .Y(n_206) );
INVx1_ASAP7_75t_L g147 ( .A(n_65), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_66), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_67), .B(n_176), .Y(n_481) );
AO32x2_ASAP7_75t_L g129 ( .A1(n_68), .A2(n_130), .A3(n_143), .B1(n_149), .B2(n_152), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_69), .B(n_142), .Y(n_505) );
INVx1_ASAP7_75t_L g239 ( .A(n_70), .Y(n_239) );
INVx1_ASAP7_75t_L g174 ( .A(n_71), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_72), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_73), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_75), .A2(n_447), .B(n_464), .C(n_468), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_76), .B(n_139), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_77), .Y(n_524) );
INVx1_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_79), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_80), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_81), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_83), .B(n_132), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_84), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_85), .B(n_139), .Y(n_179) );
INVx2_ASAP7_75t_L g145 ( .A(n_86), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_87), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_88), .B(n_136), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_89), .B(n_139), .Y(n_212) );
OR2x2_ASAP7_75t_L g430 ( .A(n_91), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g730 ( .A(n_91), .Y(n_730) );
OR2x2_ASAP7_75t_L g749 ( .A(n_91), .B(n_743), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_92), .A2(n_101), .B1(n_139), .B2(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_93), .B(n_444), .Y(n_475) );
INVx1_ASAP7_75t_L g480 ( .A(n_94), .Y(n_480) );
INVxp67_ASAP7_75t_L g527 ( .A(n_95), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_96), .B(n_139), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_97), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g465 ( .A(n_98), .Y(n_465) );
INVx1_ASAP7_75t_L g501 ( .A(n_99), .Y(n_501) );
AND2x2_ASAP7_75t_L g517 ( .A(n_100), .B(n_144), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_106), .Y(n_763) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO221x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_744), .B1(n_747), .B2(n_756), .C(n_758), .Y(n_114) );
OAI222xp33_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_119), .B1(n_731), .B2(n_732), .C1(n_738), .C2(n_739), .Y(n_115) );
INVx1_ASAP7_75t_L g731 ( .A(n_116), .Y(n_731) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_428), .B1(n_434), .B2(n_727), .Y(n_120) );
INVx1_ASAP7_75t_L g734 ( .A(n_121), .Y(n_734) );
INVx2_ASAP7_75t_L g427 ( .A(n_122), .Y(n_427) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_123), .B(n_752), .Y(n_751) );
AND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_346), .C(n_394), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_274), .C(n_319), .D(n_333), .Y(n_124) );
OAI311xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_190), .A3(n_217), .B1(n_227), .C1(n_242), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_154), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g227 ( .A1(n_127), .A2(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g335 ( .A(n_127), .B(n_262), .Y(n_335) );
AND2x2_ASAP7_75t_L g392 ( .A(n_127), .B(n_278), .Y(n_392) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g285 ( .A(n_128), .B(n_183), .Y(n_285) );
AND2x2_ASAP7_75t_L g342 ( .A(n_128), .B(n_290), .Y(n_342) );
INVx1_ASAP7_75t_L g383 ( .A(n_128), .Y(n_383) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_129), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_129), .B(n_183), .Y(n_292) );
AND2x2_ASAP7_75t_L g296 ( .A(n_129), .B(n_184), .Y(n_296) );
INVx1_ASAP7_75t_L g308 ( .A(n_129), .Y(n_308) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_136), .B1(n_138), .B2(n_142), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g135 ( .A(n_133), .Y(n_135) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
AND2x6_ASAP7_75t_L g447 ( .A(n_133), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_135), .Y(n_482) );
INVx2_ASAP7_75t_L g544 ( .A(n_135), .Y(n_544) );
INVx2_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_136), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_136), .A2(n_187), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g543 ( .A(n_136), .Y(n_543) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
INVx1_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
AND2x2_ASAP7_75t_L g445 ( .A(n_137), .B(n_204), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_137), .Y(n_448) );
INVx2_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_141), .Y(n_467) );
INVx5_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx1_ASAP7_75t_L g454 ( .A(n_143), .Y(n_454) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_144), .A2(n_156), .B(n_166), .Y(n_155) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_144), .A2(n_171), .B(n_182), .Y(n_170) );
INVx1_ASAP7_75t_L g457 ( .A(n_144), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_144), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_144), .A2(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_L g153 ( .A(n_145), .B(n_146), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_149), .B(n_223), .C(n_226), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_149), .A2(n_235), .B(n_238), .Y(n_234) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_150), .A2(n_157), .B(n_162), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_150), .A2(n_172), .B(n_177), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_150), .A2(n_196), .B(n_201), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_150), .A2(n_210), .B(n_213), .Y(n_209) );
AND2x4_ASAP7_75t_L g444 ( .A(n_150), .B(n_445), .Y(n_444) );
INVx4_ASAP7_75t_SL g469 ( .A(n_150), .Y(n_469) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_150), .B(n_445), .Y(n_502) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_152), .A2(n_209), .B(n_216), .Y(n_208) );
INVx4_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_152), .A2(n_492), .B(n_493), .Y(n_491) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_152), .Y(n_521) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_167), .Y(n_154) );
AND2x2_ASAP7_75t_L g229 ( .A(n_155), .B(n_183), .Y(n_229) );
INVx2_ASAP7_75t_L g263 ( .A(n_155), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_155), .B(n_184), .Y(n_278) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_155), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_155), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g298 ( .A(n_155), .B(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g310 ( .A(n_155), .Y(n_310) );
INVx1_ASAP7_75t_L g351 ( .A(n_155), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_155), .B(n_251), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_L g238 ( .A1(n_165), .A2(n_202), .B(n_239), .C(n_240), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g228 ( .A(n_169), .B(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_169), .Y(n_256) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_169), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g313 ( .A(n_169), .B(n_183), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_169), .B(n_308), .Y(n_371) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g261 ( .A(n_170), .Y(n_261) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_170), .Y(n_277) );
OR2x2_ASAP7_75t_L g350 ( .A(n_170), .B(n_351), .Y(n_350) );
O2A1O1Ixp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
INVx2_ASAP7_75t_L g187 ( .A(n_176), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_176), .A2(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_176), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g200 ( .A(n_180), .Y(n_200) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g451 ( .A(n_181), .Y(n_451) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx2_ASAP7_75t_L g257 ( .A(n_184), .Y(n_257) );
AND2x2_ASAP7_75t_L g262 ( .A(n_184), .B(n_263), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_187), .A2(n_202), .B(n_205), .C(n_206), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_187), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g194 ( .A(n_189), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_189), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_190), .B(n_245), .Y(n_408) );
INVx1_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g378 ( .A(n_191), .B(n_219), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_208), .Y(n_191) );
AND2x2_ASAP7_75t_L g254 ( .A(n_192), .B(n_245), .Y(n_254) );
INVx2_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
AND2x2_ASAP7_75t_L g300 ( .A(n_192), .B(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g367 ( .A(n_192), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_193), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g247 ( .A(n_193), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g287 ( .A(n_193), .B(n_208), .Y(n_287) );
AND2x2_ASAP7_75t_L g304 ( .A(n_193), .B(n_305), .Y(n_304) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_207), .Y(n_193) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_234), .B(n_241), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .C(n_200), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_198), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_198), .A2(n_505), .B(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_200), .A2(n_465), .B(n_466), .C(n_467), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_202), .A2(n_450), .B(n_452), .Y(n_449) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g230 ( .A(n_208), .B(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
AND2x2_ASAP7_75t_L g253 ( .A(n_208), .B(n_233), .Y(n_253) );
AND2x2_ASAP7_75t_L g326 ( .A(n_208), .B(n_305), .Y(n_326) );
AND2x2_ASAP7_75t_L g391 ( .A(n_208), .B(n_381), .Y(n_391) );
OAI311xp33_ASAP7_75t_L g274 ( .A1(n_217), .A2(n_275), .A3(n_279), .B1(n_281), .C1(n_301), .Y(n_274) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g286 ( .A(n_218), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g345 ( .A(n_218), .B(n_253), .Y(n_345) );
AND2x2_ASAP7_75t_L g419 ( .A(n_218), .B(n_300), .Y(n_419) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_219), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g354 ( .A(n_219), .Y(n_354) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g245 ( .A(n_220), .Y(n_245) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_220), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g374 ( .A(n_220), .B(n_248), .Y(n_374) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
AO21x1_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_226), .B(n_271), .Y(n_270) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_226), .A2(n_462), .B(n_471), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_226), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_226), .B(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_226), .A2(n_500), .B(n_507), .Y(n_499) );
INVx3_ASAP7_75t_L g529 ( .A(n_226), .Y(n_529) );
AND2x2_ASAP7_75t_L g249 ( .A(n_229), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g302 ( .A(n_229), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g382 ( .A(n_229), .B(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_230), .A2(n_262), .B1(n_282), .B2(n_286), .C(n_288), .Y(n_281) );
INVx1_ASAP7_75t_L g406 ( .A(n_231), .Y(n_406) );
OR2x2_ASAP7_75t_L g372 ( .A(n_232), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g267 ( .A(n_233), .B(n_248), .Y(n_267) );
OR2x2_ASAP7_75t_L g269 ( .A(n_233), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g294 ( .A(n_233), .Y(n_294) );
INVx2_ASAP7_75t_L g305 ( .A(n_233), .Y(n_305) );
AND2x2_ASAP7_75t_L g332 ( .A(n_233), .B(n_270), .Y(n_332) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_233), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B1(n_252), .B2(n_255), .C(n_258), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g343 ( .A(n_245), .B(n_253), .Y(n_343) );
AND2x2_ASAP7_75t_L g393 ( .A(n_245), .B(n_247), .Y(n_393) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g280 ( .A(n_247), .B(n_251), .Y(n_280) );
AND2x2_ASAP7_75t_L g359 ( .A(n_247), .B(n_332), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_248), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g318 ( .A(n_248), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_249), .A2(n_329), .B(n_331), .Y(n_328) );
OR2x2_ASAP7_75t_L g272 ( .A(n_250), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_298), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_250), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g315 ( .A(n_251), .B(n_284), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_251), .B(n_398), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_252), .B(n_278), .Y(n_388) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g311 ( .A(n_253), .B(n_266), .Y(n_311) );
INVx1_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B1(n_268), .B2(n_272), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g290 ( .A(n_261), .Y(n_290) );
INVx1_ASAP7_75t_L g303 ( .A(n_261), .Y(n_303) );
INVx1_ASAP7_75t_L g273 ( .A(n_262), .Y(n_273) );
AND2x2_ASAP7_75t_L g344 ( .A(n_262), .B(n_290), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_262), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
OR2x2_ASAP7_75t_L g268 ( .A(n_265), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_265), .B(n_381), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_265), .B(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g415 ( .A(n_267), .B(n_367), .Y(n_415) );
INVx1_ASAP7_75t_SL g381 ( .A(n_269), .Y(n_381) );
AND2x2_ASAP7_75t_L g321 ( .A(n_270), .B(n_305), .Y(n_321) );
INVx1_ASAP7_75t_L g368 ( .A(n_270), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_275), .A2(n_365), .B1(n_410), .B2(n_411), .C1(n_414), .C2(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
AND2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_278), .B(n_383), .Y(n_410) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_280), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g385 ( .A(n_282), .Y(n_385) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g323 ( .A(n_285), .Y(n_323) );
AND2x2_ASAP7_75t_L g402 ( .A(n_285), .B(n_363), .Y(n_402) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_309), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_287), .B(n_321), .Y(n_320) );
OAI32xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .A3(n_293), .B1(n_295), .B2(n_299), .Y(n_288) );
BUFx2_ASAP7_75t_L g363 ( .A(n_290), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_291), .B(n_309), .Y(n_390) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_292), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g397 ( .A(n_292), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g386 ( .A(n_293), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g357 ( .A(n_296), .B(n_330), .Y(n_357) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OAI221xp5_ASAP7_75t_SL g319 ( .A1(n_298), .A2(n_320), .B1(n_322), .B2(n_324), .C(n_328), .Y(n_319) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g337 ( .A(n_300), .B(n_321), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B1(n_306), .B2(n_311), .C(n_312), .Y(n_301) );
INVx1_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_303), .B(n_397), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_304), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_309), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
BUFx3_ASAP7_75t_L g398 ( .A(n_310), .Y(n_398) );
INVx1_ASAP7_75t_SL g339 ( .A(n_311), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_311), .B(n_353), .Y(n_352) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_313), .A2(n_414), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_321), .Y(n_360) );
INVx1_ASAP7_75t_L g424 ( .A(n_318), .Y(n_424) );
INVx2_ASAP7_75t_L g413 ( .A(n_321), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_321), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B1(n_338), .B2(n_339), .C(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_342), .A2(n_404), .B1(n_405), .B2(n_407), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_345), .A2(n_422), .B(n_425), .Y(n_421) );
NOR4xp25_ASAP7_75t_SL g346 ( .A(n_347), .B(n_355), .C(n_364), .D(n_384), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B1(n_361), .B2(n_362), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B1(n_372), .B2(n_375), .C(n_376), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_379), .B(n_382), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .C(n_389), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_389) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_393), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_409), .C(n_417), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_395) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g735 ( .A(n_429), .Y(n_735) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g729 ( .A(n_431), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g743 ( .A(n_431), .Y(n_743) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g736 ( .A(n_435), .Y(n_736) );
AND3x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_631), .C(n_688), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_576), .C(n_612), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_485), .B(n_531), .C(n_563), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_458), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g534 ( .A(n_440), .B(n_535), .Y(n_534) );
INVx5_ASAP7_75t_L g562 ( .A(n_440), .Y(n_562) );
AND2x2_ASAP7_75t_L g635 ( .A(n_440), .B(n_551), .Y(n_635) );
AND2x2_ASAP7_75t_L g673 ( .A(n_440), .B(n_579), .Y(n_673) );
AND2x2_ASAP7_75t_L g693 ( .A(n_440), .B(n_536), .Y(n_693) );
OR2x6_ASAP7_75t_L g440 ( .A(n_441), .B(n_455), .Y(n_440) );
AOI21xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_446), .B(n_454), .Y(n_441) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
INVx2_ASAP7_75t_L g453 ( .A(n_451), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_453), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_453), .A2(n_482), .B(n_515), .C(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_458), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_473), .Y(n_458) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_459), .Y(n_574) );
AND2x2_ASAP7_75t_L g588 ( .A(n_459), .B(n_535), .Y(n_588) );
INVx1_ASAP7_75t_L g611 ( .A(n_459), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_459), .B(n_562), .Y(n_650) );
OR2x2_ASAP7_75t_L g687 ( .A(n_459), .B(n_533), .Y(n_687) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_460), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_460), .B(n_536), .Y(n_630) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_536), .Y(n_551) );
BUFx2_ASAP7_75t_L g579 ( .A(n_461), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_469), .A2(n_478), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g538 ( .A1(n_469), .A2(n_478), .B(n_539), .C(n_540), .Y(n_538) );
INVx5_ASAP7_75t_L g533 ( .A(n_473), .Y(n_533) );
BUFx2_ASAP7_75t_L g555 ( .A(n_473), .Y(n_555) );
AND2x2_ASAP7_75t_L g712 ( .A(n_473), .B(n_566), .Y(n_712) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_518), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_487), .A2(n_613), .B1(n_620), .B2(n_621), .C(n_624), .Y(n_612) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
AND2x2_ASAP7_75t_L g519 ( .A(n_488), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_488), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g547 ( .A(n_489), .B(n_498), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_489), .B(n_499), .Y(n_557) );
OR2x2_ASAP7_75t_L g568 ( .A(n_489), .B(n_520), .Y(n_568) );
AND2x2_ASAP7_75t_L g571 ( .A(n_489), .B(n_559), .Y(n_571) );
AND2x2_ASAP7_75t_L g587 ( .A(n_489), .B(n_509), .Y(n_587) );
OR2x2_ASAP7_75t_L g603 ( .A(n_489), .B(n_499), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_489), .B(n_520), .Y(n_665) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_490), .B(n_509), .Y(n_657) );
AND2x2_ASAP7_75t_L g660 ( .A(n_490), .B(n_499), .Y(n_660) );
OR2x2_ASAP7_75t_L g581 ( .A(n_497), .B(n_568), .Y(n_581) );
INVx2_ASAP7_75t_L g607 ( .A(n_497), .Y(n_607) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_509), .Y(n_497) );
AND2x2_ASAP7_75t_L g530 ( .A(n_498), .B(n_510), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_498), .B(n_520), .Y(n_586) );
OR2x2_ASAP7_75t_L g597 ( .A(n_498), .B(n_510), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_498), .B(n_559), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g689 ( .A1(n_498), .A2(n_690), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_689) );
INVx5_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_499), .B(n_520), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_503), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_509), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_509), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g575 ( .A(n_509), .B(n_547), .Y(n_575) );
OR2x2_ASAP7_75t_L g619 ( .A(n_509), .B(n_520), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_509), .B(n_571), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_509), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g684 ( .A(n_509), .B(n_685), .Y(n_684) );
INVx5_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_SL g548 ( .A(n_510), .B(n_519), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_510), .A2(n_553), .B(n_556), .C(n_560), .Y(n_552) );
OR2x2_ASAP7_75t_L g590 ( .A(n_510), .B(n_586), .Y(n_590) );
OR2x2_ASAP7_75t_L g626 ( .A(n_510), .B(n_568), .Y(n_626) );
OAI311xp33_ASAP7_75t_L g632 ( .A1(n_510), .A2(n_571), .A3(n_633), .B1(n_636), .C1(n_643), .Y(n_632) );
AND2x2_ASAP7_75t_L g683 ( .A(n_510), .B(n_520), .Y(n_683) );
AND2x2_ASAP7_75t_L g691 ( .A(n_510), .B(n_546), .Y(n_691) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_510), .Y(n_709) );
AND2x2_ASAP7_75t_L g726 ( .A(n_510), .B(n_547), .Y(n_726) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
AND2x2_ASAP7_75t_L g554 ( .A(n_519), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g710 ( .A(n_519), .Y(n_710) );
AND2x2_ASAP7_75t_L g546 ( .A(n_520), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_520), .Y(n_602) );
INVxp67_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_528), .Y(n_520) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_529), .A2(n_537), .B(n_545), .Y(n_536) );
AND2x2_ASAP7_75t_L g719 ( .A(n_530), .B(n_567), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_546), .B1(n_548), .B2(n_549), .C(n_552), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_533), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g572 ( .A(n_533), .B(n_562), .Y(n_572) );
AND2x2_ASAP7_75t_L g580 ( .A(n_533), .B(n_535), .Y(n_580) );
OR2x2_ASAP7_75t_L g592 ( .A(n_533), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g610 ( .A(n_533), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g634 ( .A(n_533), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_533), .Y(n_654) );
AND2x2_ASAP7_75t_L g706 ( .A(n_533), .B(n_630), .Y(n_706) );
OAI31xp33_ASAP7_75t_L g714 ( .A1(n_533), .A2(n_583), .A3(n_682), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_534), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g678 ( .A(n_534), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_534), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_L g566 ( .A(n_535), .B(n_562), .Y(n_566) );
INVx1_ASAP7_75t_L g653 ( .A(n_535), .Y(n_653) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g703 ( .A(n_536), .B(n_562), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_SL g713 ( .A(n_546), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_547), .B(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_548), .A2(n_660), .B1(n_698), .B2(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g561 ( .A(n_551), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g620 ( .A(n_551), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_551), .B(n_572), .Y(n_725) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g695 ( .A(n_554), .B(n_696), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_555), .A2(n_614), .B(n_616), .Y(n_613) );
OR2x2_ASAP7_75t_L g621 ( .A(n_555), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g642 ( .A(n_555), .B(n_630), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_555), .B(n_653), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_555), .B(n_693), .Y(n_692) );
OAI221xp5_ASAP7_75t_SL g669 ( .A1(n_556), .A2(n_670), .B1(n_675), .B2(n_678), .C(n_679), .Y(n_669) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OR2x2_ASAP7_75t_L g646 ( .A(n_557), .B(n_619), .Y(n_646) );
INVx1_ASAP7_75t_L g685 ( .A(n_557), .Y(n_685) );
INVx2_ASAP7_75t_L g661 ( .A(n_558), .Y(n_661) );
INVx1_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_562), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g629 ( .A(n_562), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g717 ( .A(n_562), .B(n_687), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_567), .B1(n_569), .B2(n_572), .C1(n_573), .C2(n_575), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_566), .A2(n_616), .B1(n_644), .B2(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_566), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI21xp33_ASAP7_75t_SL g604 ( .A1(n_575), .A2(n_605), .B(n_608), .Y(n_604) );
OAI211xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_581), .B(n_582), .C(n_604), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_580), .A2(n_583), .B1(n_588), .B2(n_589), .C(n_591), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_580), .B(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_L g674 ( .A(n_580), .Y(n_674) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g676 ( .A(n_585), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g593 ( .A(n_588), .Y(n_593) );
AND2x2_ASAP7_75t_L g599 ( .A(n_588), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B1(n_598), .B2(n_601), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_595), .B(n_607), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_596), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g696 ( .A(n_600), .Y(n_696) );
AND2x2_ASAP7_75t_L g715 ( .A(n_600), .B(n_630), .Y(n_715) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_607), .B(n_664), .Y(n_723) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_610), .B(n_678), .Y(n_721) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g644 ( .A(n_622), .Y(n_644) );
BUFx2_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_627), .B(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_647), .C(n_669), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_642), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_651), .B(n_655), .C(n_658), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_648), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp67_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_SL g677 ( .A(n_657), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_666), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
AND2x2_ASAP7_75t_L g682 ( .A(n_660), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B1(n_684), .B2(n_686), .Y(n_679) );
INVx2_ASAP7_75t_SL g700 ( .A(n_687), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_704), .C(n_716), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_700), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_711), .B2(n_713), .C(n_714), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_705), .A2(n_717), .B(n_718), .C(n_720), .Y(n_716) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_724), .B2(n_726), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g737 ( .A(n_728), .Y(n_737) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_730), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g757 ( .A(n_745), .Y(n_757) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g761 ( .A(n_749), .Y(n_761) );
INVx1_ASAP7_75t_L g754 ( .A(n_751), .Y(n_754) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
endmodule