module fake_aes_5703_n_33 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_13), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI211xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_14), .B(n_18), .C(n_16), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_22), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_17), .B1(n_15), .B2(n_13), .C(n_4), .Y(n_26) );
OAI22xp33_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_27) );
AOI211xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_2), .B(n_4), .C(n_5), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI22xp5_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OAI22xp5_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_30), .B1(n_8), .B2(n_7), .Y(n_32) );
AOI22xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_33) );
endmodule