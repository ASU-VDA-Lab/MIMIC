module fake_jpeg_12189_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2x1_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_32),
.B1(n_13),
.B2(n_14),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_24),
.B1(n_15),
.B2(n_17),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_19),
.B(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_11),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_36),
.C(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_65),
.C(n_38),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_47),
.C(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_13),
.C(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_47),
.B1(n_54),
.B2(n_64),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_37),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_55),
.C(n_61),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_80),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_62),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_44),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_65),
.C(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_55),
.B1(n_61),
.B2(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_93),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_13),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_66),
.C(n_13),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_72),
.A3(n_80),
.B1(n_68),
.B2(n_73),
.C1(n_67),
.C2(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_102),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_79),
.B(n_70),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_101),
.B(n_0),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_90),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_81),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_12),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_111),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_95),
.B(n_93),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_112),
.B(n_99),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_9),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_14),
.C(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_10),
.C(n_3),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_113),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_121),
.B(n_107),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_126),
.C(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_106),
.B(n_3),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_130),
.C(n_6),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_116),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_127),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_0),
.B(n_4),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B1(n_4),
.B2(n_6),
.Y(n_136)
);


endmodule