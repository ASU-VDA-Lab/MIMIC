module fake_jpeg_30790_n_106 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.C(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_20),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_30),
.B(n_36),
.C(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_11),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_42),
.Y(n_56)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_28),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_45),
.C(n_31),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_54),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_36),
.B1(n_27),
.B2(n_28),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_18),
.C(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_53),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_46),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_38),
.B1(n_37),
.B2(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_19),
.B(n_17),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_26),
.B(n_19),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_40),
.B(n_26),
.C(n_17),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_50),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_72),
.C(n_64),
.Y(n_77)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_52),
.C(n_27),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_75),
.B(n_66),
.C(n_26),
.D(n_3),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_65),
.B1(n_64),
.B2(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_62),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_1),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_67),
.B1(n_79),
.B2(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_67),
.B1(n_93),
.B2(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_87),
.B(n_76),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_97),
.B(n_6),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_2),
.C(n_5),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_99),
.A2(n_101),
.B(n_6),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_6),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_102),
.B(n_2),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_5),
.Y(n_106)
);


endmodule