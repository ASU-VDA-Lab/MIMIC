module fake_jpeg_10393_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_8),
.B(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_8),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_23),
.B1(n_19),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_52),
.B1(n_27),
.B2(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_63),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_17),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_41),
.B1(n_24),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_77),
.B1(n_83),
.B2(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_70),
.B(n_32),
.Y(n_122)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_79),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_17),
.B1(n_21),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_28),
.B1(n_68),
.B2(n_87),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_52),
.B1(n_47),
.B2(n_55),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_15),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_89),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_21),
.B1(n_29),
.B2(n_28),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_38),
.C(n_26),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_26),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_103),
.C(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_98),
.B(n_111),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_101),
.B1(n_80),
.B2(n_61),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_76),
.B(n_91),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_38),
.B(n_26),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_108),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_26),
.C(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_33),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_1),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_115),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_60),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_95),
.B1(n_92),
.B2(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_122),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_32),
.B(n_25),
.C(n_18),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_120),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_132),
.C(n_97),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_127),
.B(n_130),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_129),
.B1(n_149),
.B2(n_121),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_93),
.B1(n_83),
.B2(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_135),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_67),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_112),
.B1(n_124),
.B2(n_107),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_107),
.B1(n_115),
.B2(n_119),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_143),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_81),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_140),
.Y(n_165)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_146),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_147),
.Y(n_177)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_111),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_151),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_11),
.C(n_13),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_103),
.B(n_100),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_163),
.B(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_172),
.B1(n_184),
.B2(n_73),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_99),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_164),
.C(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_160),
.B(n_169),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_110),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_98),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_97),
.C(n_117),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_109),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_138),
.C(n_134),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_88),
.B(n_109),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_126),
.A2(n_75),
.B1(n_25),
.B2(n_18),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_183),
.B1(n_121),
.B2(n_139),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_126),
.A2(n_18),
.B1(n_78),
.B2(n_73),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_127),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_196),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_145),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_195),
.C(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_193),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_131),
.B1(n_151),
.B2(n_135),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_204),
.B1(n_210),
.B2(n_203),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_134),
.C(n_142),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_167),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_158),
.B1(n_172),
.B2(n_166),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_1),
.C(n_2),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.C(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_1),
.C(n_2),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_178),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_155),
.B(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_161),
.B1(n_181),
.B2(n_160),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_194),
.B1(n_201),
.B2(n_208),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_163),
.B(n_179),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_162),
.C(n_185),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_195),
.C(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_180),
.B(n_170),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_231),
.B1(n_207),
.B2(n_210),
.Y(n_241)
);

AO22x1_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_182),
.B1(n_167),
.B2(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_168),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_1),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_189),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_242),
.C(n_247),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_245),
.B1(n_231),
.B2(n_227),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_235),
.B(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_198),
.C(n_209),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_218),
.C(n_224),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_223),
.B1(n_228),
.B2(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_222),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_233),
.B(n_223),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_260),
.B(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.C(n_265),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_230),
.B(n_214),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_217),
.B1(n_214),
.B2(n_229),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_225),
.C(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_247),
.C(n_239),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_274),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_276),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_236),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_245),
.C(n_222),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_263),
.B(n_7),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_267),
.B(n_260),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_284),
.B(n_285),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_261),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_263),
.B1(n_265),
.B2(n_9),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.C(n_276),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_292),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_271),
.A3(n_268),
.B1(n_269),
.B2(n_6),
.C1(n_10),
.C2(n_12),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

AOI321xp33_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_6),
.A3(n_10),
.B1(n_12),
.B2(n_2),
.C(n_4),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_298),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_293),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_297),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_4),
.A3(n_5),
.B1(n_12),
.B2(n_293),
.C1(n_300),
.C2(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_5),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_5),
.Y(n_305)
);


endmodule