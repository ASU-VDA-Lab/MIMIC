module fake_jpeg_9238_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_0),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_34),
.B1(n_21),
.B2(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_41),
.B1(n_36),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_41),
.B1(n_36),
.B2(n_44),
.Y(n_80)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_44),
.B1(n_18),
.B2(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_80),
.B1(n_28),
.B2(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_90),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_24),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_24),
.B(n_43),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_68),
.B1(n_18),
.B2(n_44),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_40),
.C(n_43),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_39),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_97),
.Y(n_103)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_89),
.C(n_43),
.Y(n_132)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_31),
.B1(n_30),
.B2(n_17),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_65),
.B1(n_59),
.B2(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_114),
.B1(n_117),
.B2(n_77),
.Y(n_133)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_126),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_59),
.B1(n_44),
.B2(n_64),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_125),
.B1(n_22),
.B2(n_28),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_38),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_84),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_27),
.B(n_22),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_90),
.B(n_97),
.C(n_88),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_95),
.B1(n_30),
.B2(n_32),
.Y(n_147)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_101),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_145),
.C(n_149),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_135),
.B1(n_146),
.B2(n_107),
.Y(n_154)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_89),
.B1(n_77),
.B2(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_43),
.C(n_92),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_78),
.B1(n_86),
.B2(n_28),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_116),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_86),
.C(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_152),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_31),
.A3(n_30),
.B1(n_17),
.B2(n_20),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_153),
.B1(n_123),
.B2(n_31),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_171),
.B1(n_105),
.B2(n_141),
.Y(n_195)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_159),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_119),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_124),
.B1(n_114),
.B2(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_115),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_162),
.C(n_180),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_112),
.C(n_121),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_118),
.C(n_126),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_105),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_129),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_189),
.B(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_139),
.B1(n_152),
.B2(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_193),
.B1(n_158),
.B2(n_154),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_127),
.B1(n_138),
.B2(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_20),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_141),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_99),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_110),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_120),
.C(n_136),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_21),
.B(n_29),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_120),
.B(n_104),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_26),
.B(n_157),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_19),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_82),
.C(n_26),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_172),
.B1(n_167),
.B2(n_29),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_179),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_234),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_232),
.B1(n_233),
.B2(n_182),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_222),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_82),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_82),
.B1(n_20),
.B2(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_186),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_193),
.C(n_9),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_190),
.C(n_200),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_245),
.C(n_251),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_190),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_202),
.C(n_199),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_188),
.B1(n_197),
.B2(n_198),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_254),
.B1(n_224),
.B2(n_219),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_196),
.C(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_225),
.C(n_219),
.Y(n_265)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_7),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_256),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_262),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_230),
.B1(n_218),
.B2(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_239),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_268),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_270),
.B1(n_8),
.B2(n_14),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_226),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_235),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_217),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_217),
.B1(n_220),
.B2(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_241),
.B(n_220),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_8),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.C(n_242),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_0),
.C(n_1),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

FAx1_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_244),
.CI(n_249),
.CON(n_281),
.SN(n_281)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_287),
.Y(n_300)
);

NOR2x1_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_238),
.C(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_286),
.C(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_251),
.C(n_255),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_257),
.CI(n_240),
.CON(n_288),
.SN(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_265),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_10),
.B1(n_14),
.B2(n_4),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_259),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_293),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_297),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.C(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_258),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_275),
.C(n_2),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_8),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_1),
.C(n_2),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_6),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_11),
.B1(n_14),
.B2(n_5),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_283),
.C(n_288),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_281),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_300),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_287),
.C(n_12),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_15),
.C(n_1),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_15),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_298),
.B1(n_12),
.B2(n_6),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_300),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_10),
.B(n_13),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_313),
.B(n_15),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_306),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_326),
.B(n_320),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_316),
.B(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.C(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_324),
.B(n_3),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_3),
.B(n_308),
.Y(n_332)
);


endmodule