module fake_jpeg_6837_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_43),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_19),
.B1(n_23),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_31),
.B1(n_25),
.B2(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_22),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_33),
.B2(n_26),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_24),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_78),
.B(n_93),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_84),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_42),
.B(n_27),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_67),
.B1(n_48),
.B2(n_61),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_42),
.C(n_43),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_67),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_46),
.B1(n_49),
.B2(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_0),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_58),
.B1(n_66),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_102),
.B1(n_103),
.B2(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_107),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_66),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_114),
.C(n_76),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_46),
.B1(n_67),
.B2(n_54),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_67),
.B1(n_54),
.B2(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_45),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_53),
.B1(n_49),
.B2(n_61),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_94),
.B1(n_72),
.B2(n_79),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_86),
.B(n_68),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_124),
.B(n_138),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_69),
.C(n_76),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_130),
.C(n_131),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_68),
.B(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_133),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_76),
.C(n_93),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_51),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_84),
.B(n_87),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_140),
.B(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_139),
.B1(n_120),
.B2(n_96),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_85),
.B1(n_48),
.B2(n_57),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_87),
.B(n_34),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_11),
.C(n_16),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_149),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_32),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_79),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_117),
.B1(n_115),
.B2(n_113),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_166),
.B1(n_180),
.B2(n_126),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_106),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_173),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_167),
.B(n_2),
.Y(n_203)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_106),
.B(n_107),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_177),
.CI(n_136),
.CON(n_182),
.SN(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_108),
.B1(n_120),
.B2(n_96),
.Y(n_166)
);

NAND2x1_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_147),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_120),
.B1(n_119),
.B2(n_111),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_111),
.B1(n_90),
.B2(n_70),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_34),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_119),
.C(n_90),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_123),
.C(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_1),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_70),
.B1(n_91),
.B2(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_190),
.Y(n_215)
);

NOR4xp25_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_140),
.C(n_138),
.D(n_128),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_165),
.B(n_179),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_131),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_191),
.C(n_202),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_135),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_125),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_151),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_133),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_204),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_160),
.C(n_159),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_169),
.B(n_5),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_166),
.B1(n_177),
.B2(n_156),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_220),
.B(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_196),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_172),
.B1(n_175),
.B2(n_160),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_214),
.B1(n_187),
.B2(n_200),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_163),
.B1(n_157),
.B2(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_174),
.B(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_174),
.C(n_155),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_154),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_169),
.C(n_5),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_181),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_4),
.C(n_6),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_217),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_237),
.Y(n_253)
);

OAI321xp33_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_183),
.A3(n_192),
.B1(n_182),
.B2(n_194),
.C(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_182),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_236),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_185),
.B1(n_205),
.B2(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_186),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_243),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_192),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_199),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_215),
.B1(n_205),
.B2(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_209),
.B1(n_222),
.B2(n_211),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_260),
.B(n_261),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_226),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_209),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_245),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_225),
.C(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_216),
.C(n_184),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_236),
.B1(n_231),
.B2(n_243),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_268),
.B1(n_269),
.B2(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_274),
.C(n_253),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_239),
.B(n_235),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_239),
.B(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_188),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_230),
.B(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_219),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_249),
.B(n_256),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_276),
.B(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_228),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_260),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_283),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_216),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_251),
.B1(n_238),
.B2(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_275),
.A3(n_280),
.B1(n_259),
.B2(n_206),
.C1(n_229),
.C2(n_12),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_293),
.A3(n_294),
.B1(n_295),
.B2(n_286),
.C1(n_290),
.C2(n_289),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_287),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_12),
.A3(n_15),
.B1(n_9),
.B2(n_10),
.C1(n_16),
.C2(n_13),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_9),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_6),
.C2(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_14),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.Y(n_301)
);


endmodule