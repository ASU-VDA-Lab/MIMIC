module fake_ariane_1174_n_978 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_978);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_978;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_928;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_933;
wire n_774;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_931;
wire n_827;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_23),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_17),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_178),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_19),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_55),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_32),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_103),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_99),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_109),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_136),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_204),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_94),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_191),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_54),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_188),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_127),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_118),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_36),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_143),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_201),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_160),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_84),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_93),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_135),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_164),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_56),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_182),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_154),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_77),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_61),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_15),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_157),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_20),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_172),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_189),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_116),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_69),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_105),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_161),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_163),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_141),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_180),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_59),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_72),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_166),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_203),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_221),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_211),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_226),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_215),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_223),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_209),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_229),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_225),
.B(n_232),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_274),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_252),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_290),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_235),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_225),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_273),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_210),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_279),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_210),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_269),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_0),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_216),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_227),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_230),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_231),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_220),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_222),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_234),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_237),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_238),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_243),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_228),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_270),
.B(n_1),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_236),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_239),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_271),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_240),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

OR2x2_ASAP7_75t_SL g358 ( 
.A(n_305),
.B(n_246),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_293),
.B(n_284),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_217),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_344),
.B(n_249),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_344),
.B(n_246),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_247),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_265),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_259),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_319),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_265),
.B(n_260),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_299),
.B(n_242),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_213),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_213),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_350),
.B(n_241),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_352),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_R g412 ( 
.A(n_402),
.B(n_316),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_245),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_301),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_301),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_400),
.B(n_213),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_315),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_394),
.B1(n_381),
.B2(n_398),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_315),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_398),
.A2(n_296),
.B1(n_295),
.B2(n_292),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_374),
.B(n_248),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_251),
.B1(n_258),
.B2(n_276),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_400),
.B(n_251),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_250),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_373),
.B(n_253),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_256),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_251),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_251),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_289),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_393),
.B(n_258),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_397),
.B(n_257),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

BUFx6f_ASAP7_75t_SL g446 ( 
.A(n_370),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_361),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_370),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_368),
.B(n_261),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

AND2x2_ASAP7_75t_SL g455 ( 
.A(n_371),
.B(n_258),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_262),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_383),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_354),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_382),
.B(n_263),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_382),
.B(n_264),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_258),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_266),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_376),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_395),
.B(n_288),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_276),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_366),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_395),
.B(n_267),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_276),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_385),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_369),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_355),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_359),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_383),
.B(n_276),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_390),
.B(n_369),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_375),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_390),
.B(n_1),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_375),
.B(n_286),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_379),
.A2(n_247),
.B(n_268),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_390),
.B(n_2),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_372),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_457),
.B(n_402),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_416),
.A2(n_406),
.B1(n_404),
.B2(n_402),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_422),
.A2(n_473),
.B1(n_431),
.B2(n_413),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_436),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_486),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_404),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_433),
.B(n_385),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

AO22x2_ASAP7_75t_L g499 ( 
.A1(n_424),
.A2(n_406),
.B1(n_403),
.B2(n_407),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_403),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_465),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_404),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_410),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_458),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g509 ( 
.A1(n_424),
.A2(n_407),
.B1(n_408),
.B2(n_410),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_417),
.A2(n_408),
.B1(n_405),
.B2(n_367),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_454),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_385),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_417),
.A2(n_399),
.B1(n_365),
.B2(n_358),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_421),
.A2(n_358),
.B1(n_380),
.B2(n_387),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_480),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_421),
.A2(n_485),
.B1(n_479),
.B2(n_484),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_391),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_433),
.B(n_399),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_426),
.B(n_386),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_455),
.A2(n_399),
.B1(n_388),
.B2(n_387),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_388),
.B1(n_386),
.B2(n_362),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_455),
.B(n_399),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_477),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_362),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_486),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_442),
.A2(n_409),
.B1(n_399),
.B2(n_362),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_486),
.Y(n_535)
);

AO22x2_ASAP7_75t_L g536 ( 
.A1(n_442),
.A2(n_409),
.B1(n_399),
.B2(n_362),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_412),
.A2(n_409),
.B1(n_399),
.B2(n_5),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_446),
.B(n_409),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_412),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_419),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_456),
.B(n_379),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_272),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

AO22x2_ASAP7_75t_L g545 ( 
.A1(n_419),
.A2(n_430),
.B1(n_444),
.B2(n_429),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_430),
.A2(n_429),
.B1(n_434),
.B2(n_460),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_472),
.A2(n_283),
.B1(n_282),
.B2(n_281),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_478),
.B(n_7),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_449),
.Y(n_554)
);

AO22x2_ASAP7_75t_L g555 ( 
.A1(n_449),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_478),
.A2(n_280),
.B1(n_275),
.B2(n_11),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_415),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_459),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_459),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_461),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_482),
.B(n_247),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_469),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_438),
.B(n_247),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_425),
.B(n_247),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_467),
.B(n_12),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

OAI221xp5_ASAP7_75t_L g570 ( 
.A1(n_471),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.C(n_18),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_569),
.B(n_438),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_504),
.B(n_494),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_568),
.B(n_462),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_504),
.B(n_471),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_494),
.B(n_464),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_441),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_512),
.B(n_441),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_502),
.B(n_415),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_560),
.B(n_418),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_490),
.B(n_418),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_493),
.B(n_463),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_512),
.B(n_441),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_441),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_505),
.B(n_420),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_493),
.B(n_463),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_525),
.B(n_463),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_488),
.B(n_420),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_538),
.B(n_519),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_519),
.B(n_427),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_506),
.B(n_427),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_542),
.B(n_247),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_497),
.B(n_435),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_530),
.B(n_435),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_487),
.B(n_483),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_489),
.B(n_463),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_500),
.B(n_435),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_513),
.B(n_435),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_556),
.B(n_435),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_552),
.B(n_526),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_491),
.B(n_483),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_495),
.B(n_437),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_496),
.B(n_437),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_538),
.B(n_463),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_498),
.B(n_437),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_503),
.B(n_507),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_543),
.B(n_437),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_508),
.B(n_437),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_514),
.B(n_14),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_515),
.B(n_517),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_522),
.B(n_16),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_557),
.B(n_20),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_511),
.B(n_21),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_501),
.B(n_21),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_529),
.B(n_22),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_520),
.B(n_22),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_SL g617 ( 
.A(n_562),
.B(n_23),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_524),
.B(n_24),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_533),
.B(n_24),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_537),
.B(n_468),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_518),
.B(n_25),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_541),
.B(n_492),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_565),
.B(n_25),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_559),
.B(n_26),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_521),
.B(n_26),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_535),
.B(n_27),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_518),
.B(n_27),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_559),
.B(n_28),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_546),
.B(n_28),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_548),
.B(n_29),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_563),
.B(n_29),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_SL g632 ( 
.A(n_566),
.B(n_30),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_564),
.B(n_31),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_527),
.B(n_468),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_571),
.B(n_554),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_561),
.B(n_31),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_532),
.B(n_468),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_528),
.B(n_32),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_622),
.B(n_593),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_581),
.A2(n_549),
.B(n_545),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_615),
.A2(n_567),
.B(n_570),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_531),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_601),
.A2(n_544),
.A3(n_551),
.B(n_550),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_589),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_606),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_637),
.A2(n_547),
.B(n_545),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_635),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_589),
.B(n_499),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_574),
.A2(n_540),
.B(n_537),
.C(n_539),
.Y(n_649)
);

CKINVDCx11_ASAP7_75t_R g650 ( 
.A(n_607),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_607),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_572),
.A2(n_549),
.B(n_536),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_600),
.A2(n_638),
.B(n_628),
.C(n_624),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_604),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_611),
.A2(n_553),
.B(n_468),
.Y(n_655)
);

AO21x2_ASAP7_75t_L g656 ( 
.A1(n_592),
.A2(n_534),
.B(n_536),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_602),
.A2(n_534),
.B(n_540),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_SL g658 ( 
.A(n_575),
.B(n_539),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_573),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_621),
.B(n_499),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_576),
.A2(n_553),
.B(n_555),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_603),
.A2(n_558),
.B(n_555),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_595),
.A2(n_558),
.B(n_510),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_620),
.B(n_516),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_605),
.A2(n_608),
.B(n_598),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_582),
.A2(n_510),
.A3(n_509),
.B(n_516),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_617),
.A2(n_509),
.B(n_468),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_623),
.A2(n_37),
.B(n_38),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_636),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_627),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_596),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_629),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_597),
.A2(n_39),
.B(n_40),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_634),
.A2(n_42),
.B(n_43),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_632),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_620),
.B(n_588),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_585),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_577),
.A2(n_580),
.B(n_586),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_594),
.B(n_48),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_614),
.A2(n_609),
.B(n_616),
.C(n_618),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_579),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_49),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_630),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_631),
.A2(n_58),
.B(n_60),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_587),
.A2(n_62),
.B(n_63),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_599),
.B(n_64),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_633),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_584),
.Y(n_689)
);

AND3x4_ASAP7_75t_L g690 ( 
.A(n_591),
.B(n_68),
.C(n_70),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_578),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_612),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_619),
.A2(n_75),
.B(n_76),
.C(n_78),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_583),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_642),
.A2(n_626),
.B1(n_625),
.B2(n_81),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_639),
.A2(n_79),
.B(n_80),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_663),
.A2(n_82),
.B(n_83),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_645),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_642),
.B(n_208),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_665),
.A2(n_86),
.B(n_87),
.Y(n_700)
);

OA21x2_ASAP7_75t_L g701 ( 
.A1(n_640),
.A2(n_89),
.B(n_90),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_643),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_674),
.A2(n_91),
.B(n_92),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_646),
.A2(n_95),
.B(n_96),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_658),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_653),
.A2(n_107),
.B(n_108),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_647),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_680),
.A2(n_641),
.B(n_649),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_640),
.A2(n_673),
.B(n_686),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_678),
.A2(n_110),
.B(n_111),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_662),
.A2(n_112),
.B(n_113),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_681),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_641),
.A2(n_119),
.B(n_121),
.C(n_122),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_672),
.A2(n_684),
.B1(n_687),
.B2(n_676),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_679),
.A2(n_123),
.B(n_124),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_644),
.B(n_125),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_660),
.B(n_128),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_670),
.B(n_129),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_650),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_643),
.Y(n_720)
);

AOI21xp33_ASAP7_75t_SL g721 ( 
.A1(n_690),
.A2(n_130),
.B(n_131),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_677),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_664),
.A2(n_132),
.B1(n_134),
.B2(n_137),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_694),
.Y(n_724)
);

AO31x2_ASAP7_75t_L g725 ( 
.A1(n_652),
.A2(n_139),
.A3(n_144),
.B(n_145),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_664),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_676),
.B(n_150),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_651),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_659),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_689),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_661),
.A2(n_152),
.B1(n_156),
.B2(n_159),
.Y(n_731)
);

OAI21x1_ASAP7_75t_L g732 ( 
.A1(n_657),
.A2(n_162),
.B(n_165),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_668),
.A2(n_167),
.B(n_168),
.C(n_169),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_648),
.B(n_170),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_651),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_669),
.A2(n_171),
.B(n_174),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_675),
.A2(n_176),
.B(n_177),
.Y(n_737)
);

OA21x2_ASAP7_75t_L g738 ( 
.A1(n_685),
.A2(n_179),
.B(n_181),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_654),
.B(n_207),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

NOR2x1_ASAP7_75t_SL g741 ( 
.A(n_671),
.B(n_183),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_691),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_651),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_682),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_656),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_702),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_702),
.A2(n_667),
.B(n_655),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_709),
.A2(n_692),
.B(n_688),
.Y(n_748)
);

OA21x2_ASAP7_75t_L g749 ( 
.A1(n_709),
.A2(n_655),
.B(n_693),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_744),
.B(n_666),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_708),
.Y(n_751)
);

AO21x2_ASAP7_75t_L g752 ( 
.A1(n_720),
.A2(n_656),
.B(n_688),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_720),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_745),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_744),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_698),
.B(n_666),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_696),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_745),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_745),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_707),
.B(n_727),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_728),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_725),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_697),
.A2(n_683),
.B(n_643),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_711),
.A2(n_683),
.B(n_666),
.Y(n_766)
);

CKINVDCx6p67_ASAP7_75t_R g767 ( 
.A(n_719),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_710),
.A2(n_184),
.B(n_185),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_740),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_725),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_701),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_714),
.A2(n_187),
.B1(n_190),
.B2(n_193),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_725),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_701),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_735),
.B(n_194),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_711),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_728),
.B(n_195),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_732),
.B(n_197),
.Y(n_779)
);

AND2x6_ASAP7_75t_L g780 ( 
.A(n_727),
.B(n_198),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_705),
.A2(n_202),
.B1(n_206),
.B2(n_706),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_722),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_742),
.B(n_743),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_696),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_704),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_724),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_743),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_699),
.B(n_717),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_731),
.B(n_705),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_716),
.B(n_734),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_738),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_721),
.B(n_695),
.Y(n_794)
);

AO31x2_ASAP7_75t_L g795 ( 
.A1(n_713),
.A2(n_733),
.A3(n_741),
.B(n_712),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_710),
.A2(n_737),
.B(n_703),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_738),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_731),
.B(n_726),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_738),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_715),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_723),
.B(n_726),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_787),
.B(n_718),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_R g803 ( 
.A(n_751),
.B(n_739),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_780),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_767),
.Y(n_805)
);

XNOR2xp5_ASAP7_75t_L g806 ( 
.A(n_756),
.B(n_723),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_780),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_780),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_761),
.B(n_713),
.Y(n_809)
);

XNOR2xp5_ASAP7_75t_L g810 ( 
.A(n_756),
.B(n_776),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_756),
.B(n_736),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_R g812 ( 
.A(n_767),
.B(n_733),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_762),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_784),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_761),
.B(n_695),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_762),
.B(n_751),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_784),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_783),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_R g819 ( 
.A(n_801),
.B(n_798),
.Y(n_819)
);

XOR2xp5_ASAP7_75t_L g820 ( 
.A(n_791),
.B(n_750),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_788),
.B(n_791),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_762),
.B(n_788),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_783),
.B(n_789),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_R g824 ( 
.A(n_801),
.B(n_798),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_780),
.B(n_794),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_789),
.B(n_769),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_757),
.B(n_790),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_790),
.B(n_753),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_778),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_780),
.B(n_794),
.Y(n_831)
);

BUFx10_ASAP7_75t_L g832 ( 
.A(n_780),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_753),
.B(n_778),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_778),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_R g835 ( 
.A(n_778),
.B(n_766),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_753),
.B(n_759),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_780),
.B(n_775),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_754),
.B(n_760),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_R g839 ( 
.A(n_766),
.B(n_759),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_752),
.B(n_747),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_754),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_795),
.B(n_781),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_747),
.Y(n_843)
);

CKINVDCx8_ASAP7_75t_R g844 ( 
.A(n_766),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_R g845 ( 
.A(n_749),
.B(n_755),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_747),
.Y(n_846)
);

OAI222xp33_ASAP7_75t_L g847 ( 
.A1(n_815),
.A2(n_781),
.B1(n_773),
.B2(n_764),
.C1(n_770),
.C2(n_763),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_816),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_818),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_827),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_828),
.B(n_793),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_813),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_830),
.B(n_793),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_833),
.B(n_755),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_829),
.B(n_773),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_842),
.B(n_793),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_814),
.B(n_793),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_817),
.B(n_797),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_829),
.B(n_825),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_821),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_829),
.B(n_770),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_836),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_841),
.B(n_752),
.Y(n_863)
);

OR2x2_ASAP7_75t_SL g864 ( 
.A(n_834),
.B(n_749),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_805),
.B(n_800),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_836),
.B(n_797),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_823),
.B(n_810),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_822),
.B(n_752),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_820),
.B(n_752),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_838),
.Y(n_870)
);

AOI221xp5_ASAP7_75t_L g871 ( 
.A1(n_809),
.A2(n_764),
.B1(n_763),
.B2(n_799),
.C(n_772),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_838),
.B(n_799),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_811),
.B(n_747),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_844),
.B(n_777),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_R g875 ( 
.A(n_803),
.B(n_765),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_843),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_840),
.B(n_846),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_804),
.B(n_777),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_840),
.B(n_746),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_871),
.A2(n_824),
.B1(n_819),
.B2(n_806),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_851),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_852),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_850),
.B(n_837),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_847),
.B(n_748),
.C(n_758),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_876),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_848),
.A2(n_812),
.B1(n_826),
.B2(n_831),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_869),
.A2(n_808),
.B1(n_832),
.B2(n_804),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_851),
.B(n_808),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_877),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_877),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_879),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_879),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_852),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_860),
.B(n_802),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_853),
.B(n_832),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_874),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_848),
.Y(n_897)
);

OAI31xp33_ASAP7_75t_SL g898 ( 
.A1(n_856),
.A2(n_748),
.A3(n_835),
.B(n_807),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_873),
.B(n_746),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_875),
.B(n_807),
.Y(n_900)
);

OAI31xp33_ASAP7_75t_L g901 ( 
.A1(n_867),
.A2(n_779),
.A3(n_782),
.B(n_771),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_897),
.B(n_859),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_856),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_896),
.B(n_859),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_891),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_896),
.B(n_853),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_883),
.B(n_858),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_885),
.Y(n_908)
);

AND3x2_ASAP7_75t_L g909 ( 
.A(n_898),
.B(n_874),
.C(n_863),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_881),
.B(n_872),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_896),
.B(n_872),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_882),
.B(n_857),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_888),
.B(n_857),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_888),
.B(n_858),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_868),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_908),
.Y(n_916)
);

OAI221xp5_ASAP7_75t_L g917 ( 
.A1(n_915),
.A2(n_880),
.B1(n_901),
.B2(n_884),
.C(n_887),
.Y(n_917)
);

NOR2x1_ASAP7_75t_L g918 ( 
.A(n_903),
.B(n_894),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_907),
.B(n_889),
.Y(n_919)
);

NAND2xp33_ASAP7_75t_SL g920 ( 
.A(n_903),
.B(n_882),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_914),
.B(n_890),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_910),
.B(n_890),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_905),
.Y(n_923)
);

NOR2x1_ASAP7_75t_L g924 ( 
.A(n_918),
.B(n_902),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_921),
.B(n_904),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_916),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_919),
.B(n_922),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_923),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_917),
.B(n_885),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_920),
.Y(n_930)
);

XNOR2xp5_ASAP7_75t_L g931 ( 
.A(n_924),
.B(n_880),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_926),
.B(n_914),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_924),
.B(n_886),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_929),
.A2(n_904),
.B(n_906),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_928),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_932),
.B(n_925),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_935),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_933),
.B(n_930),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_937),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_938),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_936),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_937),
.Y(n_942)
);

OA22x2_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_931),
.B1(n_934),
.B2(n_909),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_SL g944 ( 
.A(n_942),
.B(n_927),
.C(n_901),
.Y(n_944)
);

AOI211xp5_ASAP7_75t_L g945 ( 
.A1(n_940),
.A2(n_900),
.B(n_893),
.C(n_909),
.Y(n_945)
);

NOR5xp2_ASAP7_75t_L g946 ( 
.A(n_939),
.B(n_870),
.C(n_786),
.D(n_862),
.E(n_865),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_941),
.B(n_911),
.Y(n_947)
);

AOI211xp5_ASAP7_75t_L g948 ( 
.A1(n_944),
.A2(n_895),
.B(n_878),
.C(n_912),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_945),
.B(n_768),
.C(n_765),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_947),
.B(n_913),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_943),
.B(n_768),
.C(n_899),
.Y(n_951)
);

AOI211xp5_ASAP7_75t_SL g952 ( 
.A1(n_946),
.A2(n_758),
.B(n_786),
.C(n_800),
.Y(n_952)
);

AND3x4_ASAP7_75t_L g953 ( 
.A(n_949),
.B(n_863),
.C(n_892),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_950),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_952),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_951),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_948),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_957),
.B(n_758),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_891),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_SL g960 ( 
.A(n_956),
.B(n_800),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_953),
.B(n_845),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_954),
.B(n_839),
.C(n_862),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_SL g963 ( 
.A(n_959),
.B(n_779),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_958),
.B(n_866),
.Y(n_964)
);

XNOR2x1_ASAP7_75t_L g965 ( 
.A(n_960),
.B(n_863),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_SL g966 ( 
.A1(n_962),
.A2(n_792),
.B(n_749),
.Y(n_966)
);

XNOR2xp5_ASAP7_75t_L g967 ( 
.A(n_961),
.B(n_864),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_963),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_964),
.B(n_795),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_968),
.A2(n_967),
.B1(n_966),
.B2(n_965),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_971),
.A2(n_849),
.B1(n_749),
.B2(n_785),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_972),
.A2(n_970),
.B1(n_785),
.B2(n_849),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_973),
.A2(n_796),
.B1(n_774),
.B2(n_782),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_973),
.A2(n_796),
.B(n_861),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_975),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_976),
.A2(n_974),
.B1(n_774),
.B2(n_782),
.C(n_771),
.Y(n_977)
);

AOI211xp5_ASAP7_75t_L g978 ( 
.A1(n_977),
.A2(n_855),
.B(n_795),
.C(n_854),
.Y(n_978)
);


endmodule