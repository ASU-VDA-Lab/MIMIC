module fake_netlist_6_2962_n_170 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_170);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_170;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_151;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_2),
.C(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_28),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_8),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_45),
.B(n_41),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_39),
.B(n_33),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_37),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_62),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_48),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_42),
.C(n_41),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_34),
.B(n_50),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_59),
.B(n_67),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_18),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_57),
.B1(n_69),
.B2(n_64),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_58),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_87),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_71),
.B(n_75),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_61),
.B(n_72),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_61),
.B(n_72),
.C(n_70),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_74),
.B1(n_44),
.B2(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_71),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_58),
.B(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_83),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_82),
.Y(n_112)
);

OAI221xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_93),
.B1(n_101),
.B2(n_86),
.C(n_97),
.Y(n_113)
);

OAI221xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_82),
.B1(n_79),
.B2(n_99),
.C(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_99),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_95),
.C(n_88),
.Y(n_117)
);

OAI221xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_90),
.B1(n_68),
.B2(n_56),
.C(n_59),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_104),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_107),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_111),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_114),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_113),
.B1(n_107),
.B2(n_106),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_109),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_109),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

OAI222xp33_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_118),
.B1(n_67),
.B2(n_60),
.C1(n_65),
.C2(n_68),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_108),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_65),
.C(n_130),
.Y(n_142)
);

NAND4xp25_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_124),
.C(n_136),
.D(n_125),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_133),
.Y(n_144)
);

NAND4xp25_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_133),
.C(n_131),
.D(n_128),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_134),
.C(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_134),
.Y(n_147)
);

NAND4xp25_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_109),
.C(n_92),
.D(n_14),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_89),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_137),
.B1(n_135),
.B2(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_71),
.B1(n_88),
.B2(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_142),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_153),
.B1(n_156),
.B2(n_155),
.C(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_160),
.C(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

NAND2x1p5_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_162),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_167),
.B1(n_168),
.B2(n_162),
.C(n_110),
.Y(n_170)
);


endmodule