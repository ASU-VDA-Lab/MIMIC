module fake_jpeg_4627_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_21),
.B1(n_17),
.B2(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_22),
.B1(n_12),
.B2(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_12),
.B1(n_23),
.B2(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_36),
.B1(n_21),
.B2(n_24),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_46),
.C(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_28),
.B1(n_14),
.B2(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_28),
.C(n_29),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_41),
.C(n_57),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_6),
.C(n_8),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_42),
.C(n_7),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_45),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_50),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_79),
.B(n_62),
.Y(n_82)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_29),
.C(n_20),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_69),
.B1(n_59),
.B2(n_64),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_79),
.B(n_65),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_90),
.C(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_84),
.B1(n_69),
.B2(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_77),
.C(n_61),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_78),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_99),
.B(n_1),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_83),
.B1(n_67),
.B2(n_20),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_5),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_5),
.B1(n_8),
.B2(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_99),
.C(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

AO21x2_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);


endmodule