module real_jpeg_12106_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_292, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_292;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_215;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_29),
.B1(n_32),
.B2(n_45),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_4),
.A2(n_45),
.B1(n_71),
.B2(n_72),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_71),
.B1(n_72),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_132),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_132),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_132),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_53),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_31),
.B1(n_71),
.B2(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_7),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_7),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_10),
.A2(n_70),
.B(n_71),
.C(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_10),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_81),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_146),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_99),
.B1(n_100),
.B2(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_10),
.B(n_87),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_71),
.B1(n_72),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_11),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_155),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_155),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_155),
.Y(n_234)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_13),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_36),
.B1(n_71),
.B2(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_71),
.B1(n_72),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_79),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_79),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_79),
.Y(n_228)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_270),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_133),
.B(n_269),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_19),
.B(n_113),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_83),
.B2(n_112),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_20),
.B(n_84),
.C(n_96),
.Y(n_272)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_66),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_22),
.A2(n_23),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_26),
.A2(n_99),
.B(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_27),
.A2(n_37),
.B1(n_123),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_27),
.A2(n_37),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_28),
.A2(n_37),
.B(n_125),
.Y(n_199)
);

CKINVDCx6p67_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_32),
.B(n_49),
.C(n_146),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_32),
.B(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_33),
.A2(n_100),
.B(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_50),
.B(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_42),
.A2(n_56),
.B(n_196),
.C(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_42),
.B(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_43),
.B(n_57),
.C(n_59),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_52),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_46),
.A2(n_91),
.B(n_104),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_46),
.A2(n_51),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_46),
.A2(n_51),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_46),
.A2(n_51),
.B1(n_211),
.B2(n_221),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_46),
.A2(n_51),
.B(n_91),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_50),
.B(n_146),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_66),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_61),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_55),
.A2(n_150),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_60),
.B1(n_70),
.B2(n_75),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_59),
.A2(n_75),
.B(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g197 ( 
.A(n_60),
.B(n_146),
.CON(n_197),
.SN(n_197)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_62),
.A2(n_87),
.B1(n_149),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_62),
.A2(n_87),
.B1(n_184),
.B2(n_197),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_77),
.B(n_80),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_67),
.A2(n_76),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_78),
.B1(n_81),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_68),
.A2(n_81),
.B1(n_154),
.B2(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_68),
.B(n_111),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_69)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_76),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_96),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_95),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_128),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_88),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_90),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_95),
.B(n_274),
.CI(n_275),
.CON(n_273),
.SN(n_273)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_97),
.A2(n_98),
.B(n_107),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_99),
.A2(n_100),
.B1(n_226),
.B2(n_234),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_100),
.B(n_146),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_118),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_119),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_126),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_130),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_129),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_263),
.B(n_268),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_172),
.B1(n_188),
.B2(n_262),
.C(n_292),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_161),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_136),
.B(n_161),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_157),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_137),
.B(n_158),
.C(n_159),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.C(n_152),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_139),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B(n_151),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_150),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_171),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_186),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_173),
.B(n_186),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_174),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_178),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_182),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_261),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_256),
.B(n_260),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_212),
.B(n_255),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_207),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_192),
.B(n_207),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_200),
.C(n_204),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_199),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_210),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_250),
.B(n_254),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_240),
.B(n_249),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_229),
.B(n_239),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_222),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_288),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_273),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_273),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_284),
.B2(n_287),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);


endmodule