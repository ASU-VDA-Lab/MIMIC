module real_jpeg_28299_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_44),
.B(n_45),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_11),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_13),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_12),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OR2x2_ASAP7_75t_SL g18 ( 
.A(n_5),
.B(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_5),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

OAI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_16),
.B(n_25),
.C(n_42),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_12),
.B(n_13),
.Y(n_9)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_32),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_31),
.Y(n_44)
);

AOI221xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);


endmodule