module real_aes_238_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_746;
wire n_656;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_996;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_449;
wire n_754;
wire n_417;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_727;
wire n_649;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_0), .A2(n_166), .B1(n_790), .B2(n_791), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_1), .A2(n_132), .B1(n_457), .B2(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_2), .A2(n_206), .B1(n_520), .B2(n_521), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_3), .A2(n_122), .B1(n_457), .B2(n_507), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_4), .A2(n_15), .B1(n_461), .B2(n_505), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_5), .A2(n_121), .B1(n_603), .B2(n_678), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_6), .A2(n_105), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_7), .A2(n_336), .B1(n_446), .B2(n_449), .Y(n_445) );
AOI22xp5_ASAP7_75t_SL g562 ( .A1(n_8), .A2(n_373), .B1(n_504), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_9), .A2(n_259), .B1(n_615), .B2(n_694), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_10), .B(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_11), .A2(n_75), .B1(n_498), .B2(n_557), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_12), .A2(n_93), .B1(n_472), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_13), .A2(n_172), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_14), .A2(n_313), .B1(n_442), .B2(n_551), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_16), .A2(n_131), .B1(n_457), .B2(n_507), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_17), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g866 ( .A1(n_18), .A2(n_170), .B1(n_191), .B2(n_681), .C1(n_684), .C2(n_867), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_19), .A2(n_357), .B1(n_784), .B2(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_20), .A2(n_177), .B1(n_502), .B2(n_603), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_21), .A2(n_221), .B1(n_538), .B2(n_539), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g751 ( .A1(n_22), .A2(n_119), .B1(n_277), .B2(n_752), .C1(n_753), .C2(n_754), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_23), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_24), .A2(n_354), .B1(n_498), .B2(n_592), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_25), .A2(n_80), .B1(n_605), .B2(n_606), .Y(n_918) );
AOI222xp33_ASAP7_75t_L g768 ( .A1(n_26), .A2(n_335), .B1(n_366), .B2(n_457), .C1(n_565), .C2(n_752), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_27), .A2(n_291), .B1(n_592), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_28), .A2(n_289), .B1(n_399), .B2(n_419), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_29), .A2(n_37), .B1(n_454), .B2(n_457), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_30), .A2(n_229), .B1(n_548), .B2(n_673), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_31), .A2(n_96), .B1(n_181), .B2(n_517), .C1(n_518), .C2(n_524), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_32), .A2(n_240), .B1(n_780), .B2(n_784), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_33), .A2(n_230), .B1(n_517), .B2(n_606), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_34), .A2(n_42), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_35), .A2(n_231), .B1(n_791), .B2(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g417 ( .A(n_36), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_36), .B(n_48), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_38), .A2(n_67), .B1(n_539), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_39), .A2(n_379), .B1(n_488), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_40), .A2(n_147), .B1(n_502), .B2(n_603), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_41), .A2(n_97), .B1(n_454), .B2(n_457), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_43), .A2(n_368), .B1(n_551), .B2(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_44), .A2(n_83), .B1(n_563), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_45), .A2(n_68), .B1(n_421), .B2(n_585), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_46), .A2(n_258), .B1(n_488), .B2(n_651), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_47), .A2(n_383), .B1(n_390), .B2(n_948), .C(n_958), .Y(n_382) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_48), .A2(n_355), .B1(n_406), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_49), .A2(n_249), .B1(n_421), .B2(n_693), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_50), .A2(n_276), .B1(n_457), .B2(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_51), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_52), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_53), .A2(n_363), .B1(n_502), .B2(n_628), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_54), .A2(n_239), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_55), .A2(n_87), .B1(n_502), .B2(n_802), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_56), .A2(n_281), .B1(n_548), .B2(n_673), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_57), .A2(n_349), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_58), .A2(n_282), .B1(n_632), .B2(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g418 ( .A(n_59), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_60), .A2(n_237), .B1(n_443), .B2(n_790), .Y(n_825) );
AO22x1_ASAP7_75t_L g907 ( .A1(n_61), .A2(n_167), .B1(n_649), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_62), .A2(n_228), .B1(n_697), .B2(n_741), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_63), .A2(n_247), .B1(n_438), .B2(n_535), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_64), .B(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_65), .A2(n_114), .B1(n_605), .B2(n_606), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_66), .A2(n_136), .B1(n_442), .B2(n_790), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_69), .A2(n_356), .B1(n_548), .B2(n_673), .Y(n_759) );
AOI222xp33_ASAP7_75t_L g656 ( .A1(n_70), .A2(n_212), .B1(n_241), .B2(n_657), .C1(n_658), .C2(n_661), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_71), .A2(n_234), .B1(n_619), .B2(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_72), .B(n_478), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_73), .A2(n_150), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_74), .A2(n_252), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_76), .A2(n_341), .B1(n_421), .B2(n_548), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_77), .A2(n_124), .B1(n_594), .B2(n_675), .Y(n_871) );
AO22x2_ASAP7_75t_L g405 ( .A1(n_78), .A2(n_187), .B1(n_406), .B2(n_407), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_79), .A2(n_193), .B1(n_433), .B2(n_437), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_81), .A2(n_350), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_82), .A2(n_205), .B1(n_778), .B2(n_780), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_84), .A2(n_251), .B1(n_548), .B2(n_906), .Y(n_905) );
XOR2xp5_ASAP7_75t_L g642 ( .A(n_85), .B(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_86), .A2(n_176), .B1(n_541), .B2(n_542), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_88), .A2(n_137), .B1(n_443), .B2(n_554), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_89), .A2(n_246), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_90), .A2(n_338), .B1(n_491), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_91), .A2(n_371), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_92), .A2(n_260), .B1(n_449), .B2(n_787), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_94), .A2(n_158), .B1(n_472), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_95), .A2(n_129), .B1(n_555), .B2(n_787), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_98), .A2(n_342), .B1(n_541), .B2(n_542), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_99), .A2(n_286), .B1(n_477), .B2(n_931), .Y(n_978) );
XOR2x2_ASAP7_75t_L g665 ( .A(n_100), .B(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_101), .A2(n_333), .B1(n_554), .B2(n_619), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_102), .A2(n_199), .B1(n_532), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_103), .A2(n_154), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_104), .A2(n_321), .B1(n_434), .B2(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_106), .B(n_776), .Y(n_775) );
OA22x2_ASAP7_75t_L g839 ( .A1(n_107), .A2(n_840), .B1(n_841), .B2(n_856), .Y(n_839) );
INVx1_ASAP7_75t_L g856 ( .A(n_107), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_108), .A2(n_248), .B1(n_489), .B2(n_557), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_109), .A2(n_267), .B1(n_526), .B2(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_110), .B(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_111), .A2(n_378), .B1(n_504), .B2(n_628), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_112), .A2(n_178), .B1(n_541), .B2(n_542), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_113), .A2(n_200), .B1(n_457), .B2(n_565), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_115), .A2(n_347), .B1(n_791), .B2(n_829), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_116), .A2(n_194), .B1(n_502), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_117), .A2(n_207), .B1(n_651), .B2(n_675), .Y(n_674) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_118), .A2(n_294), .B1(n_406), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_120), .A2(n_370), .B1(n_449), .B2(n_787), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_123), .A2(n_364), .B1(n_488), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_125), .A2(n_375), .B1(n_554), .B2(n_555), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_126), .A2(n_144), .B1(n_446), .B2(n_649), .Y(n_1006) );
OA22x2_ASAP7_75t_L g736 ( .A1(n_127), .A2(n_737), .B1(n_738), .B2(n_755), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_127), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_128), .A2(n_222), .B1(n_443), .B2(n_557), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g843 ( .A1(n_130), .A2(n_226), .B1(n_274), .B2(n_778), .C1(n_822), .C2(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_133), .B(n_561), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_134), .A2(n_263), .B1(n_526), .B2(n_754), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_135), .B(n_684), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_138), .A2(n_293), .B1(n_551), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_139), .A2(n_305), .B1(n_437), .B2(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_140), .A2(n_369), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_141), .A2(n_209), .B1(n_494), .B2(n_549), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_142), .A2(n_362), .B1(n_470), .B2(n_472), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_143), .A2(n_253), .B1(n_457), .B2(n_565), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_145), .A2(n_367), .B1(n_628), .B2(n_965), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_146), .A2(n_197), .B1(n_520), .B2(n_521), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_148), .A2(n_211), .B1(n_520), .B2(n_521), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_149), .A2(n_244), .B1(n_531), .B2(n_532), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_151), .A2(n_273), .B1(n_437), .B2(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_152), .A2(n_162), .B1(n_551), .B2(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_153), .A2(n_332), .B1(n_504), .B2(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_155), .A2(n_284), .B1(n_491), .B2(n_492), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_156), .A2(n_268), .B1(n_425), .B2(n_433), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_157), .A2(n_326), .B1(n_538), .B2(n_539), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_159), .A2(n_265), .B1(n_438), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_160), .A2(n_208), .B1(n_491), .B2(n_974), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_161), .A2(n_215), .B1(n_497), .B2(n_654), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_163), .A2(n_233), .B1(n_421), .B2(n_548), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_164), .A2(n_352), .B1(n_517), .B2(n_606), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g847 ( .A1(n_165), .A2(n_192), .B1(n_632), .B2(n_820), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_168), .A2(n_960), .B1(n_961), .B2(n_979), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_168), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_169), .A2(n_287), .B1(n_681), .B2(n_709), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_171), .A2(n_214), .B1(n_526), .B2(n_527), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_173), .A2(n_175), .B1(n_470), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_174), .A2(n_198), .B1(n_427), .B2(n_697), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_179), .A2(n_182), .B1(n_494), .B2(n_495), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_180), .A2(n_306), .B1(n_669), .B2(n_747), .Y(n_872) );
INVx1_ASAP7_75t_L g634 ( .A(n_183), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_184), .A2(n_328), .B1(n_605), .B2(n_606), .Y(n_604) );
OA22x2_ASAP7_75t_L g875 ( .A1(n_185), .A2(n_876), .B1(n_877), .B2(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_185), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_186), .A2(n_325), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g956 ( .A(n_187), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_188), .A2(n_323), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_189), .A2(n_256), .B1(n_526), .B2(n_527), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_190), .A2(n_318), .B1(n_541), .B2(n_542), .Y(n_923) );
INVx1_ASAP7_75t_L g863 ( .A(n_195), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_196), .A2(n_381), .B1(n_693), .B2(n_694), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_201), .A2(n_262), .B1(n_464), .B2(n_778), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_202), .A2(n_250), .B1(n_654), .B2(n_671), .Y(n_670) );
OAI22x1_ASAP7_75t_SL g772 ( .A1(n_203), .A2(n_773), .B1(n_793), .B2(n_794), .Y(n_772) );
INVx1_ASAP7_75t_L g793 ( .A(n_203), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_204), .A2(n_264), .B1(n_746), .B2(n_747), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_210), .A2(n_307), .B1(n_632), .B2(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_213), .B(n_657), .Y(n_920) );
XNOR2x1_ASAP7_75t_L g982 ( .A(n_216), .B(n_983), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_216), .Y(n_1013) );
AO22x2_ASAP7_75t_L g813 ( .A1(n_217), .A2(n_814), .B1(n_815), .B2(n_830), .Y(n_813) );
INVx1_ASAP7_75t_L g830 ( .A(n_217), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_218), .A2(n_242), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g894 ( .A(n_219), .Y(n_894) );
INVx2_ASAP7_75t_L g389 ( .A(n_220), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_223), .A2(n_279), .B1(n_531), .B2(n_532), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_224), .A2(n_308), .B1(n_437), .B2(n_441), .Y(n_436) );
OA22x2_ASAP7_75t_L g608 ( .A1(n_225), .A2(n_609), .B1(n_610), .B2(n_638), .Y(n_608) );
INVx1_ASAP7_75t_L g638 ( .A(n_225), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_227), .A2(n_317), .B1(n_681), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_232), .A2(n_330), .B1(n_681), .B2(n_867), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_235), .A2(n_243), .B1(n_551), .B2(n_697), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_236), .A2(n_346), .B1(n_592), .B2(n_697), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_238), .A2(n_275), .B1(n_761), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_245), .A2(n_288), .B1(n_457), .B2(n_507), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_254), .A2(n_309), .B1(n_534), .B2(n_535), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_255), .B(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_257), .A2(n_324), .B1(n_520), .B2(n_521), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_261), .A2(n_299), .B1(n_502), .B2(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_266), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_269), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_270), .A2(n_339), .B1(n_419), .B2(n_615), .Y(n_788) );
INVx1_ASAP7_75t_L g633 ( .A(n_271), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_272), .B(n_457), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_278), .B(n_776), .Y(n_817) );
AO22x1_ASAP7_75t_L g927 ( .A1(n_280), .A2(n_928), .B1(n_942), .B2(n_943), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_280), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_283), .Y(n_989) );
XNOR2x1_ASAP7_75t_L g395 ( .A(n_285), .B(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_290), .A2(n_353), .B1(n_673), .B2(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_292), .A2(n_343), .B1(n_538), .B2(n_539), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_294), .B(n_955), .Y(n_954) );
OA22x2_ASAP7_75t_L g798 ( .A1(n_295), .A2(n_799), .B1(n_811), .B2(n_812), .Y(n_798) );
INVx1_ASAP7_75t_L g811 ( .A(n_295), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_296), .A2(n_337), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_297), .A2(n_377), .B1(n_461), .B2(n_464), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_298), .A2(n_348), .B1(n_489), .B2(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_300), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_301), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_302), .A2(n_358), .B1(n_628), .B2(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_303), .B(n_684), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_304), .A2(n_345), .B1(n_442), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_310), .A2(n_329), .B1(n_563), .B2(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g406 ( .A(n_311), .Y(n_406) );
XNOR2x2_ASAP7_75t_L g914 ( .A(n_312), .B(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_314), .A2(n_334), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g637 ( .A(n_315), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_316), .B(n_477), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g995 ( .A(n_319), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_320), .A2(n_340), .B1(n_495), .B2(n_615), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_322), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_327), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_331), .B(n_478), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_344), .A2(n_380), .B1(n_538), .B2(n_539), .Y(n_922) );
XNOR2x1_ASAP7_75t_L g484 ( .A(n_351), .B(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_359), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_360), .A2(n_374), .B1(n_504), .B2(n_505), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_361), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g952 ( .A(n_361), .Y(n_952) );
INVx1_ASAP7_75t_L g386 ( .A(n_365), .Y(n_386) );
AND2x2_ASAP7_75t_R g981 ( .A(n_365), .B(n_952), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_372), .B(n_388), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_376), .Y(n_992) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_385), .B(n_387), .Y(n_1012) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_386), .B(n_952), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_730), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g948 ( .A1(n_392), .A2(n_731), .B(n_949), .Y(n_948) );
XNOR2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_575), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_481), .B1(n_573), .B2(n_574), .Y(n_393) );
INVxp67_ASAP7_75t_L g573 ( .A(n_394), .Y(n_573) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_452), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_424), .C(n_436), .D(n_445), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_401), .Y(n_494) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g585 ( .A(n_402), .Y(n_585) );
INVx1_ASAP7_75t_L g693 ( .A(n_402), .Y(n_693) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_403), .Y(n_548) );
BUFx3_ASAP7_75t_L g851 ( .A(n_403), .Y(n_851) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_411), .Y(n_403) );
AND2x4_ASAP7_75t_L g451 ( .A(n_404), .B(n_435), .Y(n_451) );
AND2x2_ASAP7_75t_L g471 ( .A(n_404), .B(n_431), .Y(n_471) );
AND2x4_ASAP7_75t_L g520 ( .A(n_404), .B(n_431), .Y(n_520) );
AND2x2_ASAP7_75t_L g531 ( .A(n_404), .B(n_411), .Y(n_531) );
AND2x6_ASAP7_75t_L g539 ( .A(n_404), .B(n_435), .Y(n_539) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_404), .B(n_411), .Y(n_717) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_405), .B(n_409), .Y(n_423) );
INVx2_ASAP7_75t_L g430 ( .A(n_405), .Y(n_430) );
INVx1_ASAP7_75t_L g407 ( .A(n_406), .Y(n_407) );
INVx2_ASAP7_75t_L g410 ( .A(n_406), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_406), .Y(n_413) );
OAI22x1_ASAP7_75t_L g415 ( .A1(n_406), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_406), .Y(n_416) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g429 ( .A(n_409), .Y(n_429) );
AND2x4_ASAP7_75t_L g444 ( .A(n_409), .B(n_430), .Y(n_444) );
AND2x2_ASAP7_75t_L g448 ( .A(n_411), .B(n_428), .Y(n_448) );
AND2x4_ASAP7_75t_L g463 ( .A(n_411), .B(n_444), .Y(n_463) );
AND2x2_ASAP7_75t_L g517 ( .A(n_411), .B(n_444), .Y(n_517) );
AND2x6_ASAP7_75t_L g538 ( .A(n_411), .B(n_428), .Y(n_538) );
AND2x2_ASAP7_75t_L g605 ( .A(n_411), .B(n_444), .Y(n_605) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
BUFx2_ASAP7_75t_L g422 ( .A(n_412), .Y(n_422) );
INVx2_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
AND2x2_ASAP7_75t_L g468 ( .A(n_412), .B(n_415), .Y(n_468) );
AND2x4_ASAP7_75t_L g435 ( .A(n_414), .B(n_432), .Y(n_435) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g431 ( .A(n_415), .B(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g549 ( .A(n_420), .Y(n_549) );
INVx2_ASAP7_75t_L g694 ( .A(n_420), .Y(n_694) );
INVx2_ASAP7_75t_L g906 ( .A(n_420), .Y(n_906) );
INVx5_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
BUFx2_ASAP7_75t_L g586 ( .A(n_421), .Y(n_586) );
BUFx3_ASAP7_75t_L g673 ( .A(n_421), .Y(n_673) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
AND2x4_ASAP7_75t_L g532 ( .A(n_422), .B(n_423), .Y(n_532) );
AND2x4_ASAP7_75t_L g434 ( .A(n_423), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g458 ( .A(n_423), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_423), .B(n_459), .Y(n_527) );
AND2x4_ASAP7_75t_L g542 ( .A(n_423), .B(n_435), .Y(n_542) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_423), .B(n_459), .Y(n_754) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g488 ( .A(n_426), .Y(n_488) );
INVx3_ASAP7_75t_L g557 ( .A(n_426), .Y(n_557) );
INVx2_ASAP7_75t_L g671 ( .A(n_426), .Y(n_671) );
INVx1_ASAP7_75t_SL g829 ( .A(n_426), .Y(n_829) );
INVx6_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g592 ( .A(n_427), .Y(n_592) );
BUFx3_ASAP7_75t_L g741 ( .A(n_427), .Y(n_741) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
AND2x4_ASAP7_75t_L g440 ( .A(n_428), .B(n_435), .Y(n_440) );
AND2x2_ASAP7_75t_L g480 ( .A(n_428), .B(n_468), .Y(n_480) );
AND2x4_ASAP7_75t_L g524 ( .A(n_428), .B(n_468), .Y(n_524) );
AND2x2_ASAP7_75t_L g534 ( .A(n_428), .B(n_435), .Y(n_534) );
AND2x2_ASAP7_75t_L g541 ( .A(n_428), .B(n_431), .Y(n_541) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVxp67_ASAP7_75t_L g467 ( .A(n_430), .Y(n_467) );
AND2x2_ASAP7_75t_L g456 ( .A(n_431), .B(n_444), .Y(n_456) );
AND2x4_ASAP7_75t_L g526 ( .A(n_431), .B(n_444), .Y(n_526) );
BUFx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
BUFx3_ASAP7_75t_L g558 ( .A(n_434), .Y(n_558) );
BUFx3_ASAP7_75t_L g697 ( .A(n_434), .Y(n_697) );
BUFx2_ASAP7_75t_SL g971 ( .A(n_434), .Y(n_971) );
AND2x4_ASAP7_75t_L g443 ( .A(n_435), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g535 ( .A(n_435), .B(n_444), .Y(n_535) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g497 ( .A(n_439), .Y(n_497) );
INVx3_ASAP7_75t_L g551 ( .A(n_439), .Y(n_551) );
INVx2_ASAP7_75t_SL g675 ( .A(n_439), .Y(n_675) );
INVx3_ASAP7_75t_SL g761 ( .A(n_439), .Y(n_761) );
INVx2_ASAP7_75t_L g790 ( .A(n_439), .Y(n_790) );
INVx8_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g622 ( .A(n_442), .Y(n_622) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g489 ( .A(n_443), .Y(n_489) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_443), .Y(n_552) );
INVx2_ASAP7_75t_L g595 ( .A(n_443), .Y(n_595) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_443), .Y(n_941) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g491 ( .A(n_447), .Y(n_491) );
INVx2_ASAP7_75t_L g554 ( .A(n_447), .Y(n_554) );
INVx3_ASAP7_75t_L g618 ( .A(n_447), .Y(n_618) );
INVx2_ASAP7_75t_L g908 ( .A(n_447), .Y(n_908) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g669 ( .A(n_448), .Y(n_669) );
BUFx2_ASAP7_75t_L g746 ( .A(n_448), .Y(n_746) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g492 ( .A(n_450), .Y(n_492) );
INVx2_ASAP7_75t_L g555 ( .A(n_450), .Y(n_555) );
INVx2_ASAP7_75t_L g619 ( .A(n_450), .Y(n_619) );
INVx2_ASAP7_75t_SL g649 ( .A(n_450), .Y(n_649) );
INVx2_ASAP7_75t_SL g699 ( .A(n_450), .Y(n_699) );
INVx2_ASAP7_75t_L g747 ( .A(n_450), .Y(n_747) );
INVx2_ASAP7_75t_L g974 ( .A(n_450), .Y(n_974) );
INVx8_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .C(n_469), .D(n_476), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g704 ( .A(n_455), .Y(n_704) );
INVx2_ASAP7_75t_L g931 ( .A(n_455), .Y(n_931) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx5_ASAP7_75t_L g507 ( .A(n_456), .Y(n_507) );
BUFx3_ASAP7_75t_L g565 ( .A(n_456), .Y(n_565) );
BUFx3_ASAP7_75t_L g660 ( .A(n_456), .Y(n_660) );
INVx2_ASAP7_75t_L g636 ( .A(n_457), .Y(n_636) );
BUFx12f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g567 ( .A(n_458), .Y(n_567) );
BUFx4f_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g996 ( .A(n_462), .Y(n_996) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
BUFx3_ASAP7_75t_L g681 ( .A(n_463), .Y(n_681) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g505 ( .A(n_465), .Y(n_505) );
INVx1_ASAP7_75t_L g563 ( .A(n_465), .Y(n_563) );
INVx2_ASAP7_75t_L g709 ( .A(n_465), .Y(n_709) );
INVx2_ASAP7_75t_L g780 ( .A(n_465), .Y(n_780) );
INVx2_ASAP7_75t_SL g867 ( .A(n_465), .Y(n_867) );
INVx2_ASAP7_75t_L g933 ( .A(n_465), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_465), .A2(n_995), .B1(n_996), .B2(n_997), .Y(n_994) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g518 ( .A(n_467), .B(n_468), .Y(n_518) );
AND2x2_ASAP7_75t_L g606 ( .A(n_467), .B(n_468), .Y(n_606) );
AND2x4_ASAP7_75t_L g473 ( .A(n_468), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g521 ( .A(n_468), .B(n_474), .Y(n_521) );
BUFx6f_ASAP7_75t_SL g784 ( .A(n_470), .Y(n_784) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_471), .Y(n_502) );
INVx3_ASAP7_75t_L g679 ( .A(n_471), .Y(n_679) );
INVxp67_ASAP7_75t_L g993 ( .A(n_472), .Y(n_993) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g570 ( .A(n_473), .Y(n_570) );
BUFx6f_ASAP7_75t_SL g603 ( .A(n_473), .Y(n_603) );
INVx2_ASAP7_75t_L g629 ( .A(n_473), .Y(n_629) );
BUFx3_ASAP7_75t_L g802 ( .A(n_473), .Y(n_802) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g635 ( .A(n_477), .Y(n_635) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g845 ( .A(n_478), .Y(n_845) );
INVx3_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx4_ASAP7_75t_SL g561 ( .A(n_479), .Y(n_561) );
INVx4_ASAP7_75t_SL g657 ( .A(n_479), .Y(n_657) );
INVx3_ASAP7_75t_L g684 ( .A(n_479), .Y(n_684) );
INVx6_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g574 ( .A(n_481), .Y(n_574) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AO22x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_509), .B2(n_510), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_500), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .C(n_493), .D(n_496), .Y(n_486) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g654 ( .A(n_499), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_506), .D(n_508), .Y(n_500) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_502), .Y(n_626) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OA22x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_544), .B2(n_572), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
XOR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_543), .Y(n_512) );
NAND2x1_ASAP7_75t_SL g513 ( .A(n_514), .B(n_528), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx2_ASAP7_75t_SL g598 ( .A(n_524), .Y(n_598) );
BUFx2_ASAP7_75t_L g752 ( .A(n_524), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_526), .Y(n_753) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_536), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_533), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g589 ( .A(n_538), .Y(n_589) );
INVx1_ASAP7_75t_SL g572 ( .A(n_544), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_571), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_559), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_553), .D(n_556), .Y(n_546) );
INVx1_ASAP7_75t_L g1005 ( .A(n_552), .Y(n_1005) );
NAND4xp25_ASAP7_75t_SL g559 ( .A(n_560), .B(n_562), .C(n_564), .D(n_568), .Y(n_559) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_565), .Y(n_632) );
BUFx2_ASAP7_75t_L g820 ( .A(n_566), .Y(n_820) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g661 ( .A(n_567), .Y(n_661) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI22x1_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_639), .B1(n_728), .B2(n_729), .Y(n_575) );
INVxp33_ASAP7_75t_SL g728 ( .A(n_576), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_578), .B1(n_607), .B2(n_608), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_582), .B(n_596), .Y(n_581) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_585), .Y(n_615) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g651 ( .A(n_595), .Y(n_651) );
INVx1_ASAP7_75t_L g853 ( .A(n_595), .Y(n_853) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_601), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B(n_600), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_598), .A2(n_702), .B(n_703), .C(n_705), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_623), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_630), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g823 ( .A(n_629), .Y(n_823) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_634), .B2(n_635), .C1(n_636), .C2(n_637), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g729 ( .A(n_639), .Y(n_729) );
OA22x2_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_662), .B1(n_663), .B2(n_727), .Y(n_639) );
INVx1_ASAP7_75t_L g727 ( .A(n_640), .Y(n_727) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND4xp75_ASAP7_75t_SL g643 ( .A(n_644), .B(n_647), .C(n_652), .D(n_656), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
BUFx2_ASAP7_75t_L g776 ( .A(n_657), .Y(n_776) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_661), .Y(n_782) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_685), .B1(n_725), .B2(n_726), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g726 ( .A(n_665), .Y(n_726) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_667), .B(n_676), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .C(n_672), .D(n_674), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .C(n_682), .D(n_683), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g966 ( .A(n_679), .Y(n_966) );
INVx4_ASAP7_75t_L g991 ( .A(n_679), .Y(n_991) );
INVx1_ASAP7_75t_L g779 ( .A(n_681), .Y(n_779) );
INVx2_ASAP7_75t_L g725 ( .A(n_685), .Y(n_725) );
OA22x2_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_711), .B2(n_724), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_710), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_700), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_695), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_697), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_706), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g724 ( .A(n_711), .Y(n_724) );
XNOR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_723), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_719), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .C(n_716), .D(n_718), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .C(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_733), .B1(n_834), .B2(n_947), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_795), .B1(n_796), .B2(n_833), .Y(n_733) );
INVx1_ASAP7_75t_SL g833 ( .A(n_734), .Y(n_833) );
XNOR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_772), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_756), .B1(n_770), .B2(n_771), .Y(n_735) );
INVx1_ASAP7_75t_L g770 ( .A(n_736), .Y(n_770) );
INVxp67_ASAP7_75t_L g857 ( .A(n_736), .Y(n_857) );
BUFx2_ASAP7_75t_L g858 ( .A(n_736), .Y(n_858) );
INVx2_ASAP7_75t_L g755 ( .A(n_738), .Y(n_755) );
NAND4xp75_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .C(n_748), .D(n_751), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
BUFx3_ASAP7_75t_L g787 ( .A(n_746), .Y(n_787) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_SL g771 ( .A(n_756), .Y(n_771) );
XOR2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_769), .Y(n_756) );
NAND4xp75_ASAP7_75t_L g757 ( .A(n_758), .B(n_762), .C(n_765), .D(n_768), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_SL g794 ( .A(n_773), .Y(n_794) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_785), .Y(n_773) );
NAND4xp25_ASAP7_75t_SL g774 ( .A(n_775), .B(n_777), .C(n_781), .D(n_783), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND4xp25_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .C(n_789), .D(n_792), .Y(n_785) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_813), .B1(n_831), .B2(n_832), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_798), .Y(n_831) );
INVx1_ASAP7_75t_L g812 ( .A(n_799), .Y(n_812) );
NOR2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_806), .Y(n_799) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .C(n_804), .D(n_805), .Y(n_800) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .C(n_809), .D(n_810), .Y(n_806) );
INVx4_ASAP7_75t_L g832 ( .A(n_813), .Y(n_832) );
INVx2_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_824), .Y(n_815) );
NAND4xp25_ASAP7_75t_SL g816 ( .A(n_817), .B(n_818), .C(n_819), .D(n_821), .Y(n_816) );
INVx1_ASAP7_75t_L g977 ( .A(n_820), .Y(n_977) );
INVx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .C(n_827), .D(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g947 ( .A(n_834), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B1(n_911), .B2(n_912), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
XNOR2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_859), .Y(n_836) );
OAI22xp5_ASAP7_75t_SL g837 ( .A1(n_838), .A2(n_839), .B1(n_857), .B2(n_858), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_848), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_846), .C(n_847), .Y(n_842) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND4xp25_ASAP7_75t_L g848 ( .A(n_849), .B(n_852), .C(n_854), .D(n_855), .Y(n_848) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_892), .B1(n_909), .B2(n_910), .Y(n_860) );
INVx2_ASAP7_75t_L g910 ( .A(n_861), .Y(n_910) );
AOI22x1_ASAP7_75t_SL g861 ( .A1(n_862), .A2(n_875), .B1(n_890), .B2(n_891), .Y(n_861) );
INVx1_ASAP7_75t_SL g891 ( .A(n_862), .Y(n_891) );
XNOR2x1_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
OR2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_870), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .C(n_869), .Y(n_865) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .C(n_873), .D(n_874), .Y(n_870) );
INVx3_ASAP7_75t_L g890 ( .A(n_875), .Y(n_890) );
AO22x2_ASAP7_75t_L g926 ( .A1(n_875), .A2(n_890), .B1(n_927), .B2(n_944), .Y(n_926) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR2x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_884), .Y(n_878) );
NAND4xp25_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .C(n_882), .D(n_883), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_888), .C(n_889), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
INVx2_ASAP7_75t_L g909 ( .A(n_892), .Y(n_909) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
XNOR2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
NAND2xp5_ASAP7_75t_SL g895 ( .A(n_896), .B(n_901), .Y(n_895) );
AND4x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .C(n_899), .D(n_900), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_907), .Y(n_901) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .C(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
OA22x2_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_926), .B1(n_945), .B2(n_946), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g945 ( .A(n_914), .Y(n_945) );
OR2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_921), .Y(n_915) );
NAND4xp25_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .C(n_919), .D(n_920), .Y(n_916) );
NAND4xp25_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .C(n_924), .D(n_925), .Y(n_921) );
INVx1_ASAP7_75t_L g946 ( .A(n_926), .Y(n_946) );
INVx1_ASAP7_75t_SL g944 ( .A(n_927), .Y(n_944) );
INVx1_ASAP7_75t_SL g943 ( .A(n_928), .Y(n_943) );
NOR2x1_ASAP7_75t_L g928 ( .A(n_929), .B(n_936), .Y(n_928) );
NAND4xp25_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .C(n_934), .D(n_935), .Y(n_929) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .C(n_939), .D(n_940), .Y(n_936) );
INVx1_ASAP7_75t_SL g949 ( .A(n_950), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_953), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_951), .B(n_954), .Y(n_1009) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
OAI222xp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_980), .B1(n_982), .B2(n_1007), .C1(n_1010), .C2(n_1013), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVxp33_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NOR3xp33_ASAP7_75t_SL g962 ( .A(n_963), .B(n_968), .C(n_975), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .Y(n_963) );
BUFx3_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
NAND4xp25_ASAP7_75t_SL g968 ( .A(n_969), .B(n_970), .C(n_972), .D(n_973), .Y(n_968) );
OAI21xp5_ASAP7_75t_SL g975 ( .A1(n_976), .A2(n_977), .B(n_978), .Y(n_975) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_998), .Y(n_983) );
NOR3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_988), .C(n_994), .Y(n_984) );
NAND2xp5_ASAP7_75t_SL g985 ( .A(n_986), .B(n_987), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_990), .B1(n_992), .B2(n_993), .Y(n_988) );
INVx2_ASAP7_75t_SL g990 ( .A(n_991), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1002), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1006), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_1008), .Y(n_1007) );
CKINVDCx6p67_ASAP7_75t_R g1008 ( .A(n_1009), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_1011), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_1012), .Y(n_1011) );
endmodule