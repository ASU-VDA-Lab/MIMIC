module real_jpeg_15024_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_59),
.B1(n_61),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_214)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_37),
.B1(n_64),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_59),
.B1(n_61),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_110),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_110),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_110),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_125),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_11),
.B(n_27),
.C(n_43),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_100),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_11),
.A2(n_24),
.B1(n_35),
.B2(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_106),
.Y(n_231)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_59),
.B1(n_61),
.B2(n_78),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_78),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_47),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_47),
.B1(n_64),
.B2(n_65),
.Y(n_120)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_20),
.B(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_91),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_21),
.B(n_81),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_22),
.B(n_54),
.C(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_23),
.B(n_38),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_24),
.A2(n_35),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_24),
.A2(n_35),
.B1(n_212),
.B2(n_220),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_24),
.A2(n_86),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_25),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_25),
.A2(n_34),
.B(n_87),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_29),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_26),
.B(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_35),
.A2(n_84),
.B(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_35),
.B(n_100),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B(n_48),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_39),
.A2(n_44),
.B1(n_51),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_39),
.A2(n_51),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_39),
.B(n_100),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_39),
.A2(n_51),
.B1(n_184),
.B2(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_40),
.B(n_49),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_40),
.A2(n_50),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_40),
.B(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA22x2_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_46),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_45),
.B(n_65),
.C(n_75),
.Y(n_180)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_46),
.A2(n_74),
.B(n_179),
.C(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_46),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_51),
.A2(n_90),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_51),
.A2(n_133),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_51),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_68),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_65),
.B(n_99),
.C(n_101),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_100),
.CON(n_99),
.SN(n_99)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.C(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_65),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_65),
.B(n_100),
.CON(n_179),
.SN(n_179)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_77),
.B(n_79),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_106),
.B1(n_156),
.B2(n_179),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_103),
.B1(n_104),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_76),
.A2(n_104),
.B1(n_146),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_91),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.C(n_107),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_92),
.A2(n_93),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_109),
.B1(n_125),
.B2(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_102),
.B(n_107),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_135),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_127),
.B2(n_128),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_249),
.C(n_253),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_160),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_160),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.C(n_153),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_144),
.C(n_149),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_250)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_243),
.B(n_248),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_198),
.B(n_242),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_186),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_181),
.C(n_182),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_173),
.A2(n_174),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_182),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_187),
.B(n_192),
.C(n_196),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_196),
.B2(n_197),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_236),
.B(n_241),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_226),
.B(n_235),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_215),
.B(n_225),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_221),
.B(n_224),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);


endmodule