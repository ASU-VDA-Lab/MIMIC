module fake_netlist_6_3604_n_1808 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1808);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1808;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_21),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_86),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_41),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_45),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_112),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_63),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_47),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_92),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_23),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_38),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_54),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_42),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_83),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_54),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_116),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_32),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_89),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_48),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_19),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_24),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_55),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_23),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_121),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_117),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_163),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_22),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_20),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_145),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_147),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_48),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_18),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_131),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_20),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_104),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_35),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_118),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_13),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_125),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_107),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_166),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_93),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_62),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_128),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_140),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_111),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_40),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_87),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_101),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_149),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_4),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_129),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_2),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_106),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_22),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_57),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_33),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_154),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_97),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_60),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_65),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_141),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_146),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_94),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_67),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_35),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_70),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_158),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_58),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_96),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_151),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_148),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_31),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_49),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_167),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_134),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_136),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_34),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_75),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_79),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_108),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_44),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_36),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_39),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_74),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_139),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_95),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_102),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_29),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_0),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_62),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_50),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_53),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_17),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

BUFx8_ASAP7_75t_SL g326 ( 
.A(n_91),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_113),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_61),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_28),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_47),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_30),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_52),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_14),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_85),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_50),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_66),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_169),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_169),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_169),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_326),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_217),
.B(n_1),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_172),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_170),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_192),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_178),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_184),
.B(n_1),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_169),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_184),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_185),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_175),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_248),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_186),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_180),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_169),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_190),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_249),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_176),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_177),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_173),
.B(n_4),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_187),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_191),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_301),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_194),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_246),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_228),
.B(n_5),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_199),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_204),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_171),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_171),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_206),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_196),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_228),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_196),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_227),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_213),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_263),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_219),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_263),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_227),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_262),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_183),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_221),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_240),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_240),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_190),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_224),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_246),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_211),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_225),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_229),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_230),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_275),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_237),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_275),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_276),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_220),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_276),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_239),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_241),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_220),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_247),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_251),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_252),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_262),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_254),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_340),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_352),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_349),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_370),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_267),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_368),
.B(n_258),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_368),
.B(n_259),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_195),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_267),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_342),
.B(n_189),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_362),
.B(n_243),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_348),
.B(n_321),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_367),
.B(n_261),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_353),
.B(n_360),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_267),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_375),
.A2(n_321),
.B(n_205),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_341),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_361),
.B(n_226),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_381),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_350),
.B(n_265),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_235),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_382),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_350),
.B(n_273),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_338),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_358),
.B(n_211),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_358),
.B(n_211),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_348),
.B(n_195),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_395),
.A2(n_205),
.B(n_203),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_278),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_488),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_403),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_446),
.A2(n_447),
.B1(n_488),
.B2(n_472),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_460),
.Y(n_498)
);

NOR2x1p5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_215),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_344),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_442),
.B(n_262),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_460),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_423),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_460),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_407),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_436),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_446),
.A2(n_371),
.B1(n_380),
.B2(n_374),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_467),
.B(n_359),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_R g517 ( 
.A(n_436),
.B(n_347),
.Y(n_517)
);

NAND2x1p5_ASAP7_75t_L g518 ( 
.A(n_460),
.B(n_173),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_438),
.B(n_405),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_447),
.B(n_472),
.C(n_467),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_480),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_483),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_351),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_476),
.B(n_359),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_489),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_489),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_426),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_355),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_426),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_363),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_438),
.B(n_405),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_428),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_458),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_461),
.B(n_369),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_471),
.B(n_407),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_431),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_488),
.B(n_449),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_431),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_428),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_471),
.B(n_364),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_419),
.A2(n_179),
.B(n_174),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_458),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_452),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_482),
.B(n_366),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_476),
.A2(n_416),
.B1(n_383),
.B2(n_388),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_452),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_419),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_369),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_482),
.B(n_386),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_432),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_432),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

BUFx6f_ASAP7_75t_SL g579 ( 
.A(n_442),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_424),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_443),
.B(n_280),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_424),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_458),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_445),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_424),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_492),
.A2(n_412),
.B1(n_332),
.B2(n_198),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_454),
.B(n_397),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_427),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_428),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_427),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_449),
.B(n_401),
.C(n_400),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_461),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_429),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_486),
.A2(n_279),
.B1(n_215),
.B2(n_209),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_492),
.A2(n_409),
.B1(n_404),
.B2(n_393),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_432),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_432),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_445),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_443),
.B(n_280),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_455),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_434),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_486),
.A2(n_279),
.B1(n_215),
.B2(n_209),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_434),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_455),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_486),
.A2(n_414),
.B1(n_410),
.B2(n_402),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_487),
.B(n_415),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_433),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_442),
.B(n_262),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_442),
.B(n_262),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_453),
.B(n_315),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_433),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_434),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_487),
.B(n_412),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_434),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_453),
.B(n_282),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_434),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_433),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_434),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_442),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_455),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_487),
.B(n_284),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_434),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_442),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_456),
.B(n_289),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_485),
.B(n_174),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_485),
.Y(n_632)
);

AND3x1_ASAP7_75t_L g633 ( 
.A(n_483),
.B(n_218),
.C(n_203),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_435),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_434),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_456),
.A2(n_245),
.B1(n_270),
.B2(n_269),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_461),
.B(n_396),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_469),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_456),
.B(n_253),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_435),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_456),
.B(n_382),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_440),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_628),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_497),
.A2(n_365),
.B1(n_354),
.B2(n_345),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_520),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_523),
.B(n_207),
.C(n_188),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_545),
.B(n_343),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_564),
.B(n_290),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_582),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_499),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_568),
.B(n_202),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_493),
.A2(n_309),
.B1(n_304),
.B2(n_287),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_493),
.B(n_440),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_585),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_504),
.A2(n_292),
.B1(n_302),
.B2(n_288),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_504),
.B(n_262),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_632),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_632),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_561),
.B(n_440),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_618),
.B(n_212),
.C(n_210),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_565),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_567),
.B(n_440),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_585),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_214),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_509),
.B(n_279),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_525),
.B(n_231),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_526),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_554),
.A2(n_238),
.B1(n_325),
.B2(n_302),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_515),
.B(n_233),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_574),
.B(n_293),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_554),
.B(n_440),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_529),
.B(n_440),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_598),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_524),
.A2(n_313),
.B(n_292),
.C(n_325),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_615),
.B(n_440),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_609),
.B(n_295),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_501),
.B(n_440),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_565),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_536),
.B(n_444),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_549),
.B(n_611),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_524),
.A2(n_527),
.B1(n_534),
.B2(n_533),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_496),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_L g686 ( 
.A1(n_549),
.A2(n_307),
.B1(n_317),
.B2(n_300),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_511),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_496),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_522),
.A2(n_318),
.B1(n_298),
.B2(n_306),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_583),
.B(n_236),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_522),
.A2(n_327),
.B1(n_310),
.B2(n_311),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_514),
.B(n_389),
.C(n_387),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_626),
.B(n_242),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_538),
.B(n_444),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_610),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_593),
.B(n_316),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_511),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_539),
.A2(n_334),
.B1(n_179),
.B2(n_296),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_526),
.B(n_253),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_637),
.B(n_218),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_516),
.B(n_264),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_597),
.B(n_389),
.C(n_387),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_539),
.B(n_253),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_588),
.B(n_266),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_638),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_620),
.B(n_444),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_527),
.A2(n_260),
.B(n_257),
.C(n_313),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_509),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_616),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_530),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_586),
.B(n_253),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_581),
.A2(n_317),
.B1(n_222),
.B2(n_307),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_533),
.B(n_444),
.Y(n_715)
);

BUFx12f_ASAP7_75t_SL g716 ( 
.A(n_637),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_534),
.B(n_444),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_550),
.B(n_444),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_550),
.B(n_444),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_628),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_638),
.B(n_268),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_641),
.B(n_285),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_622),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_540),
.B(n_271),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_581),
.A2(n_193),
.B1(n_222),
.B2(n_197),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_562),
.A2(n_505),
.B1(n_500),
.B2(n_498),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_542),
.B(n_272),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_631),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_581),
.A2(n_182),
.B1(n_197),
.B2(n_193),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_622),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_548),
.B(n_558),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_596),
.B(n_285),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_569),
.B(n_274),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_570),
.B(n_277),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_634),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_634),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_591),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_562),
.B(n_444),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_505),
.B(n_450),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_640),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_572),
.B(n_450),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_507),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_602),
.B(n_223),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_631),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_580),
.B(n_450),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_587),
.B(n_450),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_606),
.B(n_285),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_589),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_R g750 ( 
.A(n_517),
.B(n_283),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_513),
.A2(n_255),
.B1(n_232),
.B2(n_238),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_592),
.A2(n_309),
.B(n_304),
.C(n_182),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_602),
.B(n_223),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_631),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_544),
.Y(n_755)
);

OAI21xp33_ASAP7_75t_L g756 ( 
.A1(n_636),
.A2(n_255),
.B(n_232),
.Y(n_756)
);

AND2x6_ASAP7_75t_SL g757 ( 
.A(n_637),
.B(n_234),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_537),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_518),
.A2(n_256),
.B(n_234),
.C(n_250),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_510),
.B(n_220),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_544),
.B(n_285),
.Y(n_761)
);

OAI221xp5_ASAP7_75t_L g762 ( 
.A1(n_633),
.A2(n_256),
.B1(n_250),
.B2(n_257),
.C(n_260),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_595),
.B(n_450),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_612),
.B(n_294),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_518),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_629),
.B(n_478),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_494),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_560),
.B(n_223),
.Y(n_769)
);

O2A1O1Ixp5_ASAP7_75t_L g770 ( 
.A1(n_563),
.A2(n_451),
.B(n_457),
.C(n_435),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_518),
.A2(n_330),
.B1(n_288),
.B2(n_281),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_639),
.A2(n_200),
.B1(n_287),
.B2(n_296),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_581),
.A2(n_603),
.B1(n_571),
.B2(n_546),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_519),
.B(n_478),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_637),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_519),
.B(n_532),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_519),
.B(n_478),
.Y(n_778)
);

OAI21xp33_ASAP7_75t_L g779 ( 
.A1(n_546),
.A2(n_330),
.B(n_299),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_546),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_494),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_495),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_581),
.A2(n_200),
.B1(n_281),
.B2(n_286),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_546),
.B(n_305),
.Y(n_784)
);

AO22x2_ASAP7_75t_L g785 ( 
.A1(n_532),
.A2(n_300),
.B1(n_291),
.B2(n_286),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_571),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_608),
.Y(n_787)
);

OAI21xp33_ASAP7_75t_L g788 ( 
.A1(n_571),
.A2(n_322),
.B(n_329),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_SL g789 ( 
.A1(n_594),
.A2(n_328),
.B1(n_324),
.B2(n_323),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_625),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_508),
.B(n_291),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_535),
.B(n_478),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_625),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_502),
.A2(n_479),
.B(n_474),
.C(n_469),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_581),
.A2(n_442),
.B1(n_469),
.B2(n_474),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_603),
.A2(n_442),
.B1(n_474),
.B2(n_479),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_630),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_537),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_630),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_571),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_602),
.B(n_223),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_535),
.B(n_308),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_537),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_502),
.B(n_335),
.C(n_312),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_556),
.B(n_484),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_556),
.B(n_484),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_556),
.B(n_484),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_624),
.B(n_223),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_495),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_573),
.B(n_578),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_675),
.A2(n_512),
.B(n_503),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_687),
.Y(n_812)
);

OAI321xp33_ASAP7_75t_L g813 ( 
.A1(n_713),
.A2(n_563),
.A3(n_413),
.B1(n_406),
.B2(n_408),
.C(n_411),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_643),
.B(n_624),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_661),
.A2(n_512),
.B(n_503),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_664),
.A2(n_512),
.B(n_503),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_649),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_670),
.A2(n_573),
.B1(n_578),
.B2(n_607),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_653),
.A2(n_642),
.B(n_635),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_697),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_670),
.A2(n_603),
.B1(n_613),
.B2(n_614),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_673),
.A2(n_600),
.B(n_573),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_683),
.B(n_578),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_643),
.B(n_603),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_715),
.A2(n_642),
.B(n_635),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_717),
.A2(n_719),
.B(n_718),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_693),
.B(n_731),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_677),
.A2(n_613),
.B(n_614),
.C(n_577),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

AOI33xp33_ASAP7_75t_L g830 ( 
.A1(n_657),
.A2(n_406),
.A3(n_413),
.B1(n_411),
.B2(n_408),
.B3(n_479),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_693),
.B(n_603),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_683),
.B(n_669),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_750),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_738),
.A2(n_739),
.B(n_726),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_680),
.A2(n_642),
.B(n_635),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_643),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_731),
.B(n_600),
.Y(n_837)
);

BUFx4f_ASAP7_75t_L g838 ( 
.A(n_701),
.Y(n_838)
);

BUFx4f_ASAP7_75t_L g839 ( 
.A(n_701),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_682),
.A2(n_531),
.B(n_541),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_SL g841 ( 
.A(n_651),
.B(n_594),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_649),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_720),
.B(n_624),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_659),
.B(n_600),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_660),
.B(n_607),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_671),
.B(n_607),
.Y(n_846)
);

AOI33xp33_ASAP7_75t_L g847 ( 
.A1(n_657),
.A2(n_220),
.A3(n_303),
.B1(n_475),
.B2(n_470),
.B3(n_331),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_750),
.A2(n_303),
.B1(n_244),
.B2(n_336),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_663),
.B(n_623),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_694),
.A2(n_543),
.B(n_575),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_681),
.B(n_623),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_751),
.A2(n_579),
.B1(n_262),
.B2(n_244),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_743),
.B(n_623),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_244),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_720),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_745),
.A2(n_579),
.B1(n_576),
.B2(n_619),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_654),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_707),
.A2(n_531),
.B(n_575),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_678),
.A2(n_531),
.B(n_575),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_743),
.B(n_537),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_654),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_737),
.Y(n_862)
);

BUFx2_ASAP7_75t_SL g863 ( 
.A(n_755),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_744),
.A2(n_521),
.B(n_506),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_768),
.B(n_508),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_726),
.A2(n_552),
.B(n_506),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_655),
.Y(n_867)
);

O2A1O1Ixp5_ASAP7_75t_L g868 ( 
.A1(n_744),
.A2(n_576),
.B(n_543),
.C(n_619),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_751),
.A2(n_484),
.B(n_314),
.C(n_320),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_766),
.A2(n_576),
.B(n_543),
.Y(n_870)
);

AND2x4_ASAP7_75t_SL g871 ( 
.A(n_720),
.B(n_303),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_720),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_655),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_645),
.B(n_541),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_658),
.A2(n_684),
.B(n_777),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_684),
.A2(n_521),
.B(n_528),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_665),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_656),
.B(n_541),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_765),
.A2(n_619),
.B1(n_579),
.B2(n_627),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_745),
.B(n_537),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_810),
.A2(n_627),
.B(n_621),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_754),
.B(n_599),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_665),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_671),
.B(n_599),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_754),
.B(n_599),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_SL g886 ( 
.A1(n_686),
.A2(n_551),
.B(n_590),
.C(n_584),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_685),
.B(n_599),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_753),
.A2(n_627),
.B(n_621),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_674),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_771),
.B(n_599),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_771),
.B(n_605),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_666),
.B(n_303),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_770),
.A2(n_551),
.B(n_528),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_753),
.A2(n_778),
.B(n_775),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_676),
.Y(n_895)
);

O2A1O1Ixp5_ASAP7_75t_L g896 ( 
.A1(n_722),
.A2(n_555),
.B(n_552),
.C(n_553),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_801),
.A2(n_557),
.B(n_553),
.C(n_555),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_808),
.A2(n_547),
.B(n_559),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_774),
.B(n_627),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_666),
.B(n_605),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_647),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_695),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_792),
.A2(n_557),
.B(n_547),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_SL g904 ( 
.A1(n_752),
.A2(n_601),
.B(n_590),
.C(n_584),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_695),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_668),
.B(n_605),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_668),
.B(n_605),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_688),
.B(n_605),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_700),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_710),
.B(n_617),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_690),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_758),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_708),
.A2(n_601),
.B(n_577),
.C(n_559),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_700),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_805),
.A2(n_621),
.B(n_617),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_760),
.B(n_333),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_711),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_806),
.A2(n_617),
.B(n_566),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_807),
.A2(n_617),
.B(n_566),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_741),
.A2(n_566),
.B(n_508),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_711),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_746),
.A2(n_566),
.B(n_508),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_747),
.A2(n_566),
.B(n_508),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_730),
.B(n_448),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_735),
.B(n_448),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_758),
.Y(n_926)
);

AOI21xp33_ASAP7_75t_L g927 ( 
.A1(n_705),
.A2(n_244),
.B(n_336),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_763),
.A2(n_803),
.B(n_798),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_709),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_667),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_721),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_798),
.A2(n_421),
.B(n_464),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_705),
.A2(n_448),
.B(n_462),
.Y(n_933)
);

AND2x6_ASAP7_75t_L g934 ( 
.A(n_795),
.B(n_244),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_462),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_803),
.A2(n_421),
.B(n_459),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_723),
.B(n_336),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_723),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_712),
.B(n_5),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_728),
.A2(n_421),
.B(n_459),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_736),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_736),
.Y(n_942)
);

O2A1O1Ixp5_ASAP7_75t_L g943 ( 
.A1(n_672),
.A2(n_462),
.B(n_451),
.C(n_457),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_690),
.B(n_470),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_701),
.B(n_336),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_742),
.A2(n_421),
.B(n_464),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_749),
.B(n_451),
.Y(n_947)
);

AOI21xp33_ASAP7_75t_L g948 ( 
.A1(n_702),
.A2(n_336),
.B(n_7),
.Y(n_948)
);

BUFx12f_ASAP7_75t_L g949 ( 
.A(n_757),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_773),
.A2(n_464),
.B(n_459),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_786),
.A2(n_451),
.B1(n_457),
.B2(n_470),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_780),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_650),
.A2(n_421),
.B(n_464),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_644),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_802),
.A2(n_421),
.B(n_459),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_662),
.B(n_64),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_692),
.B(n_470),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_734),
.B(n_451),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_767),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_721),
.Y(n_960)
);

NOR2x1p5_ASAP7_75t_L g961 ( 
.A(n_646),
.B(n_475),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_702),
.B(n_475),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_734),
.B(n_457),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_699),
.B(n_6),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_764),
.B(n_457),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_776),
.B(n_475),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_796),
.B(n_421),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_802),
.A2(n_491),
.B(n_490),
.C(n_481),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_764),
.B(n_491),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_767),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_696),
.A2(n_491),
.B(n_490),
.C(n_481),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_724),
.B(n_491),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_756),
.A2(n_762),
.B(n_779),
.C(n_759),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_648),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_716),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_724),
.B(n_491),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_L g977 ( 
.A(n_804),
.B(n_491),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_781),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_787),
.A2(n_463),
.B(n_490),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_784),
.A2(n_491),
.B(n_490),
.C(n_481),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_781),
.A2(n_463),
.B(n_490),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_800),
.B(n_491),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_703),
.B(n_490),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_761),
.B(n_6),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_727),
.B(n_490),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_652),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_782),
.A2(n_463),
.B(n_481),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_790),
.A2(n_799),
.B(n_797),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_772),
.B(n_714),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_793),
.A2(n_463),
.B(n_481),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_725),
.A2(n_490),
.B1(n_481),
.B2(n_477),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_782),
.A2(n_463),
.B(n_477),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_809),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_789),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_791),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_929),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_827),
.A2(n_729),
.B1(n_783),
.B2(n_689),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_929),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_911),
.B(n_704),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_911),
.A2(n_784),
.B(n_733),
.C(n_727),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_948),
.A2(n_769),
.B(n_679),
.C(n_748),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_862),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_820),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_873),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_986),
.A2(n_785),
.B1(n_732),
.B2(n_698),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_832),
.A2(n_788),
.B(n_733),
.C(n_794),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_832),
.B(n_691),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_984),
.A2(n_791),
.B(n_785),
.C(n_11),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_931),
.B(n_785),
.C(n_9),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_916),
.B(n_481),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_812),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_833),
.B(n_162),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_944),
.B(n_481),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_986),
.A2(n_477),
.B1(n_473),
.B2(n_468),
.Y(n_1015)
);

OR2x4_ASAP7_75t_L g1016 ( 
.A(n_984),
.B(n_477),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_817),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_889),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_964),
.A2(n_973),
.B(n_846),
.C(n_821),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_823),
.B(n_477),
.Y(n_1020)
);

CKINVDCx8_ASAP7_75t_R g1021 ( 
.A(n_863),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_889),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_824),
.A2(n_463),
.B(n_473),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_952),
.B(n_133),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_823),
.B(n_477),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_892),
.B(n_477),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_964),
.A2(n_973),
.B(n_960),
.C(n_939),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_950),
.A2(n_127),
.B(n_71),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_812),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_927),
.A2(n_8),
.B(n_9),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_884),
.B(n_477),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_846),
.A2(n_473),
.B(n_468),
.C(n_466),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_831),
.A2(n_473),
.B(n_468),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_954),
.A2(n_473),
.B1(n_468),
.B2(n_466),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_975),
.B(n_473),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_842),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_829),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_930),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_829),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_867),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_960),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_821),
.B(n_473),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_952),
.B(n_115),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_829),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_901),
.B(n_468),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_829),
.B(n_468),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_466),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_939),
.B(n_8),
.C(n_11),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_836),
.B(n_466),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_814),
.A2(n_465),
.B(n_466),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_930),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_877),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_843),
.A2(n_465),
.B(n_466),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_962),
.B(n_466),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_L g1055 ( 
.A(n_852),
.B(n_465),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_957),
.A2(n_465),
.B(n_16),
.C(n_17),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_900),
.B(n_906),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_877),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_875),
.A2(n_465),
.B(n_16),
.C(n_19),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_907),
.B(n_465),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_871),
.B(n_974),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_837),
.B(n_465),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_883),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_983),
.A2(n_465),
.B1(n_161),
.B2(n_157),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_871),
.B(n_13),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_843),
.A2(n_153),
.B(n_150),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_883),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_989),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_836),
.B(n_142),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_890),
.A2(n_110),
.B1(n_100),
.B2(n_99),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_826),
.A2(n_84),
.B(n_80),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_905),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_855),
.B(n_68),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_841),
.A2(n_76),
.B1(n_26),
.B2(n_30),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_855),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_917),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_811),
.A2(n_816),
.B(n_815),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_895),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_917),
.B(n_25),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_872),
.B(n_32),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_834),
.A2(n_34),
.B(n_36),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_994),
.B(n_37),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_872),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_SL g1084 ( 
.A1(n_949),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_941),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_989),
.A2(n_44),
.B(n_45),
.C(n_49),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_887),
.B(n_51),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_908),
.B(n_52),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_869),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_941),
.B(n_874),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_852),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_891),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_978),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_835),
.A2(n_63),
.B(n_840),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_887),
.B(n_909),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_914),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_921),
.B(n_938),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_942),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_961),
.A2(n_966),
.B1(n_874),
.B2(n_878),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_978),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_869),
.A2(n_828),
.B(n_847),
.C(n_963),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_857),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_899),
.A2(n_972),
.B(n_985),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_966),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_861),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_878),
.B(n_902),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_848),
.A2(n_956),
.B1(n_899),
.B2(n_839),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_958),
.B(n_965),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_976),
.B(n_969),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_912),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_982),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_838),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_SL g1113 ( 
.A1(n_980),
.A2(n_851),
.B(n_849),
.C(n_937),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_854),
.B(n_844),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_860),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_850),
.A2(n_858),
.B(n_870),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_830),
.A2(n_847),
.B(n_822),
.C(n_813),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_819),
.A2(n_825),
.B(n_859),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_982),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_980),
.A2(n_894),
.B(n_893),
.Y(n_1120)
);

AO22x1_ASAP7_75t_L g1121 ( 
.A1(n_934),
.A2(n_995),
.B1(n_993),
.B2(n_970),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_982),
.B(n_945),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_854),
.B(n_838),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_934),
.A2(n_959),
.B1(n_933),
.B2(n_935),
.Y(n_1124)
);

OR2x6_ASAP7_75t_SL g1125 ( 
.A(n_839),
.B(n_845),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_943),
.A2(n_988),
.B(n_968),
.C(n_947),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_854),
.B(n_945),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_924),
.B(n_925),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_945),
.A2(n_880),
.B1(n_882),
.B2(n_885),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_853),
.Y(n_1130)
);

NAND3xp33_ASAP7_75t_SL g1131 ( 
.A(n_830),
.B(n_953),
.C(n_856),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_910),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_879),
.A2(n_881),
.B(n_876),
.Y(n_1133)
);

INVx6_ASAP7_75t_L g1134 ( 
.A(n_912),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_912),
.B(n_937),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_913),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_934),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_995),
.B(n_926),
.Y(n_1138)
);

OAI22x1_ASAP7_75t_L g1139 ( 
.A1(n_926),
.A2(n_967),
.B1(n_864),
.B2(n_934),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_896),
.A2(n_971),
.B(n_868),
.C(n_928),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_934),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_990),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_951),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_898),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_866),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_886),
.A2(n_904),
.B(n_818),
.C(n_967),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_886),
.A2(n_904),
.B1(n_940),
.B2(n_903),
.C(n_946),
.Y(n_1147)
);

AOI221x1_ASAP7_75t_L g1148 ( 
.A1(n_1081),
.A2(n_955),
.B1(n_915),
.B2(n_888),
.C(n_991),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1057),
.A2(n_977),
.B(n_865),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1048),
.A2(n_981),
.B1(n_987),
.B2(n_979),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1036),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_L g1152 ( 
.A(n_1019),
.B(n_919),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1109),
.A2(n_918),
.B(n_897),
.Y(n_1153)
);

INVx5_ASAP7_75t_L g1154 ( 
.A(n_1035),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1033),
.A2(n_992),
.B(n_936),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1008),
.B(n_932),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1109),
.A2(n_920),
.B(n_922),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1128),
.B(n_923),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1112),
.B(n_1104),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1051),
.B(n_1024),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1017),
.Y(n_1161)
);

OAI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1041),
.A2(n_1082),
.B1(n_1074),
.B2(n_1016),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1050),
.A2(n_1053),
.B(n_1133),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1146),
.A2(n_1028),
.B(n_1094),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1023),
.A2(n_1042),
.B(n_1142),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_996),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_999),
.B(n_1000),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_1002),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1108),
.A2(n_1047),
.B(n_1031),
.Y(n_1169)
);

AO22x2_ASAP7_75t_L g1170 ( 
.A1(n_1048),
.A2(n_1010),
.B1(n_1092),
.B2(n_997),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1059),
.A2(n_1068),
.B1(n_1089),
.B2(n_1056),
.C(n_1071),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1032),
.A2(n_1103),
.B(n_1140),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1101),
.A2(n_1126),
.A3(n_1117),
.B(n_1139),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1027),
.A2(n_1007),
.B(n_1001),
.C(n_999),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1132),
.B(n_1145),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1108),
.A2(n_1055),
.B(n_1026),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1117),
.A2(n_1025),
.A3(n_1020),
.B(n_1030),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1040),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1082),
.A2(n_1086),
.B(n_1079),
.C(n_1009),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_1054),
.B(n_1014),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_SL g1181 ( 
.A(n_1021),
.B(n_1075),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1147),
.A2(n_1060),
.B(n_1062),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1046),
.A2(n_1049),
.B(n_1138),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1091),
.A2(n_1016),
.B1(n_1005),
.B2(n_1124),
.Y(n_1184)
);

CKINVDCx8_ASAP7_75t_R g1185 ( 
.A(n_1038),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1125),
.B2(n_998),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1046),
.A2(n_1049),
.B(n_1138),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1018),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1110),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1136),
.A2(n_1088),
.A3(n_1097),
.B(n_1143),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1115),
.B(n_1130),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1075),
.B(n_1037),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_996),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1088),
.A2(n_1097),
.A3(n_1114),
.B(n_1070),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_1029),
.B(n_1012),
.C(n_998),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1113),
.A2(n_1115),
.B(n_1120),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1012),
.A2(n_1029),
.B(n_1087),
.C(n_1114),
.Y(n_1197)
);

NOR2x1_ASAP7_75t_SL g1198 ( 
.A(n_1035),
.B(n_1090),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1113),
.A2(n_1120),
.B(n_1011),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1024),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1005),
.A2(n_1064),
.B(n_1095),
.C(n_1129),
.Y(n_1202)
);

AO32x2_ASAP7_75t_L g1203 ( 
.A1(n_1141),
.A2(n_1084),
.A3(n_1039),
.B1(n_1037),
.B2(n_1091),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1090),
.A2(n_1106),
.B(n_1121),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1123),
.B(n_1095),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1122),
.B(n_1035),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1043),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1066),
.A2(n_1124),
.B(n_1022),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1122),
.A2(n_1141),
.B1(n_1015),
.B2(n_1078),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1106),
.A2(n_1131),
.B(n_1144),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1045),
.B(n_1063),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1144),
.A2(n_1015),
.B(n_1073),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1034),
.A2(n_1102),
.B(n_1105),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1043),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1110),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1080),
.A2(n_1098),
.B(n_1096),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1063),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1013),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1135),
.A2(n_1072),
.B(n_1100),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1134),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1072),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1127),
.B(n_1004),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1093),
.A2(n_1067),
.B(n_1076),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1039),
.B(n_1073),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1111),
.B(n_1119),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1052),
.A2(n_1058),
.B(n_1085),
.C(n_1119),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1069),
.A2(n_1111),
.B(n_1137),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1044),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1083),
.A2(n_1144),
.B(n_1110),
.C(n_1013),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1110),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_SL g1231 ( 
.A(n_1134),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1134),
.B(n_827),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1019),
.A2(n_1101),
.B(n_1027),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1003),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1019),
.A2(n_1000),
.B(n_827),
.C(n_1027),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1082),
.B(n_1048),
.C(n_644),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1036),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1000),
.A2(n_497),
.B(n_827),
.C(n_1027),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1061),
.B(n_931),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1019),
.A2(n_1000),
.B(n_827),
.C(n_1027),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1027),
.A2(n_523),
.B1(n_497),
.B2(n_446),
.C(n_515),
.Y(n_1241)
);

AO21x1_ASAP7_75t_L g1242 ( 
.A1(n_1027),
.A2(n_1081),
.B(n_1007),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1036),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1019),
.B(n_827),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1103),
.A2(n_1140),
.A3(n_1032),
.B(n_1133),
.Y(n_1245)
);

OAI22x1_ASAP7_75t_L g1246 ( 
.A1(n_1082),
.A2(n_960),
.B1(n_1107),
.B2(n_984),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1112),
.B(n_952),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1008),
.A2(n_651),
.B1(n_841),
.B2(n_931),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1041),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1081),
.A2(n_446),
.B(n_447),
.C(n_705),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1008),
.B(n_827),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1000),
.A2(n_497),
.B(n_827),
.C(n_1027),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1036),
.Y(n_1254)
);

BUFx2_ASAP7_75t_R g1255 ( 
.A(n_1021),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1048),
.A2(n_523),
.B1(n_497),
.B2(n_827),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1019),
.B(n_841),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1118),
.A2(n_1116),
.B(n_1077),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1002),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1008),
.B(n_827),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1008),
.B(n_827),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1036),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1035),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_996),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1027),
.A2(n_497),
.B1(n_1081),
.B2(n_1019),
.C(n_670),
.Y(n_1266)
);

NAND2xp33_ASAP7_75t_R g1267 ( 
.A(n_1013),
.B(n_750),
.Y(n_1267)
);

AO32x2_ASAP7_75t_L g1268 ( 
.A1(n_1092),
.A2(n_497),
.A3(n_652),
.B1(n_997),
.B2(n_1070),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1118),
.A2(n_1116),
.B(n_1077),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1109),
.A2(n_1108),
.B(n_1133),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1061),
.B(n_931),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1019),
.A2(n_1000),
.B(n_827),
.C(n_1027),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1008),
.B(n_827),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1061),
.B(n_931),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1118),
.A2(n_1116),
.B(n_1077),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1019),
.A2(n_1101),
.B(n_1027),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1103),
.A2(n_1140),
.A3(n_1032),
.B(n_1133),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1019),
.A2(n_670),
.B1(n_827),
.B2(n_1091),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1110),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1103),
.A2(n_1140),
.A3(n_1032),
.B(n_1133),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1036),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1000),
.A2(n_497),
.B(n_827),
.C(n_1027),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1133),
.A2(n_1032),
.B(n_968),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1008),
.B(n_931),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1036),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1118),
.A2(n_1116),
.B(n_1077),
.Y(n_1290)
);

BUFx2_ASAP7_75t_R g1291 ( 
.A(n_1021),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1057),
.A2(n_1109),
.B(n_831),
.Y(n_1292)
);

AO21x1_ASAP7_75t_L g1293 ( 
.A1(n_1027),
.A2(n_1081),
.B(n_1007),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1006),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1241),
.A2(n_1280),
.B1(n_1257),
.B2(n_1256),
.Y(n_1295)
);

AND2x4_ASAP7_75t_SL g1296 ( 
.A(n_1160),
.B(n_1247),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1234),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1151),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1257),
.A2(n_1280),
.B1(n_1256),
.B2(n_1184),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1168),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1199),
.B(n_1239),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1236),
.A2(n_1248),
.B1(n_1267),
.B2(n_1205),
.Y(n_1302)
);

CKINVDCx11_ASAP7_75t_R g1303 ( 
.A(n_1259),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1250),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1185),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1247),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1184),
.A2(n_1260),
.B1(n_1261),
.B2(n_1274),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1218),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1231),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1154),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1242),
.A2(n_1293),
.B1(n_1170),
.B2(n_1246),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1237),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1220),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1271),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1170),
.A2(n_1167),
.B1(n_1233),
.B2(n_1277),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1252),
.A2(n_1244),
.B1(n_1287),
.B2(n_1233),
.Y(n_1317)
);

BUFx8_ASAP7_75t_SL g1318 ( 
.A(n_1275),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1201),
.A2(n_1240),
.B1(n_1272),
.B2(n_1235),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1244),
.A2(n_1214),
.B1(n_1207),
.B2(n_1174),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1166),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1255),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1277),
.A2(n_1162),
.B1(n_1186),
.B2(n_1156),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1198),
.A2(n_1154),
.B1(n_1263),
.B2(n_1212),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1291),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1152),
.A2(n_1175),
.B1(n_1289),
.B2(n_1283),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1266),
.A2(n_1160),
.B1(n_1222),
.B2(n_1181),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1265),
.A2(n_1159),
.B1(n_1206),
.B2(n_1193),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1154),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1243),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1254),
.A2(n_1262),
.B1(n_1191),
.B2(n_1265),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1159),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1263),
.A2(n_1227),
.B1(n_1209),
.B2(n_1266),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1230),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1232),
.A2(n_1294),
.B1(n_1161),
.B2(n_1188),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1217),
.A2(n_1221),
.B1(n_1216),
.B2(n_1158),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1228),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1171),
.A2(n_1206),
.B1(n_1263),
.B2(n_1211),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1225),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1206),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1238),
.A2(n_1284),
.B(n_1253),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1202),
.A2(n_1209),
.B1(n_1224),
.B2(n_1229),
.Y(n_1342)
);

CKINVDCx6p67_ASAP7_75t_R g1343 ( 
.A(n_1189),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1158),
.A2(n_1251),
.B1(n_1213),
.B2(n_1210),
.Y(n_1344)
);

BUFx8_ASAP7_75t_L g1345 ( 
.A(n_1189),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1197),
.B(n_1195),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1223),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1213),
.A2(n_1227),
.B1(n_1288),
.B2(n_1286),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1219),
.A2(n_1196),
.B1(n_1204),
.B2(n_1200),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1203),
.A2(n_1179),
.B1(n_1150),
.B2(n_1219),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1215),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1249),
.A2(n_1292),
.B1(n_1273),
.B2(n_1278),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1264),
.A2(n_1150),
.B1(n_1180),
.B2(n_1172),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1172),
.A2(n_1169),
.B1(n_1176),
.B2(n_1268),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1223),
.Y(n_1355)
);

BUFx10_ASAP7_75t_L g1356 ( 
.A(n_1192),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1226),
.A2(n_1281),
.B1(n_1208),
.B2(n_1149),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1203),
.A2(n_1148),
.B1(n_1268),
.B2(n_1270),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1203),
.A2(n_1268),
.B1(n_1285),
.B2(n_1164),
.Y(n_1359)
);

INVx8_ASAP7_75t_L g1360 ( 
.A(n_1183),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1182),
.A2(n_1285),
.B1(n_1165),
.B2(n_1153),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1182),
.A2(n_1163),
.B1(n_1187),
.B2(n_1157),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1194),
.A2(n_1190),
.B1(n_1173),
.B2(n_1177),
.Y(n_1363)
);

INVx3_ASAP7_75t_SL g1364 ( 
.A(n_1194),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1177),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1290),
.A2(n_1258),
.B1(n_1276),
.B2(n_1269),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1245),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1155),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1279),
.A2(n_1257),
.B1(n_1280),
.B2(n_651),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1282),
.A2(n_436),
.B1(n_931),
.B2(n_651),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1282),
.A2(n_841),
.B1(n_651),
.B2(n_1257),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1256),
.A2(n_931),
.B1(n_827),
.B2(n_960),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1168),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1257),
.A2(n_841),
.B1(n_651),
.B2(n_750),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1234),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1199),
.B(n_1239),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1168),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1257),
.A2(n_651),
.B1(n_1167),
.B2(n_827),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1234),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1151),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1154),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1215),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1151),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_SL g1387 ( 
.A(n_1234),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1168),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1257),
.A2(n_841),
.B1(n_651),
.B2(n_750),
.Y(n_1390)
);

BUFx8_ASAP7_75t_SL g1391 ( 
.A(n_1250),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1168),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1234),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1168),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1234),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1151),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1250),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1151),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1252),
.B(n_1260),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1168),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1252),
.B(n_1260),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1234),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1252),
.B(n_1260),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1252),
.B(n_1260),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1256),
.A2(n_523),
.B(n_644),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1234),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1241),
.A2(n_1048),
.B1(n_1280),
.B2(n_1257),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1256),
.A2(n_931),
.B1(n_827),
.B2(n_960),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1236),
.A2(n_436),
.B1(n_931),
.B2(n_651),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1234),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1189),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1301),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1362),
.A2(n_1361),
.B(n_1352),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1399),
.B(n_1401),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1362),
.A2(n_1361),
.B(n_1352),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1306),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1360),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1360),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1298),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1353),
.A2(n_1357),
.B(n_1354),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1407),
.A2(n_1323),
.B(n_1373),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_R g1426 ( 
.A(n_1322),
.B(n_1400),
.Y(n_1426)
);

INVxp33_ASAP7_75t_L g1427 ( 
.A(n_1378),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1316),
.B(n_1364),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1305),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1328),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1363),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1363),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1340),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1353),
.A2(n_1354),
.B(n_1367),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1350),
.B(n_1312),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1341),
.B(n_1342),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1365),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1334),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1349),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1368),
.A2(n_1319),
.A3(n_1347),
.B(n_1355),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1346),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1313),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1348),
.A2(n_1344),
.B(n_1336),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1321),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1311),
.B(n_1384),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1312),
.B(n_1295),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1383),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1339),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1386),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1348),
.A2(n_1344),
.B(n_1336),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1337),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1396),
.Y(n_1453)
);

NAND2x1_ASAP7_75t_L g1454 ( 
.A(n_1368),
.B(n_1326),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1398),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1358),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1320),
.B(n_1327),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1358),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1359),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1345),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1295),
.B(n_1373),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1299),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1299),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1317),
.B(n_1372),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1311),
.B(n_1384),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1315),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1345),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1308),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1369),
.A2(n_1338),
.B(n_1308),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1376),
.A2(n_1402),
.B(n_1389),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1376),
.A2(n_1410),
.B(n_1379),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1369),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1379),
.B(n_1402),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1329),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1389),
.A2(n_1409),
.B1(n_1410),
.B2(n_1405),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1333),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1338),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_SL g1479 ( 
.A(n_1392),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1405),
.B(n_1409),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1296),
.B(n_1335),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1323),
.B(n_1371),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1397),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1296),
.B(n_1351),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1366),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1375),
.B(n_1390),
.C(n_1370),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1414),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1331),
.B(n_1302),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1331),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1381),
.Y(n_1490)
);

AOI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1411),
.A2(n_1324),
.B(n_1314),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1490),
.B(n_1325),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1490),
.B(n_1382),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1425),
.A2(n_1412),
.B1(n_1332),
.B2(n_1408),
.C(n_1395),
.Y(n_1494)
);

NOR2x1_ASAP7_75t_R g1495 ( 
.A(n_1419),
.B(n_1394),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_SL g1496 ( 
.A1(n_1476),
.A2(n_1310),
.B(n_1385),
.C(n_1343),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1476),
.A2(n_1413),
.B(n_1393),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_SL g1498 ( 
.A1(n_1486),
.A2(n_1464),
.B(n_1477),
.C(n_1468),
.Y(n_1498)
);

NAND2x1_ASAP7_75t_L g1499 ( 
.A(n_1436),
.B(n_1465),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1423),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_L g1501 ( 
.A(n_1457),
.B(n_1441),
.C(n_1474),
.Y(n_1501)
);

AO32x2_ASAP7_75t_L g1502 ( 
.A1(n_1452),
.A2(n_1318),
.A3(n_1300),
.B1(n_1303),
.B2(n_1380),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1457),
.A2(n_1297),
.B1(n_1377),
.B2(n_1387),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1427),
.B(n_1408),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1415),
.B(n_1413),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1436),
.A2(n_1393),
.B(n_1391),
.C(n_1387),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1428),
.B(n_1388),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1474),
.A2(n_1304),
.B1(n_1297),
.B2(n_1377),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1471),
.A2(n_1356),
.B(n_1307),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1416),
.A2(n_1356),
.B(n_1309),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1416),
.A2(n_1309),
.B(n_1403),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1459),
.B(n_1456),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1441),
.B(n_1488),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1429),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1429),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1422),
.B(n_1420),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1436),
.B(n_1491),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1438),
.Y(n_1520)
);

AO32x2_ASAP7_75t_L g1521 ( 
.A1(n_1452),
.A2(n_1487),
.A3(n_1458),
.B1(n_1456),
.B2(n_1431),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_SL g1522 ( 
.A(n_1436),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1480),
.A2(n_1482),
.B1(n_1461),
.B2(n_1435),
.C(n_1439),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1436),
.A2(n_1472),
.B(n_1470),
.Y(n_1525)
);

AND2x4_ASAP7_75t_SL g1526 ( 
.A(n_1484),
.B(n_1481),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1472),
.A2(n_1482),
.B1(n_1447),
.B2(n_1470),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1444),
.A2(n_1451),
.B(n_1472),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1420),
.B(n_1437),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1448),
.B(n_1450),
.Y(n_1530)
);

AO32x2_ASAP7_75t_L g1531 ( 
.A1(n_1487),
.A2(n_1431),
.A3(n_1432),
.B1(n_1470),
.B2(n_1440),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1491),
.B(n_1469),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1444),
.A2(n_1451),
.B(n_1469),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_SL g1534 ( 
.A1(n_1477),
.A2(n_1468),
.B(n_1462),
.C(n_1463),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1448),
.B(n_1450),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1430),
.A2(n_1417),
.B1(n_1421),
.B2(n_1447),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1454),
.B(n_1424),
.Y(n_1537)
);

AND2x2_ASAP7_75t_SL g1538 ( 
.A(n_1435),
.B(n_1478),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1430),
.B(n_1489),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1430),
.A2(n_1462),
.B1(n_1463),
.B2(n_1473),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1533),
.B(n_1432),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1424),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1501),
.B(n_1467),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1537),
.B(n_1418),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1516),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1532),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1485),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1521),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1523),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1521),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1529),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1527),
.A2(n_1478),
.B(n_1473),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1418),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1532),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1519),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1535),
.Y(n_1563)
);

AOI221x1_ASAP7_75t_SL g1564 ( 
.A1(n_1536),
.A2(n_1540),
.B1(n_1514),
.B2(n_1503),
.C(n_1518),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1539),
.B(n_1440),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1499),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1531),
.B(n_1434),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1558),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1550),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1548),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1562),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1558),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1567),
.B(n_1511),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1561),
.B(n_1513),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1548),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1566),
.B(n_1526),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1549),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1549),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1566),
.Y(n_1580)
);

NAND4xp25_ASAP7_75t_SL g1581 ( 
.A(n_1564),
.B(n_1494),
.C(n_1524),
.D(n_1525),
.Y(n_1581)
);

AND2x4_ASAP7_75t_SL g1582 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1563),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1567),
.B(n_1511),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_L g1585 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1440),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1544),
.A2(n_1498),
.A3(n_1534),
.B(n_1540),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1567),
.B(n_1531),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1542),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1546),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1531),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1559),
.A2(n_1506),
.B(n_1497),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1563),
.B(n_1513),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1566),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1552),
.B(n_1531),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1566),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1562),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1589),
.B(n_1542),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1585),
.B(n_1545),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1589),
.B(n_1542),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1553),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1570),
.B(n_1565),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1590),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1596),
.B(n_1566),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1590),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1569),
.B(n_1565),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1593),
.B(n_1565),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1556),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1578),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1587),
.B(n_1551),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1581),
.A2(n_1564),
.B1(n_1559),
.B2(n_1498),
.C(n_1544),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1579),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1572),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1592),
.A2(n_1493),
.B(n_1534),
.C(n_1496),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1605),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1622),
.B(n_1594),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1612),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1624),
.A2(n_1587),
.B(n_1592),
.C(n_1520),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1609),
.B(n_1586),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1586),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1616),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1613),
.B(n_1615),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1588),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1598),
.B(n_1588),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1613),
.A2(n_1581),
.B1(n_1522),
.B2(n_1512),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1616),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1568),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1618),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1588),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1599),
.B(n_1433),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1621),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1621),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1602),
.B(n_1591),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1625),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.B(n_1573),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1606),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1600),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1607),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1627),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1628),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1573),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1606),
.B(n_1573),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1603),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1629),
.B(n_1585),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1667),
.B(n_1608),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1671),
.B(n_1599),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1667),
.B(n_1603),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1671),
.B(n_1610),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1653),
.B(n_1622),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1653),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1670),
.B(n_1601),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1672),
.B(n_1611),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1611),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1632),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1601),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1633),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1641),
.B(n_1626),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1633),
.B(n_1492),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1641),
.B(n_1626),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1670),
.B(n_1614),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1662),
.B(n_1606),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1635),
.B(n_1495),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1639),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1635),
.B(n_1596),
.C(n_1510),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1639),
.B(n_1597),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1641),
.B(n_1600),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1639),
.B(n_1597),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1646),
.A2(n_1560),
.B(n_1547),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1632),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1433),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1662),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1656),
.B(n_1614),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1604),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1634),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1661),
.B(n_1600),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1631),
.B(n_1509),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1631),
.B(n_1509),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1642),
.B(n_1604),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1630),
.Y(n_1708)
);

OAI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1697),
.A2(n_1693),
.B1(n_1679),
.B2(n_1691),
.C(n_1681),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1700),
.A2(n_1682),
.B1(n_1706),
.B2(n_1705),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1699),
.A2(n_1507),
.B(n_1661),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1433),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1687),
.B(n_1648),
.Y(n_1713)
);

AOI21xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1673),
.A2(n_1507),
.B(n_1661),
.Y(n_1714)
);

AOI211x1_ASAP7_75t_SL g1715 ( 
.A1(n_1685),
.A2(n_1651),
.B(n_1642),
.C(n_1643),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1677),
.A2(n_1668),
.B1(n_1648),
.B2(n_1659),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1717)
);

OAI32xp33_ASAP7_75t_L g1718 ( 
.A1(n_1678),
.A2(n_1663),
.A3(n_1651),
.B1(n_1643),
.B2(n_1669),
.Y(n_1718)
);

NAND2xp33_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1572),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1686),
.B(n_1648),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1690),
.A2(n_1663),
.B(n_1669),
.Y(n_1721)
);

OAI31xp33_ASAP7_75t_L g1722 ( 
.A1(n_1690),
.A2(n_1558),
.A3(n_1445),
.B(n_1466),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1703),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1695),
.A2(n_1668),
.B1(n_1659),
.B2(n_1663),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1694),
.Y(n_1725)
);

OAI32xp33_ASAP7_75t_L g1726 ( 
.A1(n_1696),
.A2(n_1669),
.A3(n_1668),
.B1(n_1659),
.B2(n_1637),
.Y(n_1726)
);

NAND4xp25_ASAP7_75t_L g1727 ( 
.A(n_1684),
.B(n_1508),
.C(n_1541),
.D(n_1445),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1686),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1695),
.A2(n_1538),
.B1(n_1596),
.B2(n_1558),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1688),
.A2(n_1560),
.B1(n_1538),
.B2(n_1551),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1685),
.B(n_1594),
.C(n_1634),
.Y(n_1731)
);

AOI322xp5_ASAP7_75t_L g1732 ( 
.A1(n_1688),
.A2(n_1591),
.A3(n_1595),
.B1(n_1584),
.B2(n_1574),
.C1(n_1555),
.C2(n_1554),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1692),
.B(n_1640),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.B(n_1620),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1709),
.A2(n_1676),
.B(n_1698),
.C(n_1683),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1704),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1723),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1712),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1717),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1716),
.B(n_1704),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1719),
.A2(n_1680),
.B1(n_1674),
.B2(n_1702),
.C(n_1707),
.Y(n_1741)
);

AO22x2_ASAP7_75t_L g1742 ( 
.A1(n_1710),
.A2(n_1703),
.B1(n_1708),
.B2(n_1674),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1725),
.B(n_1680),
.C(n_1708),
.Y(n_1743)
);

AOI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1718),
.A2(n_1702),
.B(n_1707),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1733),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1717),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1721),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1720),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1724),
.A2(n_1594),
.B1(n_1560),
.B2(n_1596),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1734),
.Y(n_1750)
);

AOI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1726),
.A2(n_1595),
.B1(n_1666),
.B2(n_1652),
.C1(n_1664),
.C2(n_1640),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1715),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1714),
.A2(n_1701),
.B1(n_1689),
.B2(n_1666),
.C(n_1647),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1711),
.B(n_1647),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1737),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1727),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1750),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1736),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1739),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1739),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1738),
.B(n_1753),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1740),
.B(n_1731),
.Y(n_1763)
);

XNOR2x1_ASAP7_75t_SL g1764 ( 
.A(n_1742),
.B(n_1479),
.Y(n_1764)
);

NOR2x1_ASAP7_75t_SL g1765 ( 
.A(n_1745),
.B(n_1460),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1751),
.A2(n_1722),
.B(n_1729),
.C(n_1732),
.Y(n_1766)
);

NOR4xp25_ASAP7_75t_L g1767 ( 
.A(n_1761),
.B(n_1735),
.C(n_1747),
.D(n_1741),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1760),
.B(n_1748),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1763),
.B(n_1752),
.Y(n_1769)
);

NAND4xp25_ASAP7_75t_L g1770 ( 
.A(n_1762),
.B(n_1751),
.C(n_1743),
.D(n_1744),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1759),
.B(n_1755),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1755),
.Y(n_1773)
);

NOR3x1_ASAP7_75t_L g1774 ( 
.A(n_1757),
.B(n_1701),
.C(n_1689),
.Y(n_1774)
);

OAI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1766),
.A2(n_1744),
.B(n_1722),
.C(n_1754),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1758),
.B(n_1749),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1769),
.B(n_1765),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_SL g1778 ( 
.A1(n_1775),
.A2(n_1764),
.B(n_1776),
.C(n_1771),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1767),
.A2(n_1764),
.B(n_1756),
.C(n_1765),
.Y(n_1779)
);

AOI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1770),
.A2(n_1460),
.B(n_1426),
.C(n_1475),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1770),
.A2(n_1652),
.B(n_1650),
.Y(n_1781)
);

NAND4xp25_ASAP7_75t_L g1782 ( 
.A(n_1780),
.B(n_1774),
.C(n_1772),
.D(n_1768),
.Y(n_1782)
);

AOI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1779),
.A2(n_1773),
.B(n_1730),
.Y(n_1783)
);

OAI322xp33_ASAP7_75t_L g1784 ( 
.A1(n_1781),
.A2(n_1665),
.A3(n_1630),
.B1(n_1660),
.B2(n_1638),
.C1(n_1644),
.C2(n_1649),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1777),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1778),
.B(n_1502),
.C(n_1630),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1778),
.A2(n_1654),
.B1(n_1664),
.B2(n_1650),
.C(n_1658),
.Y(n_1787)
);

NOR2xp67_ASAP7_75t_L g1788 ( 
.A(n_1782),
.B(n_1654),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1785),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1786),
.Y(n_1790)
);

INVx5_ASAP7_75t_L g1791 ( 
.A(n_1783),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1787),
.B(n_1636),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1789),
.B(n_1460),
.Y(n_1793)
);

NAND4xp75_ASAP7_75t_L g1794 ( 
.A(n_1788),
.B(n_1784),
.C(n_1655),
.D(n_1657),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1792),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_SL g1796 ( 
.A(n_1795),
.B(n_1791),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1790),
.B1(n_1791),
.B2(n_1794),
.Y(n_1797)
);

OAI22x1_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1793),
.B1(n_1665),
.B2(n_1660),
.Y(n_1798)
);

AOI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1797),
.A2(n_1644),
.B(n_1638),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1798),
.B(n_1638),
.Y(n_1800)
);

OAI22x1_ASAP7_75t_L g1801 ( 
.A1(n_1799),
.A2(n_1665),
.B1(n_1660),
.B2(n_1649),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1800),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1657),
.B(n_1655),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1802),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1803),
.B1(n_1649),
.B2(n_1644),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1805),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1658),
.B1(n_1475),
.B2(n_1505),
.C(n_1504),
.Y(n_1807)
);

OAI31xp33_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1475),
.A3(n_1502),
.B(n_1446),
.Y(n_1808)
);


endmodule