module fake_jpeg_3762_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp33_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_48),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_56),
.Y(n_85)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_34),
.B1(n_21),
.B2(n_20),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_52),
.Y(n_77)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_76),
.B1(n_83),
.B2(n_88),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_27),
.C(n_31),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_3),
.C(n_6),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_78),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_17),
.B1(n_33),
.B2(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_42),
.B(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_51),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_40),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_24),
.B1(n_19),
.B2(n_34),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_84),
.B1(n_91),
.B2(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_120),
.B1(n_87),
.B2(n_90),
.Y(n_147)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_51),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_109),
.B(n_96),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_57),
.B1(n_48),
.B2(n_44),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_124),
.B(n_90),
.C(n_75),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_96),
.CI(n_75),
.CON(n_148),
.SN(n_148)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_118),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_43),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_112),
.B1(n_70),
.B2(n_80),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_44),
.B1(n_43),
.B2(n_10),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_65),
.B(n_79),
.C(n_69),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_10),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_11),
.C(n_12),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_96),
.C(n_113),
.Y(n_151)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_12),
.B1(n_69),
.B2(n_70),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_115),
.B1(n_104),
.B2(n_109),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_141),
.B1(n_152),
.B2(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_77),
.Y(n_139)
);

OAI22x1_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_98),
.B1(n_112),
.B2(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_116),
.B(n_126),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_117),
.B(n_108),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_121),
.B1(n_117),
.B2(n_106),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_149),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_138),
.B(n_140),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_163),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_140),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_122),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_161),
.C(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_108),
.C(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_133),
.B1(n_143),
.B2(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_133),
.C(n_145),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_148),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_144),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_186),
.B(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_191),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_187),
.CI(n_188),
.CON(n_198),
.SN(n_198)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_167),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_181),
.C(n_178),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_142),
.B(n_146),
.Y(n_187)
);

NOR4xp25_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_172),
.C(n_162),
.D(n_174),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_142),
.B(n_129),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_172),
.B1(n_154),
.B2(n_162),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_156),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_201),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_190),
.CI(n_176),
.CON(n_210),
.SN(n_210)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_157),
.B1(n_165),
.B2(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_202),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_170),
.B1(n_168),
.B2(n_175),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_182),
.B1(n_192),
.B2(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_189),
.B1(n_203),
.B2(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_216),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_215),
.B(n_210),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_180),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.C(n_212),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_206),
.A3(n_198),
.B1(n_200),
.B2(n_197),
.C1(n_196),
.C2(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_203),
.B1(n_202),
.B2(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_220),
.B1(n_214),
.B2(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_203),
.B1(n_194),
.B2(n_198),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_204),
.B1(n_205),
.B2(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_229),
.B(n_227),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_221),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_226),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_234),
.B(n_231),
.Y(n_238)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_224),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_238),
.B(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.Y(n_242)
);


endmodule