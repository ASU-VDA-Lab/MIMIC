module fake_jpeg_30075_n_260 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_26),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_67),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_29),
.B1(n_17),
.B2(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_85),
.B1(n_2),
.B2(n_6),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_29),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_30),
.B(n_35),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_71),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_34),
.Y(n_71)
);

BUFx2_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_87),
.B(n_90),
.C(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_75),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_34),
.B1(n_27),
.B2(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_35),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_37),
.A2(n_33),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_37),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_38),
.B(n_22),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_28),
.B1(n_2),
.B2(n_6),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_10),
.B1(n_72),
.B2(n_59),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_1),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_107),
.B1(n_121),
.B2(n_84),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_57),
.Y(n_150)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_115),
.Y(n_153)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx24_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_10),
.B1(n_92),
.B2(n_80),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_137),
.B1(n_150),
.B2(n_114),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_66),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_94),
.B1(n_70),
.B2(n_60),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_109),
.B1(n_126),
.B2(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_82),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_139),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_98),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_141),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_70),
.B1(n_94),
.B2(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_57),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_77),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_91),
.C(n_71),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_77),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_71),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_91),
.CI(n_99),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_81),
.C(n_83),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_101),
.B(n_96),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_181),
.B1(n_148),
.B2(n_156),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_171),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_107),
.B1(n_127),
.B2(n_99),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_R g203 ( 
.A1(n_168),
.A2(n_179),
.B(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_184),
.B1(n_168),
.B2(n_155),
.Y(n_191)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_129),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_174),
.Y(n_205)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_122),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_132),
.A2(n_109),
.B1(n_107),
.B2(n_120),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_184),
.B(n_169),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_108),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_96),
.B1(n_105),
.B2(n_102),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_124),
.B1(n_112),
.B2(n_99),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_108),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_144),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_132),
.B1(n_154),
.B2(n_131),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_164),
.B1(n_178),
.B2(n_176),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_158),
.C(n_143),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_195),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_146),
.C(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_156),
.B1(n_160),
.B2(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.C(n_182),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_187),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_170),
.B(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_166),
.B1(n_161),
.B2(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_212),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_172),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_170),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_216),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_192),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_188),
.C(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_195),
.Y(n_223)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_194),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_206),
.B1(n_193),
.B2(n_190),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_218),
.B1(n_217),
.B2(n_211),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_232),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_237),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_236),
.B1(n_226),
.B2(n_228),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_212),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_213),
.C(n_222),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_213),
.C(n_235),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_223),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_244),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_227),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_247),
.C(n_236),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_221),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_191),
.C(n_172),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_238),
.A3(n_228),
.B1(n_224),
.B2(n_231),
.C1(n_234),
.C2(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_225),
.B1(n_219),
.B2(n_204),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_245),
.B(n_246),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_248),
.B(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_254),
.B(n_248),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_257),
.B(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_167),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_167),
.Y(n_260)
);


endmodule