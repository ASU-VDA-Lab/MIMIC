module fake_jpeg_21673_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_11),
.B(n_30),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_58),
.B1(n_77),
.B2(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_98),
.B1(n_53),
.B2(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_61),
.C(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_84),
.B1(n_88),
.B2(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_108),
.B1(n_92),
.B2(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_74),
.B1(n_63),
.B2(n_68),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_58),
.B1(n_83),
.B2(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_112),
.B1(n_64),
.B2(n_66),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_50),
.B1(n_81),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_129),
.B1(n_60),
.B2(n_1),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_124),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_76),
.B(n_53),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_56),
.B(n_70),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_64),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_71),
.B1(n_68),
.B2(n_63),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_75),
.B1(n_59),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_72),
.B1(n_73),
.B2(n_57),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_136),
.B1(n_140),
.B2(n_129),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_69),
.B1(n_65),
.B2(n_62),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_4),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_5),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_145),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_115),
.A3(n_121),
.B1(n_23),
.B2(n_48),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_154),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_21),
.B(n_47),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_127),
.B1(n_7),
.B2(n_8),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_18),
.B(n_43),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_137),
.CI(n_143),
.CON(n_159),
.SN(n_159)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_146),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_159),
.C(n_157),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_160),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_158),
.B1(n_155),
.B2(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_154),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_136),
.B(n_7),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_16),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_22),
.B(n_41),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_14),
.B(n_40),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_44),
.B(n_36),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_26),
.B(n_8),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_6),
.Y(n_175)
);


endmodule