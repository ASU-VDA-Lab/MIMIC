module fake_jpeg_1486_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_67),
.B1(n_64),
.B2(n_53),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_70),
.B1(n_52),
.B2(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_54),
.B1(n_65),
.B2(n_58),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_88),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

NAND2xp67_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_68),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_73),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_72),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_76),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_69),
.B(n_70),
.C(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_99),
.B1(n_59),
.B2(n_4),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_58),
.B1(n_60),
.B2(n_55),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_80),
.B1(n_55),
.B2(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_118),
.B1(n_121),
.B2(n_2),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_1),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_1),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_59),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_103),
.C(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_59),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_96),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_37),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_19),
.C(n_47),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_144),
.C(n_146),
.Y(n_166)
);

CKINVDCx12_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_10),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_2),
.B(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_49),
.B(n_45),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_147),
.B(n_34),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_10),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_44),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_108),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_43),
.B(n_41),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_125),
.B1(n_118),
.B2(n_111),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_151),
.B1(n_161),
.B2(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_153),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_124),
.B1(n_7),
.B2(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_6),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_147),
.B1(n_137),
.B2(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_9),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.C(n_14),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_159),
.B1(n_166),
.B2(n_13),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_35),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_33),
.B(n_29),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_165),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_187)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_176),
.B(n_175),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_149),
.B1(n_151),
.B2(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_159),
.B(n_12),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.B(n_177),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_193),
.B1(n_185),
.B2(n_172),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_185),
.C(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_196),
.C(n_191),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_181),
.B(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_188),
.B(n_190),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_198),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_11),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_15),
.C(n_16),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_202),
.B(n_17),
.CI(n_18),
.CON(n_203),
.SN(n_203)
);


endmodule