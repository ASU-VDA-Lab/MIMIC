module fake_jpeg_16370_n_375 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_38),
.B(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_61),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_56),
.Y(n_86)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_16),
.B(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_65),
.Y(n_100)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_37),
.B1(n_15),
.B2(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_76),
.B1(n_81),
.B2(n_85),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_18),
.B1(n_16),
.B2(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_89),
.B1(n_44),
.B2(n_51),
.Y(n_129)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_17),
.B1(n_32),
.B2(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_66),
.B1(n_61),
.B2(n_56),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_36),
.B(n_32),
.C(n_25),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_83),
.A2(n_26),
.B(n_19),
.C(n_21),
.Y(n_154)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_36),
.B1(n_24),
.B2(n_20),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_24),
.B1(n_20),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_87),
.A2(n_93),
.B1(n_34),
.B2(n_26),
.Y(n_136)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_30),
.B1(n_19),
.B2(n_34),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_30),
.B1(n_34),
.B2(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_112),
.Y(n_126)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_13),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_108),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_41),
.B(n_12),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_31),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_50),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_116),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_55),
.B1(n_46),
.B2(n_62),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_136),
.B1(n_164),
.B2(n_137),
.Y(n_180)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_128),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_90),
.B1(n_99),
.B2(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_123),
.A2(n_138),
.B1(n_167),
.B2(n_21),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_132),
.Y(n_184)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_130),
.A2(n_150),
.B1(n_159),
.B2(n_109),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_134),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_62),
.B1(n_58),
.B2(n_26),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_140),
.Y(n_195)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx6p67_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_31),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_31),
.Y(n_145)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_155),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_101),
.B1(n_111),
.B2(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_74),
.Y(n_151)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_91),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

OR2x4_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_9),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_12),
.C(n_2),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g209 ( 
.A(n_156),
.B(n_160),
.Y(n_209)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_96),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_1),
.C(n_2),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_31),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_58),
.B1(n_21),
.B2(n_4),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_73),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_183),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_73),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_189),
.B(n_139),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_125),
.B(n_73),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_175),
.B(n_201),
.Y(n_251)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_186),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_72),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_206),
.B(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_121),
.A2(n_67),
.B1(n_116),
.B2(n_75),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_210),
.B(n_206),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_162),
.C(n_131),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_181),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_198),
.B1(n_158),
.B2(n_146),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_80),
.C(n_104),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_154),
.Y(n_183)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_83),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_109),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_161),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_141),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_118),
.B(n_166),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_5),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_129),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_205),
.B1(n_211),
.B2(n_130),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_119),
.A2(n_54),
.B1(n_21),
.B2(n_10),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_7),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_124),
.B(n_9),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_119),
.A2(n_10),
.B1(n_148),
.B2(n_122),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_149),
.A2(n_10),
.B(n_124),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_219),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_230),
.B(n_250),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_226),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_234),
.B(n_235),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_222),
.A2(n_237),
.B1(n_248),
.B2(n_195),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_230),
.B(n_233),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_232),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_139),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_174),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_169),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_142),
.B(n_118),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_148),
.B(n_143),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_146),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_143),
.C(n_161),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_236),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_196),
.B(n_179),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_244),
.B(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_184),
.A2(n_143),
.B1(n_140),
.B2(n_127),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_249),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_178),
.B1(n_189),
.B2(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_168),
.B(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_172),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_188),
.A2(n_206),
.B1(n_211),
.B2(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_182),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_213),
.B1(n_203),
.B2(n_190),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_192),
.B1(n_190),
.B2(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_200),
.B(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_192),
.B(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_229),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_254),
.B(n_255),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_209),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_272),
.C(n_275),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_215),
.A2(n_195),
.B1(n_170),
.B2(n_187),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_276),
.B1(n_230),
.B2(n_220),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_252),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_267),
.B(n_285),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_176),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_268),
.B(n_282),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_274),
.B1(n_238),
.B2(n_244),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_280),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_186),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_170),
.B1(n_234),
.B2(n_222),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_236),
.A2(n_243),
.B1(n_226),
.B2(n_232),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_235),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_279),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_248),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_230),
.A2(n_227),
.B1(n_246),
.B2(n_223),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_233),
.B(n_283),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_247),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_241),
.B1(n_242),
.B2(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_277),
.B1(n_265),
.B2(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_218),
.B(n_228),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_293),
.B(n_303),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_294),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_239),
.B(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_259),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_296),
.C(n_308),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_251),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_276),
.B1(n_285),
.B2(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_305),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_263),
.B1(n_254),
.B2(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_270),
.A2(n_258),
.B1(n_283),
.B2(n_286),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_307),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_256),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_280),
.B(n_279),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_303),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_255),
.A2(n_261),
.B1(n_260),
.B2(n_257),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_271),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_319),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_330),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_327),
.C(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_295),
.C(n_296),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_297),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_311),
.C(n_301),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_332),
.C(n_290),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_298),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_318),
.B1(n_331),
.B2(n_333),
.Y(n_334)
);

OAI22x1_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_346),
.B1(n_287),
.B2(n_316),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_313),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_293),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_345),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_324),
.B(n_302),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_326),
.B(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_340),
.B(n_344),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_294),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_348),
.B(n_341),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_300),
.CI(n_288),
.CON(n_344),
.SN(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_325),
.B1(n_322),
.B2(n_328),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_317),
.B(n_309),
.Y(n_347)
);

NAND4xp25_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_344),
.C(n_336),
.D(n_334),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_287),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_SL g350 ( 
.A(n_348),
.B(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_357),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_352),
.A2(n_353),
.B(n_349),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_343),
.A2(n_323),
.B(n_327),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_316),
.C(n_337),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_337),
.C(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_344),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_360),
.B(n_364),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_346),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_363),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_342),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_365),
.A2(n_352),
.B(n_357),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_362),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_355),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_369),
.A2(n_370),
.B(n_367),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_371),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_365),
.B(n_364),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_362),
.C(n_353),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_354),
.Y(n_375)
);


endmodule