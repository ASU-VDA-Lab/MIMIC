module fake_jpeg_29625_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_20),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_22),
.Y(n_64)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_38),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_68),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_39),
.B1(n_29),
.B2(n_40),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_76),
.B1(n_71),
.B2(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_66),
.Y(n_85)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_77),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_13),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_25),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_74),
.B(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_33),
.B(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_76)
);

FAx1_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_33),
.CI(n_28),
.CON(n_77),
.SN(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_56),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_42),
.B(n_56),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_88),
.B1(n_77),
.B2(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_91),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_60),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_11),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_81),
.C(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_77),
.C(n_74),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_106),
.C(n_82),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_105),
.B1(n_83),
.B2(n_85),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_76),
.B1(n_69),
.B2(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_0),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_85),
.B(n_79),
.C(n_84),
.D(n_91),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_88),
.B1(n_80),
.B2(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_6),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_115),
.B(n_10),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_106),
.C(n_101),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_119),
.C(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_121),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_103),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_98),
.B1(n_109),
.B2(n_110),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_104),
.B1(n_99),
.B2(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_10),
.C(n_2),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_132),
.A3(n_130),
.B1(n_119),
.B2(n_127),
.C1(n_3),
.C2(n_1),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_135),
.Y(n_139)
);


endmodule