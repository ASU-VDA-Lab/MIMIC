module real_aes_18219_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_884;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g118 ( .A(n_0), .B(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_1), .A2(n_4), .B1(n_291), .B2(n_292), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_2), .A2(n_44), .B1(n_162), .B2(n_191), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_3), .A2(n_24), .B1(n_191), .B2(n_272), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_5), .A2(n_16), .B1(n_552), .B2(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_6), .A2(n_30), .B1(n_146), .B2(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_6), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_7), .A2(n_60), .B1(n_199), .B2(n_228), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_8), .A2(n_17), .B1(n_162), .B2(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_10), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_11), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_12), .A2(n_18), .B1(n_573), .B2(n_574), .Y(n_572) );
OR2x2_ASAP7_75t_L g126 ( .A(n_13), .B(n_38), .Y(n_126) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_14), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_15), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_19), .A2(n_101), .B1(n_292), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_20), .A2(n_39), .B1(n_234), .B2(n_609), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_21), .B(n_233), .Y(n_606) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_22), .A2(n_58), .B(n_175), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_23), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_25), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_26), .B(n_167), .Y(n_247) );
INVx4_ASAP7_75t_R g215 ( .A(n_27), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_28), .A2(n_48), .B1(n_169), .B2(n_289), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_29), .A2(n_54), .B1(n_169), .B2(n_552), .Y(n_562) );
INVx1_ASAP7_75t_L g146 ( .A(n_30), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_31), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_32), .B(n_609), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_33), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_34), .B(n_191), .Y(n_254) );
INVx1_ASAP7_75t_L g296 ( .A(n_35), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_SL g269 ( .A1(n_36), .A2(n_162), .B(n_166), .C(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_37), .A2(n_55), .B1(n_162), .B2(n_169), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_40), .A2(n_87), .B1(n_162), .B2(n_618), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_41), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_42), .A2(n_47), .B1(n_162), .B2(n_164), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_43), .A2(n_144), .B1(n_145), .B2(n_148), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_43), .Y(n_148) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_45), .A2(n_68), .B1(n_887), .B2(n_888), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_45), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_46), .A2(n_59), .B1(n_552), .B2(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g251 ( .A(n_49), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_50), .B(n_162), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_51), .Y(n_189) );
INVx2_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
INVx1_ASAP7_75t_L g124 ( .A(n_53), .Y(n_124) );
BUFx3_ASAP7_75t_L g139 ( .A(n_53), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_56), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_57), .A2(n_89), .B1(n_162), .B2(n_169), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_61), .A2(n_75), .B1(n_289), .B2(n_554), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_62), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_63), .A2(n_78), .B1(n_162), .B2(n_164), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_64), .A2(n_99), .B1(n_552), .B2(n_574), .Y(n_595) );
INVx1_ASAP7_75t_L g175 ( .A(n_65), .Y(n_175) );
AND2x4_ASAP7_75t_L g177 ( .A(n_66), .B(n_178), .Y(n_177) );
OA22x2_ASAP7_75t_L g141 ( .A1(n_67), .A2(n_142), .B1(n_143), .B2(n_149), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_67), .Y(n_142) );
INVx1_ASAP7_75t_L g887 ( .A(n_68), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_69), .A2(n_92), .B1(n_169), .B2(n_289), .Y(n_288) );
AO22x1_ASAP7_75t_L g231 ( .A1(n_70), .A2(n_76), .B1(n_232), .B2(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g178 ( .A(n_71), .Y(n_178) );
AND2x2_ASAP7_75t_L g273 ( .A(n_72), .B(n_185), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_73), .B(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_74), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_77), .B(n_191), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g882 ( .A1(n_79), .A2(n_128), .B1(n_883), .B2(n_884), .Y(n_882) );
CKINVDCx14_ASAP7_75t_R g883 ( .A(n_79), .Y(n_883) );
INVx2_ASAP7_75t_L g167 ( .A(n_80), .Y(n_167) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_81), .B(n_185), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_82), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_83), .A2(n_100), .B1(n_169), .B2(n_199), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_84), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_85), .B(n_173), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_86), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_88), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_90), .Y(n_866) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_91), .B(n_185), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_93), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_94), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_95), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g539 ( .A(n_95), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g610 ( .A(n_96), .B(n_233), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_97), .A2(n_171), .B(n_199), .C(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g219 ( .A(n_98), .B(n_220), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_102), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_877), .Y(n_103) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_132), .B1(n_873), .B2(n_874), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_110), .B(n_116), .Y(n_115) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_111), .B(n_120), .Y(n_131) );
INVx1_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_111), .B(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_112), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_127), .Y(n_112) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_120), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x4_ASAP7_75t_L g130 ( .A(n_116), .B(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g875 ( .A(n_118), .B(n_876), .Y(n_875) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx5_ASAP7_75t_L g876 ( .A(n_121), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_121), .Y(n_880) );
CKINVDCx8_ASAP7_75t_R g892 ( .A(n_121), .Y(n_892) );
AND2x6_ASAP7_75t_SL g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_125), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2x1_ASAP7_75t_L g872 ( .A(n_126), .B(n_139), .Y(n_872) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_127), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_128), .Y(n_884) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI21xp33_ASAP7_75t_L g877 ( .A1(n_132), .A2(n_874), .B(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_865), .Y(n_133) );
BUFx12f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_864), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_141), .B(n_150), .Y(n_864) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_536), .B1(n_540), .B2(n_861), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_445), .Y(n_151) );
NOR3xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_361), .C(n_392), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_327), .Y(n_153) );
AOI211x1_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_239), .B(n_282), .C(n_313), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_203), .Y(n_156) );
AND2x2_ASAP7_75t_L g468 ( .A(n_157), .B(n_343), .Y(n_468) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_182), .Y(n_157) );
INVx1_ASAP7_75t_L g353 ( .A(n_158), .Y(n_353) );
OR2x2_ASAP7_75t_L g474 ( .A(n_158), .B(n_325), .Y(n_474) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g310 ( .A(n_159), .B(n_183), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_159), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g342 ( .A(n_159), .Y(n_342) );
OR2x2_ASAP7_75t_L g373 ( .A(n_159), .B(n_204), .Y(n_373) );
AND2x2_ASAP7_75t_L g387 ( .A(n_159), .B(n_204), .Y(n_387) );
AND2x2_ASAP7_75t_L g424 ( .A(n_159), .B(n_380), .Y(n_424) );
AO31x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_172), .A3(n_176), .B(n_179), .Y(n_159) );
OAI22x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_165), .B1(n_168), .B2(n_170), .Y(n_160) );
INVx4_ASAP7_75t_L g164 ( .A(n_162), .Y(n_164) );
INVx1_ASAP7_75t_L g554 ( .A(n_162), .Y(n_554) );
INVx1_ASAP7_75t_L g574 ( .A(n_162), .Y(n_574) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx1_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx1_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_163), .Y(n_233) );
INVx1_ASAP7_75t_L g235 ( .A(n_163), .Y(n_235) );
INVx1_ASAP7_75t_L g266 ( .A(n_163), .Y(n_266) );
INVx2_ASAP7_75t_L g272 ( .A(n_163), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_164), .A2(n_189), .B(n_190), .C(n_192), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_L g604 ( .A1(n_164), .A2(n_166), .B(n_605), .C(n_606), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_165), .A2(n_225), .B1(n_277), .B2(n_278), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_165), .A2(n_170), .B1(n_288), .B2(n_290), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_165), .A2(n_551), .B1(n_553), .B2(n_555), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_165), .A2(n_555), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_165), .A2(n_572), .B1(n_575), .B2(n_576), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_165), .A2(n_555), .B1(n_587), .B2(n_588), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_165), .A2(n_576), .B1(n_595), .B2(n_596), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_165), .A2(n_608), .B(n_610), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_165), .A2(n_170), .B1(n_617), .B2(n_619), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_165), .A2(n_555), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_166), .A2(n_196), .B(n_198), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_166), .B(n_231), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_166), .A2(n_224), .B(n_231), .C(n_237), .Y(n_326) );
BUFx8_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
INVx2_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
INVx1_ASAP7_75t_L g250 ( .A(n_167), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_169), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g291 ( .A(n_169), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_170), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_SL g576 ( .A(n_171), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_172), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_172), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g181 ( .A(n_173), .Y(n_181) );
INVx2_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
OAI21xp33_ASAP7_75t_L g237 ( .A1(n_173), .A2(n_229), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_174), .Y(n_186) );
INVx2_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_176), .A2(n_260), .A3(n_571), .B(n_577), .Y(n_570) );
AO31x2_ASAP7_75t_L g585 ( .A1(n_176), .A2(n_279), .A3(n_586), .B(n_589), .Y(n_585) );
AO31x2_ASAP7_75t_L g631 ( .A1(n_176), .A2(n_615), .A3(n_632), .B(n_636), .Y(n_631) );
BUFx10_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx10_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
INVx1_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
INVx1_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx2_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
BUFx2_ASAP7_75t_L g260 ( .A(n_181), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_181), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_181), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g304 ( .A(n_182), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_182), .B(n_221), .Y(n_355) );
AND2x2_ASAP7_75t_L g498 ( .A(n_182), .B(n_204), .Y(n_498) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx3_ASAP7_75t_L g322 ( .A(n_183), .Y(n_322) );
AND2x2_ASAP7_75t_L g341 ( .A(n_183), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g378 ( .A(n_183), .Y(n_378) );
AND2x2_ASAP7_75t_L g402 ( .A(n_183), .B(n_204), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_184), .B(n_187), .Y(n_183) );
NOR2x1_ASAP7_75t_L g200 ( .A(n_185), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g279 ( .A(n_185), .Y(n_279) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g255 ( .A(n_186), .B(n_202), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_186), .B(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_186), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g602 ( .A(n_186), .Y(n_602) );
BUFx3_ASAP7_75t_L g615 ( .A(n_186), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_186), .B(n_637), .Y(n_636) );
OAI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_195), .B(n_200), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_191), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx3_ASAP7_75t_L g226 ( .A(n_194), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g214 ( .A1(n_197), .A2(n_215), .B1(n_216), .B2(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g289 ( .A(n_197), .Y(n_289) );
INVx1_ASAP7_75t_L g609 ( .A(n_197), .Y(n_609) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AO31x2_ASAP7_75t_L g275 ( .A1(n_202), .A2(n_276), .A3(n_279), .B(n_280), .Y(n_275) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_203), .Y(n_302) );
AND2x2_ASAP7_75t_L g363 ( .A(n_203), .B(n_352), .Y(n_363) );
INVx2_ASAP7_75t_L g495 ( .A(n_203), .Y(n_495) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_221), .Y(n_203) );
INVx1_ASAP7_75t_L g300 ( .A(n_204), .Y(n_300) );
AND2x4_ASAP7_75t_L g312 ( .A(n_204), .B(n_222), .Y(n_312) );
INVx2_ASAP7_75t_L g380 ( .A(n_204), .Y(n_380) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_208), .B(n_219), .Y(n_204) );
AO31x2_ASAP7_75t_L g548 ( .A1(n_205), .A2(n_549), .A3(n_550), .B(n_556), .Y(n_548) );
AO31x2_ASAP7_75t_L g559 ( .A1(n_205), .A2(n_293), .A3(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_SL g577 ( .A(n_207), .B(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_207), .B(n_621), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_213), .B(n_218), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
INVx1_ASAP7_75t_L g635 ( .A(n_216), .Y(n_635) );
INVx1_ASAP7_75t_L g549 ( .A(n_218), .Y(n_549) );
AND2x2_ASAP7_75t_L g379 ( .A(n_221), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g386 ( .A(n_221), .Y(n_386) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g464 ( .A(n_222), .B(n_380), .Y(n_464) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_230), .B(n_236), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_229), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_225), .A2(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g555 ( .A(n_226), .Y(n_555) );
INVx1_ASAP7_75t_L g573 ( .A(n_228), .Y(n_573) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g552 ( .A(n_233), .Y(n_552) );
OAI21xp33_ASAP7_75t_SL g246 ( .A1(n_234), .A2(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_238), .A2(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
OR2x2_ASAP7_75t_L g369 ( .A(n_241), .B(n_257), .Y(n_369) );
AND2x2_ASAP7_75t_L g507 ( .A(n_241), .B(n_451), .Y(n_507) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g389 ( .A(n_242), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_242), .B(n_331), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_242), .B(n_307), .Y(n_444) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
AND2x2_ASAP7_75t_L g317 ( .A(n_243), .B(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_SL g330 ( .A(n_243), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g338 ( .A(n_243), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_243), .B(n_307), .Y(n_409) );
AND2x2_ASAP7_75t_L g457 ( .A(n_243), .B(n_286), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_243), .B(n_285), .Y(n_500) );
BUFx2_ASAP7_75t_L g519 ( .A(n_243), .Y(n_519) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_255), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_250), .Y(n_268) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g303 ( .A(n_257), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g416 ( .A(n_257), .Y(n_416) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_274), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_258), .B(n_286), .Y(n_319) );
INVx2_ASAP7_75t_L g331 ( .A(n_258), .Y(n_331) );
AND2x2_ASAP7_75t_L g367 ( .A(n_258), .B(n_275), .Y(n_367) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AOI21x1_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_273), .Y(n_259) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_260), .A2(n_287), .A3(n_293), .B(n_295), .Y(n_286) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_260), .A2(n_549), .A3(n_594), .B(n_597), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_268), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g292 ( .A(n_266), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_SL g618 ( .A(n_272), .Y(n_618) );
INVx1_ASAP7_75t_L g391 ( .A(n_274), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_274), .B(n_286), .Y(n_408) );
INVx2_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
OR2x2_ASAP7_75t_L g350 ( .A(n_275), .B(n_286), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_275), .B(n_286), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_303), .B1(n_305), .B2(n_309), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_297), .B1(n_301), .B2(n_302), .Y(n_283) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_284), .B(n_367), .Y(n_381) );
AND2x2_ASAP7_75t_L g415 ( .A(n_284), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g333 ( .A(n_286), .Y(n_333) );
INVx1_ASAP7_75t_L g339 ( .A(n_286), .Y(n_339) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_293), .A2(n_615), .A3(n_616), .B(n_620), .Y(n_614) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_SL g611 ( .A(n_294), .Y(n_611) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g473 ( .A(n_299), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
AND3x1_ASAP7_75t_L g458 ( .A(n_300), .B(n_321), .C(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g414 ( .A(n_301), .Y(n_414) );
AND2x4_ASAP7_75t_L g450 ( .A(n_301), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g488 ( .A(n_304), .Y(n_488) );
INVx1_ASAP7_75t_L g492 ( .A(n_305), .Y(n_492) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
OR2x2_ASAP7_75t_L g465 ( .A(n_306), .B(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_306), .Y(n_513) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g413 ( .A(n_307), .B(n_391), .Y(n_413) );
AND2x2_ASAP7_75t_L g455 ( .A(n_307), .B(n_322), .Y(n_455) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_307), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_310), .A2(n_311), .B(n_375), .C(n_381), .Y(n_374) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_310), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_310), .B(n_468), .Y(n_514) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_312), .B(n_341), .Y(n_360) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_315), .B(n_320), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx2_ASAP7_75t_L g336 ( .A(n_318), .Y(n_336) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_319), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_320), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_321), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_321), .B(n_387), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_321), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_321), .B(n_379), .Y(n_535) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g518 ( .A(n_322), .Y(n_518) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g344 ( .A(n_325), .Y(n_344) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_340), .B(n_345), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
OAI33xp33_ASAP7_75t_L g394 ( .A1(n_330), .A2(n_335), .A3(n_395), .B1(n_396), .B2(n_398), .B3(n_399), .Y(n_394) );
OR2x2_ASAP7_75t_L g526 ( .A(n_330), .B(n_350), .Y(n_526) );
INVx2_ASAP7_75t_L g528 ( .A(n_330), .Y(n_528) );
INVx1_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
OR2x2_ASAP7_75t_L g390 ( .A(n_331), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g398 ( .A(n_335), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_335), .B(n_517), .C(n_519), .Y(n_516) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_336), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_336), .B(n_500), .Y(n_504) );
AND2x4_ASAP7_75t_L g533 ( .A(n_336), .B(n_534), .Y(n_533) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
OR2x2_ASAP7_75t_L g365 ( .A(n_338), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g478 ( .A(n_338), .B(n_413), .Y(n_478) );
INVx1_ASAP7_75t_L g534 ( .A(n_338), .Y(n_534) );
AND2x4_ASAP7_75t_SL g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
INVx1_ASAP7_75t_L g400 ( .A(n_342), .Y(n_400) );
AND2x2_ASAP7_75t_L g441 ( .A(n_342), .B(n_344), .Y(n_441) );
INVx1_ASAP7_75t_L g481 ( .A(n_343), .Y(n_481) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g372 ( .A(n_344), .B(n_373), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_351), .B1(n_358), .B2(n_360), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
INVx2_ASAP7_75t_L g451 ( .A(n_350), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_355), .C(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g395 ( .A(n_352), .Y(n_395) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_353), .B(n_378), .Y(n_480) );
OR2x2_ASAP7_75t_L g496 ( .A(n_353), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g509 ( .A(n_353), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_355), .B(n_423), .Y(n_484) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_382), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_368), .B2(n_370), .C(n_374), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI32xp33_ASAP7_75t_L g531 ( .A1(n_365), .A2(n_462), .A3(n_480), .B1(n_532), .B2(n_535), .Y(n_531) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g501 ( .A(n_367), .Y(n_501) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_370), .A2(n_383), .B(n_388), .Y(n_382) );
NAND2x1_ASAP7_75t_L g530 ( .A(n_371), .B(n_518), .Y(n_530) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
AND2x2_ASAP7_75t_L g524 ( .A(n_377), .B(n_405), .Y(n_524) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g472 ( .A(n_378), .Y(n_472) );
INVx2_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g401 ( .A(n_385), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_410), .C(n_421), .D(n_432), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_401), .B1(n_403), .B2(n_406), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_395), .A2(n_523), .B1(n_525), .B2(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g505 ( .A(n_400), .B(n_464), .Y(n_505) );
AND2x2_ASAP7_75t_L g508 ( .A(n_402), .B(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_403), .A2(n_422), .B1(n_426), .B2(n_429), .Y(n_421) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
OR2x2_ASAP7_75t_L g443 ( .A(n_408), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g427 ( .A(n_409), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_415), .B(n_417), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_411), .A2(n_516), .B(n_520), .C(n_522), .Y(n_515) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
AND2x4_ASAP7_75t_L g483 ( .A(n_416), .B(n_457), .Y(n_483) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_423), .A2(n_449), .B(n_452), .Y(n_448) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g454 ( .A(n_424), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_424), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g430 ( .A(n_428), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_430), .A2(n_461), .B1(n_465), .B2(n_467), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_439), .B2(n_442), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_437), .Y(n_453) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_510), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_469), .C(n_485), .D(n_502), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g512 ( .A(n_450), .B(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_456), .B2(n_458), .Y(n_452) );
INVxp67_ASAP7_75t_L g476 ( .A(n_456), .Y(n_476) );
BUFx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g466 ( .A(n_457), .Y(n_466) );
AND2x2_ASAP7_75t_L g489 ( .A(n_457), .B(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_475), .B(n_477), .Y(n_469) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x6_ASAP7_75t_L g494 ( .A(n_472), .B(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g491 ( .A(n_473), .Y(n_491) );
OAI32xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .A3(n_481), .B1(n_482), .B2(n_484), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B1(n_491), .B2(n_492), .C(n_493), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_499), .Y(n_493) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g525 ( .A(n_504), .Y(n_525) );
INVx1_ASAP7_75t_L g521 ( .A(n_505), .Y(n_521) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OAI211xp5_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_514), .B(n_515), .C(n_527), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVxp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_531), .Y(n_527) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
BUFx8_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g871 ( .A(n_538), .B(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g863 ( .A(n_539), .Y(n_863) );
XNOR2x1_ASAP7_75t_L g885 ( .A(n_540), .B(n_886), .Y(n_885) );
AND3x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_723), .C(n_777), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_683), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_622), .C(n_665), .Y(n_542) );
OAI21xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_565), .B(n_580), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g715 ( .A(n_546), .B(n_626), .Y(n_715) );
INVx2_ASAP7_75t_L g741 ( .A(n_546), .Y(n_741) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_558), .Y(n_546) );
INVx1_ASAP7_75t_L g640 ( .A(n_547), .Y(n_640) );
INVx2_ASAP7_75t_L g755 ( .A(n_547), .Y(n_755) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g568 ( .A(n_548), .Y(n_568) );
AND2x4_ASAP7_75t_L g698 ( .A(n_548), .B(n_660), .Y(n_698) );
INVx1_ASAP7_75t_L g751 ( .A(n_558), .Y(n_751) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g579 ( .A(n_559), .Y(n_579) );
AND2x4_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_559), .Y(n_657) );
INVx2_ASAP7_75t_L g660 ( .A(n_559), .Y(n_660) );
OR2x2_ASAP7_75t_L g674 ( .A(n_559), .B(n_631), .Y(n_674) );
AND2x2_ASAP7_75t_L g776 ( .A(n_559), .B(n_570), .Y(n_776) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g831 ( .A(n_566), .B(n_832), .Y(n_831) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
OR2x2_ASAP7_75t_L g658 ( .A(n_567), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_567), .B(n_677), .Y(n_722) );
AND2x2_ASAP7_75t_L g787 ( .A(n_567), .B(n_763), .Y(n_787) );
INVx4_ASAP7_75t_L g821 ( .A(n_567), .Y(n_821) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g656 ( .A(n_568), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g694 ( .A(n_568), .B(n_628), .Y(n_694) );
AND2x2_ASAP7_75t_L g804 ( .A(n_568), .B(n_631), .Y(n_804) );
AND2x2_ASAP7_75t_L g838 ( .A(n_568), .B(n_660), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_579), .Y(n_569) );
INVx4_ASAP7_75t_SL g628 ( .A(n_570), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_570), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g739 ( .A(n_570), .B(n_631), .Y(n_739) );
BUFx2_ASAP7_75t_L g757 ( .A(n_570), .Y(n_757) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_579), .A2(n_666), .B1(n_671), .B2(n_672), .C1(n_675), .C2(n_679), .Y(n_665) );
INVx1_ASAP7_75t_L g796 ( .A(n_579), .Y(n_796) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_591), .Y(n_580) );
AND2x2_ASAP7_75t_L g833 ( .A(n_581), .B(n_645), .Y(n_833) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g854 ( .A(n_582), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g663 ( .A(n_583), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_583), .B(n_646), .Y(n_802) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_584), .B(n_650), .Y(n_692) );
AND2x2_ASAP7_75t_L g720 ( .A(n_584), .B(n_600), .Y(n_720) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g649 ( .A(n_585), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g682 ( .A(n_585), .B(n_614), .Y(n_682) );
INVx1_ASAP7_75t_L g710 ( .A(n_585), .Y(n_710) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_585), .Y(n_816) );
AOI222xp33_ASAP7_75t_L g765 ( .A1(n_591), .A2(n_708), .B1(n_766), .B2(n_767), .C1(n_769), .C2(n_771), .Y(n_765) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_599), .Y(n_591) );
INVx1_ASAP7_75t_L g700 ( .A(n_592), .Y(n_700) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g646 ( .A(n_593), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_593), .B(n_614), .Y(n_651) );
AND2x2_ASAP7_75t_L g711 ( .A(n_593), .B(n_613), .Y(n_711) );
AND2x2_ASAP7_75t_L g699 ( .A(n_599), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g794 ( .A(n_599), .B(n_710), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_599), .B(n_801), .Y(n_800) );
AND3x1_ASAP7_75t_L g859 ( .A(n_599), .B(n_629), .C(n_860), .Y(n_859) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_613), .Y(n_599) );
AND2x2_ASAP7_75t_L g680 ( .A(n_600), .B(n_646), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_600), .B(n_782), .Y(n_829) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g643 ( .A(n_601), .Y(n_643) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_612), .Y(n_601) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_602), .A2(n_603), .B(n_612), .Y(n_650) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_611), .Y(n_603) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g645 ( .A(n_614), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g678 ( .A(n_614), .B(n_664), .Y(n_678) );
INVx1_ASAP7_75t_L g688 ( .A(n_614), .Y(n_688) );
BUFx2_ASAP7_75t_L g782 ( .A(n_614), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_641), .B(n_647), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_625), .B(n_638), .Y(n_624) );
AOI221xp5_ASAP7_75t_SL g705 ( .A1(n_625), .A2(n_706), .B1(n_712), .B2(n_716), .C(n_721), .Y(n_705) );
AND2x4_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_627), .B(n_640), .Y(n_826) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_628), .B(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g668 ( .A(n_628), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g704 ( .A(n_628), .Y(n_704) );
INVx1_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
AND2x2_ASAP7_75t_L g733 ( .A(n_628), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g745 ( .A(n_628), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_628), .B(n_751), .Y(n_858) );
INVx2_ASAP7_75t_L g693 ( .A(n_629), .Y(n_693) );
AND2x2_ASAP7_75t_L g703 ( .A(n_629), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_629), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_629), .B(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g654 ( .A(n_631), .Y(n_654) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_631), .Y(n_697) );
INVx1_ASAP7_75t_L g734 ( .A(n_631), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_631), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g673 ( .A(n_639), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_639), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_640), .Y(n_732) );
NOR2xp33_ASAP7_75t_R g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_643), .B(n_713), .C(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g744 ( .A(n_643), .B(n_651), .Y(n_744) );
AND2x2_ASAP7_75t_L g773 ( .A(n_643), .B(n_743), .Y(n_773) );
OR2x2_ASAP7_75t_L g840 ( .A(n_643), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g766 ( .A(n_645), .B(n_649), .Y(n_766) );
INVx2_ASAP7_75t_SL g850 ( .A(n_645), .Y(n_850) );
INVx2_ASAP7_75t_L g677 ( .A(n_646), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_646), .B(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g719 ( .A(n_646), .Y(n_719) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_646), .Y(n_792) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_652), .A3(n_655), .B1(n_658), .B2(n_661), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g671 ( .A(n_649), .B(n_651), .Y(n_671) );
AND2x2_ASAP7_75t_L g729 ( .A(n_649), .B(n_711), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_649), .B(n_711), .Y(n_737) );
INVx1_ASAP7_75t_L g664 ( .A(n_650), .Y(n_664) );
AND2x4_ASAP7_75t_SL g662 ( .A(n_651), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g806 ( .A(n_651), .Y(n_806) );
INVx2_ASAP7_75t_L g841 ( .A(n_651), .Y(n_841) );
AND2x2_ASAP7_75t_L g853 ( .A(n_651), .B(n_720), .Y(n_853) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_652), .B(n_774), .C(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g669 ( .A(n_654), .Y(n_669) );
AOI321xp33_ASAP7_75t_L g852 ( .A1(n_655), .A2(n_714), .A3(n_853), .B1(n_854), .B2(n_856), .C(n_859), .Y(n_852) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g670 ( .A(n_657), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_659), .A2(n_678), .B1(n_857), .B2(n_858), .Y(n_856) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g759 ( .A(n_663), .B(n_718), .Y(n_759) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g793 ( .A(n_668), .Y(n_793) );
NAND2x1_ASAP7_75t_L g820 ( .A(n_668), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_668), .B(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g818 ( .A(n_670), .B(n_804), .Y(n_818) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g758 ( .A(n_674), .Y(n_758) );
OR2x2_ASAP7_75t_L g825 ( .A(n_674), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_677), .B(n_678), .Y(n_702) );
NOR2x1p5_ASAP7_75t_L g743 ( .A(n_677), .B(n_682), .Y(n_743) );
INVx1_ASAP7_75t_L g813 ( .A(n_677), .Y(n_813) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_678), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_680), .Y(n_857) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_695), .C(n_705), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_693), .C(n_694), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g835 ( .A(n_689), .Y(n_835) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g727 ( .A(n_692), .Y(n_727) );
INVx1_ASAP7_75t_L g763 ( .A(n_692), .Y(n_763) );
NAND2xp33_ASAP7_75t_L g767 ( .A(n_693), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g771 ( .A(n_693), .Y(n_771) );
INVx1_ASAP7_75t_L g797 ( .A(n_694), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_699), .B(n_701), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx3_ASAP7_75t_L g746 ( .A(n_698), .Y(n_746) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g823 ( .A(n_710), .B(n_813), .Y(n_823) );
AND2x2_ASAP7_75t_L g726 ( .A(n_711), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g791 ( .A(n_711), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
OR2x2_ASAP7_75t_L g749 ( .A(n_714), .B(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g728 ( .A(n_715), .Y(n_728) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g762 ( .A(n_719), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g851 ( .A(n_720), .Y(n_851) );
NOR2xp67_ASAP7_75t_L g723 ( .A(n_724), .B(n_760), .Y(n_723) );
NAND3xp33_ASAP7_75t_SL g724 ( .A(n_725), .B(n_735), .C(n_747), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g768 ( .A(n_733), .Y(n_768) );
AND2x2_ASAP7_75t_L g843 ( .A(n_733), .B(n_754), .Y(n_843) );
INVx1_ASAP7_75t_L g790 ( .A(n_734), .Y(n_790) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI32xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .A3(n_740), .B1(n_742), .B2(n_745), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g770 ( .A(n_739), .Y(n_770) );
NAND2x1_ASAP7_75t_L g808 ( .A(n_739), .B(n_809), .Y(n_808) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g769 ( .A(n_741), .B(n_770), .Y(n_769) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OAI211xp5_ASAP7_75t_SL g795 ( .A1(n_746), .A2(n_789), .B(n_796), .C(n_797), .Y(n_795) );
INVx2_ASAP7_75t_L g809 ( .A(n_746), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_752), .B(n_759), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_753), .Y(n_764) );
NAND2x1_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx2_ASAP7_75t_L g847 ( .A(n_754), .Y(n_847) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g855 ( .A(n_755), .B(n_790), .Y(n_855) );
AND2x2_ASAP7_75t_L g860 ( .A(n_755), .B(n_816), .Y(n_860) );
AND2x4_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g785 ( .A(n_758), .Y(n_785) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .B(n_765), .C(n_772), .Y(n_760) );
INVxp67_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_762), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_810), .C(n_839), .Y(n_777) );
OAI211xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_783), .B(n_786), .C(n_798), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_784), .A2(n_823), .B1(n_824), .B2(n_827), .Y(n_822) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_794), .B2(n_795), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_791), .B1(n_792), .B2(n_793), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_789), .B(n_821), .Y(n_832) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g803 ( .A(n_796), .B(n_804), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_803), .B1(n_805), .B2(n_807), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OR2x2_ASAP7_75t_L g828 ( .A(n_802), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI211xp5_ASAP7_75t_SL g810 ( .A1(n_811), .A2(n_817), .B(n_822), .C(n_830), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_833), .B1(n_834), .B2(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OAI211xp5_ASAP7_75t_SL g839 ( .A1(n_840), .A2(n_842), .B(n_844), .C(n_852), .Y(n_839) );
INVxp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OR2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVx4_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx5_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
BUFx10_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
CKINVDCx16_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
AOI211xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_881), .B(n_889), .C(n_890), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
XNOR2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .Y(n_881) );
NOR2xp67_ASAP7_75t_SL g890 ( .A(n_891), .B(n_892), .Y(n_890) );
endmodule