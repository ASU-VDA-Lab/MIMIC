module fake_jpeg_12302_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_49),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_51),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_52),
.B1(n_56),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_58),
.B1(n_50),
.B2(n_21),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_51),
.Y(n_87)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_45),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_46),
.B(n_1),
.C(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_73),
.C(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_13),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_22),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_91),
.C(n_96),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_9),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_23),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_98),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_25),
.B(n_37),
.C(n_36),
.Y(n_96)
);

AOI22x1_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_11),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_26),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.C(n_40),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_27),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_31),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_119),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.C(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_105),
.B(n_113),
.C(n_112),
.D(n_110),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_127),
.C(n_116),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_119),
.C(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_128),
.B(n_122),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_118),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_101),
.Y(n_137)
);


endmodule