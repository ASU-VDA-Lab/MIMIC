module real_jpeg_25383_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_38),
.B(n_54),
.C(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_23),
.C(n_26),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_18),
.B1(n_19),
.B2(n_55),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_41),
.B(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_23),
.B1(n_28),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_23),
.B1(n_28),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_46),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_42),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_78),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_77),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_51),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_15),
.B(n_51),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.C(n_40),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_16),
.A2(n_34),
.B1(n_35),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_29),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_18),
.A2(n_19),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_18),
.A2(n_39),
.B(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_84),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_55),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_28),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_30),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_32),
.B(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_40),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_50),
.Y(n_63)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_63),
.B(n_92),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_64),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_63),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_106),
.B(n_111),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_94),
.B(n_105),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_90),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_101),
.B(n_104),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_110),
.Y(n_111)
);


endmodule