module fake_jpeg_25297_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_24),
.Y(n_65)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_27),
.B1(n_22),
.B2(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_73),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_27),
.B1(n_46),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_82),
.B1(n_57),
.B2(n_47),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_77),
.B1(n_28),
.B2(n_18),
.Y(n_132)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_76),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_86),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_41),
.B(n_26),
.C(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_17),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_17),
.B1(n_16),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_95),
.B1(n_21),
.B2(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_19),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_21),
.B1(n_32),
.B2(n_16),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_98),
.B1(n_57),
.B2(n_28),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_19),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_22),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_34),
.CI(n_18),
.CON(n_130),
.SN(n_130)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_72),
.B1(n_77),
.B2(n_82),
.Y(n_135)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_121),
.Y(n_140)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_103),
.B(n_94),
.Y(n_138)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_75),
.B(n_70),
.C(n_89),
.Y(n_136)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_45),
.B1(n_34),
.B2(n_18),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_88),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_164),
.B1(n_124),
.B2(n_131),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_148),
.B(n_133),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_75),
.B1(n_68),
.B2(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_68),
.B(n_91),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_149),
.B(n_151),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_130),
.B1(n_132),
.B2(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_98),
.B1(n_97),
.B2(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_147),
.B(n_157),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_89),
.B(n_79),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_123),
.B(n_129),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_69),
.B1(n_98),
.B2(n_74),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_159),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_104),
.B(n_87),
.C(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_96),
.B1(n_90),
.B2(n_76),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_83),
.B1(n_37),
.B2(n_43),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_38),
.B(n_28),
.C(n_13),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_39),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_39),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_110),
.C(n_43),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_159),
.C(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_169),
.B(n_180),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_173),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_110),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_178),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_106),
.B1(n_121),
.B2(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_148),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_112),
.B(n_126),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_179),
.A2(n_183),
.B(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_189),
.B(n_4),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_149),
.B(n_137),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_116),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_190),
.C(n_198),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_133),
.B1(n_114),
.B2(n_112),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_4),
.B(n_5),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_160),
.B(n_141),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_114),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_146),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_199),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_34),
.B1(n_18),
.B2(n_25),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_135),
.A2(n_34),
.B1(n_31),
.B2(n_25),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_145),
.B1(n_162),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_158),
.B1(n_156),
.B2(n_31),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_156),
.B1(n_25),
.B2(n_20),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_20),
.C(n_15),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_213),
.C(n_198),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_223),
.B1(n_181),
.B2(n_180),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_4),
.B(n_5),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_212),
.B(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_14),
.C(n_13),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_191),
.B(n_185),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_220),
.B(n_224),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_6),
.B(n_7),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_6),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_225),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_179),
.A2(n_178),
.B(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_8),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_234),
.B1(n_207),
.B2(n_209),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_176),
.B1(n_185),
.B2(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_233),
.A2(n_244),
.B1(n_249),
.B2(n_201),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_197),
.B1(n_171),
.B2(n_188),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_177),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_237),
.B(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_240),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_167),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_246),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_217),
.B(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_228),
.B1(n_223),
.B2(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_206),
.B(n_172),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_254),
.CI(n_214),
.CON(n_266),
.SN(n_266)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_229),
.B1(n_224),
.B2(n_218),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_211),
.A2(n_171),
.B(n_187),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_235),
.B(n_249),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_196),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_168),
.C(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_225),
.C(n_210),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_213),
.B(n_200),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_268),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_260),
.B1(n_269),
.B2(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_202),
.B1(n_212),
.B2(n_215),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_267),
.C(n_241),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_239),
.C(n_247),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_272),
.B1(n_231),
.B2(n_230),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_233),
.A2(n_209),
.B1(n_203),
.B2(n_227),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_8),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_250),
.B1(n_235),
.B2(n_252),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_236),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_9),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_279),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_265),
.Y(n_294)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_282),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_267),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_253),
.C(n_232),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_292),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_230),
.B1(n_214),
.B2(n_10),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_289),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_8),
.CI(n_9),
.CON(n_286),
.SN(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_8),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_9),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_266),
.C(n_264),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_286),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_276),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_307),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_273),
.B1(n_274),
.B2(n_257),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_305),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_275),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_277),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_279),
.A2(n_256),
.B(n_260),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_308),
.B(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_290),
.B1(n_287),
.B2(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_259),
.C(n_280),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_317),
.C(n_304),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_290),
.C(n_258),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_300),
.B1(n_307),
.B2(n_299),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_324),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_293),
.B(n_300),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_312),
.B(n_315),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_308),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_303),
.B1(n_295),
.B2(n_11),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_330),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_316),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_318),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_322),
.B(n_326),
.C(n_331),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_325),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_321),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_319),
.B(n_10),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_10),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);


endmodule