module fake_aes_8533_n_436 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_436);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_436;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_134;
wire n_429;
wire n_233;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_103), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_76), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_58), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_37), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_50), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_75), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_73), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_89), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_106), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_74), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_57), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_54), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_104), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_55), .Y(n_134) );
INVxp67_ASAP7_75t_SL g135 ( .A(n_92), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_13), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_35), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_35), .Y(n_138) );
INVxp67_ASAP7_75t_SL g139 ( .A(n_102), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_66), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_4), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_67), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_15), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_90), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_70), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g148 ( .A(n_25), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_60), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_65), .Y(n_150) );
CKINVDCx14_ASAP7_75t_R g151 ( .A(n_42), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_17), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_77), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_12), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_72), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_31), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_34), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_79), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_107), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_68), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_23), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_38), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_85), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_53), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_43), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_155), .A2(n_45), .B(n_44), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_153), .B(n_46), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_108), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_150), .B(n_0), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_108), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_151), .B(n_0), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_109), .B(n_116), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_116), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_117), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_165), .B(n_1), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_117), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_120), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_148), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_120), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
XOR2xp5_ASAP7_75t_L g191 ( .A(n_141), .B(n_2), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_122), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_123), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_123), .B(n_5), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_174), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_195), .Y(n_197) );
NAND3xp33_ASAP7_75t_L g198 ( .A(n_171), .B(n_126), .C(n_124), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_195), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_177), .Y(n_201) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_179), .B(n_164), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_188), .A2(n_127), .B1(n_128), .B2(n_126), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_195), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_175), .B(n_164), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_179), .B(n_167), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_182), .B(n_110), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_175), .B(n_136), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_184), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_170), .B(n_127), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_174), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_188), .A2(n_129), .B1(n_130), .B2(n_128), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_180), .B(n_130), .C(n_129), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_184), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_180), .B(n_111), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_181), .B(n_131), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_181), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_181), .B(n_131), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_114), .B1(n_115), .B2(n_110), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_199), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_205), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_213), .A2(n_183), .B1(n_170), .B2(n_185), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_214), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_218), .B(n_191), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_214), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_208), .A2(n_172), .B(n_188), .C(n_186), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_202), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_214), .Y(n_234) );
INVx5_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_203), .B(n_189), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_204), .B(n_172), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_201), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_197), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_213), .A2(n_192), .B1(n_193), .B2(n_190), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_223), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_202), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_204), .A2(n_194), .B1(n_115), .B2(n_119), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_210), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_214), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
BUFx4f_ASAP7_75t_SL g248 ( .A(n_222), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_207), .B(n_113), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_207), .B(n_169), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_221), .B(n_118), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_220), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_228), .A2(n_204), .B1(n_217), .B2(n_215), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_229), .B(n_215), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_198), .B(n_219), .C(n_209), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_232), .A2(n_222), .B(n_224), .C(n_206), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_238), .B(n_225), .C(n_219), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_233), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_233), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_254), .A2(n_204), .B1(n_217), .B2(n_225), .Y(n_265) );
BUFx12f_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_229), .Y(n_267) );
OR2x6_ASAP7_75t_L g268 ( .A(n_237), .B(n_217), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_233), .B(n_211), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_240), .A2(n_144), .B1(n_163), .B2(n_154), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_231), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_231), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_231), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
INVx5_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_227), .Y(n_276) );
OR2x6_ASAP7_75t_L g277 ( .A(n_243), .B(n_241), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_242), .A2(n_200), .B(n_196), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_112), .B(n_139), .C(n_135), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_248), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_242), .A2(n_200), .B(n_196), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_121), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_239), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_245), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_245), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_244), .A2(n_132), .B1(n_146), .B2(n_125), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_249), .B(n_243), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_251), .Y(n_289) );
INVx8_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_290), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_280), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_284), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_290), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_284), .Y(n_295) );
AOI22xp33_ASAP7_75t_SL g296 ( .A1(n_270), .A2(n_247), .B1(n_246), .B2(n_159), .Y(n_296) );
NAND2x1_ASAP7_75t_L g297 ( .A(n_259), .B(n_252), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_290), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_275), .B(n_247), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_268), .A2(n_247), .B1(n_256), .B2(n_255), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_265), .A2(n_256), .B1(n_157), .B2(n_187), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_257), .A2(n_157), .B1(n_187), .B2(n_152), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
CKINVDCx6p67_ASAP7_75t_R g304 ( .A(n_266), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_289), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_262), .A2(n_157), .B1(n_161), .B2(n_137), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_258), .A2(n_134), .B(n_133), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_277), .B(n_138), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_275), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_279), .B(n_145), .C(n_143), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_278), .A2(n_200), .B(n_196), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_283), .A2(n_140), .B1(n_147), .B2(n_142), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_286), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_287), .A2(n_166), .B(n_168), .C(n_162), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_282), .B(n_6), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_276), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_281), .A2(n_200), .B(n_196), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_261), .A2(n_264), .B(n_263), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_263), .B(n_160), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_269), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_260), .A2(n_173), .B(n_176), .C(n_178), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_309), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_308), .A2(n_273), .B1(n_271), .B2(n_267), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_313), .A2(n_288), .B1(n_274), .B2(n_272), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_304), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_318), .A2(n_212), .B(n_216), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_216), .B1(n_9), .B2(n_10), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_8), .B1(n_11), .B2(n_12), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_315), .A2(n_216), .B1(n_14), .B2(n_16), .Y(n_331) );
AO31x2_ASAP7_75t_L g332 ( .A1(n_314), .A2(n_18), .A3(n_19), .B(n_20), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_321), .A2(n_19), .B(n_21), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_319), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_299), .A2(n_317), .B(n_311), .Y(n_338) );
OAI221xp5_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_26), .B1(n_27), .B2(n_28), .C(n_29), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_291), .B(n_30), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_296), .A2(n_32), .B1(n_33), .B2(n_36), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_307), .A2(n_297), .B(n_305), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_320), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_298), .B(n_39), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_310), .A2(n_40), .B(n_41), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_325), .B(n_309), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_324), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_344), .B(n_316), .Y(n_350) );
NOR2xp33_ASAP7_75t_R g351 ( .A(n_326), .B(n_292), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_322), .B(n_309), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_343), .Y(n_353) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_338), .A2(n_306), .B(n_312), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_322), .B(n_294), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_339), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_51), .B(n_52), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_340), .A2(n_59), .B1(n_61), .B2(n_63), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_334), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_336), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_323), .B(n_69), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_332), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_78), .B(n_80), .C(n_81), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_330), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_327), .A2(n_333), .B(n_345), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_330), .A2(n_97), .B1(n_98), .B2(n_100), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_341), .A2(n_329), .B(n_337), .C(n_335), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_347), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_366), .B(n_342), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_356), .B(n_360), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_360), .B(n_361), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_346), .B(n_349), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_348), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_367), .A2(n_369), .B1(n_353), .B2(n_370), .C(n_350), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_362), .B(n_358), .Y(n_379) );
NAND4xp25_ASAP7_75t_SL g380 ( .A(n_359), .B(n_364), .C(n_351), .D(n_357), .Y(n_380) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_354), .B(n_358), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_368), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_368), .B(n_363), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_363), .B(n_365), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_363), .B(n_365), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_363), .A2(n_366), .B(n_365), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_365), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_365), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_348), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_363), .B(n_365), .Y(n_392) );
AO21x2_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_366), .B(n_365), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_373), .B(n_374), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_379), .Y(n_396) );
OR2x6_ASAP7_75t_L g397 ( .A(n_379), .B(n_375), .Y(n_397) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_371), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_386), .B(n_387), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_386), .B(n_387), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_389), .B(n_392), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_378), .Y(n_402) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_380), .B(n_377), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_389), .B(n_392), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_390), .B(n_385), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_388), .B(n_393), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_382), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_393), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_372), .B(n_383), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_403), .A2(n_384), .B(n_381), .Y(n_411) );
AND2x4_ASAP7_75t_SL g412 ( .A(n_402), .B(n_400), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_399), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_409), .B(n_376), .C(n_391), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_406), .B(n_401), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_406), .B(n_401), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_404), .B(n_394), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_415), .B(n_410), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_417), .B(n_410), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_413), .B(n_407), .Y(n_420) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_411), .A2(n_396), .B1(n_397), .B2(n_408), .C(n_405), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_417), .B(n_405), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_416), .B(n_398), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_412), .B(n_395), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_418), .B(n_420), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_424), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_426), .A2(n_421), .B1(n_423), .B2(n_424), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_427), .A2(n_425), .B1(n_419), .B2(n_422), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_428), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_429), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_430), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_430), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_431), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_432), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_433), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_435), .A2(n_434), .B1(n_433), .B2(n_414), .Y(n_436) );
endmodule