module fake_netlist_5_597_n_967 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_967);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_967;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_947;
wire n_757;
wire n_820;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_964;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_928;
wire n_858;
wire n_829;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_781;
wire n_711;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_893;
wire n_502;
wire n_892;
wire n_736;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_18),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_35),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_112),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_27),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_41),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_61),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_10),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_14),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_7),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_102),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_7),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_163),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_33),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_88),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_108),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_101),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_157),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

CKINVDCx6p67_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_3),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_37),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_81),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_63),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_133),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_96),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_19),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_10),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_119),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_15),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_124),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_5),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_71),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_87),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_171),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_212),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_261),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_212),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_227),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_194),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_195),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_247),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_200),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_208),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_223),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_196),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_1),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_214),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_197),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_198),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_216),
.B(n_1),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_231),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_199),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_202),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_221),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_192),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_219),
.B(n_2),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_224),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_256),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_204),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_276),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_244),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_296),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_299),
.B(n_222),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_226),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_305),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_279),
.A2(n_268),
.B1(n_273),
.B2(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_232),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_277),
.B(n_226),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_306),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_308),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_311),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_316),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_248),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_297),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_268),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_R g365 ( 
.A(n_272),
.B(n_230),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_266),
.B(n_253),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_284),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_303),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_286),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_298),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_368),
.B(n_253),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_216),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_340),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_250),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_255),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_257),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_234),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_329),
.Y(n_388)
);

OR2x6_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_258),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_265),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_339),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_365),
.Y(n_393)
);

OAI22x1_ASAP7_75t_L g394 ( 
.A1(n_319),
.A2(n_271),
.B1(n_269),
.B2(n_311),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_263),
.B1(n_260),
.B2(n_240),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_240),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_226),
.B1(n_230),
.B2(n_264),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_321),
.B(n_205),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_206),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

BUFx8_ASAP7_75t_SL g417 ( 
.A(n_336),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_374),
.B(n_207),
.Y(n_420)
);

NAND2x1p5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_215),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_218),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_337),
.B(n_220),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_331),
.B(n_229),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_345),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_357),
.B(n_26),
.Y(n_431)
);

CKINVDCx8_ASAP7_75t_R g432 ( 
.A(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_323),
.B(n_236),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_373),
.B(n_242),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_323),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_243),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_333),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_322),
.B(n_245),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_325),
.B(n_246),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_364),
.B(n_269),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_320),
.B(n_2),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_325),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_328),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_328),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_362),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_332),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_332),
.Y(n_453)
);

AND2x6_ASAP7_75t_SL g454 ( 
.A(n_444),
.B(n_271),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_386),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_445),
.A2(n_371),
.B1(n_249),
.B2(n_251),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_396),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_439),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_390),
.B(n_341),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_371),
.B1(n_252),
.B2(n_262),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_341),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_383),
.B(n_362),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_411),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_382),
.A2(n_347),
.B1(n_343),
.B2(n_342),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_382),
.B(n_347),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_382),
.B(n_385),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_336),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_423),
.B(n_342),
.Y(n_477)
);

O2A1O1Ixp5_ASAP7_75t_L g478 ( 
.A1(n_377),
.A2(n_93),
.B(n_189),
.C(n_187),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_450),
.A2(n_343),
.B1(n_4),
.B2(n_5),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_387),
.B(n_3),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_6),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_379),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_408),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_382),
.B(n_29),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

BUFx6f_ASAP7_75t_SL g488 ( 
.A(n_444),
.Y(n_488)
);

O2A1O1Ixp5_ASAP7_75t_L g489 ( 
.A1(n_377),
.A2(n_97),
.B(n_184),
.C(n_183),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_382),
.B(n_30),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_385),
.B(n_31),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_429),
.B(n_32),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_380),
.B(n_8),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_34),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_408),
.B(n_9),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_389),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_428),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_424),
.B(n_11),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_443),
.B(n_434),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_403),
.B(n_11),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_395),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_442),
.Y(n_505)
);

NAND2x1_ASAP7_75t_L g506 ( 
.A(n_381),
.B(n_36),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_434),
.B(n_15),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_421),
.B(n_16),
.Y(n_508)
);

BUFx8_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_418),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_17),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_421),
.B(n_18),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_383),
.B(n_19),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_428),
.B(n_20),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_395),
.B(n_21),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_441),
.B(n_21),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_409),
.B(n_39),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_40),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_186),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_413),
.B(n_42),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_448),
.B(n_181),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_43),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_397),
.Y(n_527)
);

AND2x4_ASAP7_75t_SL g528 ( 
.A(n_446),
.B(n_44),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_451),
.B(n_22),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_433),
.B(n_45),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_437),
.B(n_22),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_435),
.B(n_23),
.Y(n_532)
);

BUFx5_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_46),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_407),
.B(n_47),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_505),
.A2(n_449),
.B1(n_451),
.B2(n_446),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_393),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_509),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_407),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_462),
.B(n_407),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_468),
.B(n_393),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_474),
.A2(n_381),
.B(n_384),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_473),
.B(n_388),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_483),
.B(n_407),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_502),
.A2(n_384),
.B(n_414),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_519),
.A2(n_414),
.B(n_426),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_452),
.B(n_442),
.Y(n_550)
);

OAI21xp33_ASAP7_75t_L g551 ( 
.A1(n_496),
.A2(n_383),
.B(n_389),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_494),
.B(n_422),
.Y(n_552)
);

O2A1O1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_517),
.A2(n_422),
.B(n_447),
.C(n_399),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_459),
.B(n_407),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_459),
.B(n_511),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_520),
.A2(n_426),
.B(n_438),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_532),
.A2(n_444),
.B(n_431),
.C(n_394),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_458),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_522),
.A2(n_438),
.B(n_427),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_431),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_526),
.A2(n_427),
.B(n_425),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_497),
.B(n_431),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_465),
.B(n_431),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_530),
.A2(n_534),
.B(n_491),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_480),
.B(n_416),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_485),
.A2(n_425),
.B(n_416),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_485),
.A2(n_425),
.B(n_416),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_500),
.B(n_425),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_456),
.A2(n_432),
.B1(n_48),
.B2(n_51),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_457),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_461),
.B(n_24),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_535),
.A2(n_115),
.B(n_52),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_464),
.B(n_24),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_466),
.B(n_56),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_500),
.A2(n_57),
.B(n_58),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_527),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_471),
.B(n_59),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_535),
.A2(n_60),
.B(n_62),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_518),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_453),
.B(n_417),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_478),
.A2(n_67),
.B(n_69),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_515),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_475),
.B(n_417),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_456),
.B(n_70),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_492),
.A2(n_72),
.B(n_73),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_503),
.A2(n_74),
.B(n_75),
.Y(n_590)
);

AOI21xp33_ASAP7_75t_L g591 ( 
.A1(n_477),
.A2(n_76),
.B(n_77),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_533),
.B(n_78),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_463),
.B(n_79),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_489),
.A2(n_80),
.B(n_83),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_487),
.Y(n_595)
);

AOI22x1_ASAP7_75t_SL g596 ( 
.A1(n_454),
.A2(n_84),
.B1(n_85),
.B2(n_90),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_512),
.B(n_91),
.Y(n_597)
);

NAND2x1p5_ASAP7_75t_L g598 ( 
.A(n_498),
.B(n_94),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_549),
.A2(n_506),
.B(n_495),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_543),
.A2(n_486),
.B(n_490),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_508),
.B(n_513),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_574),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_541),
.A2(n_521),
.B(n_524),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_560),
.A2(n_528),
.B(n_527),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_569),
.B(n_529),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_556),
.A2(n_514),
.B(n_523),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_597),
.A2(n_527),
.B(n_510),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_554),
.A2(n_484),
.B(n_501),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_550),
.A2(n_463),
.B1(n_531),
.B2(n_529),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_583),
.A2(n_594),
.B(n_588),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_559),
.A2(n_499),
.B(n_516),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_584),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_585),
.Y(n_614)
);

AO21x1_ASAP7_75t_L g615 ( 
.A1(n_590),
.A2(n_484),
.B(n_504),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_542),
.B(n_504),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_576),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_469),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_507),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_563),
.A2(n_533),
.B(n_472),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_551),
.A2(n_557),
.B(n_553),
.C(n_590),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_593),
.A2(n_479),
.B(n_533),
.C(n_454),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_547),
.B(n_479),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_561),
.A2(n_533),
.B(n_99),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_572),
.A2(n_533),
.B(n_488),
.C(n_509),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

AO21x1_ASAP7_75t_L g629 ( 
.A1(n_591),
.A2(n_98),
.B(n_100),
.Y(n_629)
);

NOR2x1_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_488),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_555),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_106),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_540),
.A2(n_107),
.B(n_109),
.C(n_110),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_537),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_558),
.Y(n_635)
);

AO31x2_ASAP7_75t_L g636 ( 
.A1(n_571),
.A2(n_111),
.A3(n_113),
.B(n_114),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_573),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_116),
.B(n_117),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_536),
.B(n_120),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_552),
.A2(n_123),
.B(n_125),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_548),
.A2(n_126),
.B(n_127),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_575),
.B(n_579),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_581),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_581),
.A2(n_132),
.B(n_136),
.C(n_137),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_578),
.A2(n_138),
.B(n_139),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_546),
.A2(n_140),
.B(n_141),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_578),
.B(n_143),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_544),
.B(n_538),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_562),
.A2(n_566),
.B(n_567),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_562),
.A2(n_144),
.B(n_146),
.C(n_148),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_538),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_628),
.B(n_587),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_613),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_624),
.B(n_582),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_616),
.B(n_598),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_638),
.B(n_539),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_638),
.B(n_580),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_610),
.A2(n_568),
.B1(n_589),
.B2(n_577),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_618),
.B(n_596),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

BUFx2_ASAP7_75t_SL g662 ( 
.A(n_635),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_611),
.A2(n_149),
.B(n_150),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_637),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_602),
.Y(n_665)
);

BUFx2_ASAP7_75t_R g666 ( 
.A(n_649),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_606),
.A2(n_622),
.B(n_623),
.C(n_611),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_614),
.Y(n_668)
);

O2A1O1Ixp5_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_626),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_605),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_SL g672 ( 
.A1(n_644),
.A2(n_156),
.B(n_158),
.C(n_159),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_619),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_620),
.A2(n_166),
.B(n_167),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_634),
.B(n_168),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_630),
.B(n_169),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_621),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_605),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_621),
.B(n_170),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_606),
.B(n_176),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_607),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_644),
.A2(n_632),
.B1(n_640),
.B2(n_601),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_612),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_632),
.A2(n_173),
.B1(n_175),
.B2(n_629),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_652),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_605),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_651),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_627),
.B(n_643),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_648),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_643),
.B(n_604),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_631),
.B(n_648),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_603),
.A2(n_650),
.B(n_600),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_636),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_646),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_608),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_636),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_639),
.A2(n_641),
.B1(n_647),
.B2(n_642),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_636),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_599),
.A2(n_611),
.B(n_603),
.Y(n_699)
);

NAND2x1p5_ASAP7_75t_L g700 ( 
.A(n_625),
.B(n_538),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_605),
.Y(n_701)
);

AOI222xp33_ASAP7_75t_L g702 ( 
.A1(n_616),
.A2(n_445),
.B1(n_496),
.B2(n_408),
.C1(n_606),
.C2(n_624),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_609),
.B(n_649),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_616),
.B(n_542),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_681),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_696),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_702),
.B(n_704),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_702),
.A2(n_655),
.B1(n_687),
.B2(n_691),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_687),
.A2(n_691),
.B1(n_688),
.B2(n_660),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_703),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_683),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_667),
.A2(n_682),
.B(n_690),
.Y(n_712)
);

AOI21x1_ASAP7_75t_L g713 ( 
.A1(n_699),
.A2(n_692),
.B(n_698),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_677),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_700),
.A2(n_694),
.B(n_674),
.Y(n_716)
);

AOI21x1_ASAP7_75t_L g717 ( 
.A1(n_698),
.A2(n_690),
.B(n_659),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_671),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_671),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_658),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_656),
.A2(n_703),
.B1(n_653),
.B2(n_689),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_700),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_703),
.B(n_661),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_SL g724 ( 
.A1(n_695),
.A2(n_677),
.B(n_673),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_677),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_687),
.A2(n_691),
.B1(n_680),
.B2(n_653),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_674),
.A2(n_697),
.B(n_659),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_664),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_679),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_671),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_668),
.B(n_670),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_666),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_665),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_693),
.Y(n_735)
);

CKINVDCx11_ASAP7_75t_R g736 ( 
.A(n_678),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_701),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_672),
.A2(n_663),
.B(n_669),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_691),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_657),
.A2(n_673),
.B1(n_684),
.B2(n_676),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_686),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_701),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_701),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_678),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_675),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_662),
.B(n_702),
.Y(n_747)
);

CKINVDCx11_ASAP7_75t_R g748 ( 
.A(n_654),
.Y(n_748)
);

AOI21x1_ASAP7_75t_L g749 ( 
.A1(n_699),
.A2(n_692),
.B(n_698),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_661),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_696),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_696),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_654),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_702),
.A2(n_606),
.B1(n_615),
.B2(n_518),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_702),
.B(n_704),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_704),
.A2(n_542),
.B(n_525),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_702),
.B(n_704),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_692),
.A2(n_625),
.B(n_699),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_681),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_696),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_704),
.A2(n_610),
.B1(n_408),
.B2(n_616),
.Y(n_762)
);

AO21x2_ASAP7_75t_L g763 ( 
.A1(n_699),
.A2(n_692),
.B(n_698),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_705),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_753),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_750),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_713),
.A2(n_749),
.B(n_717),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_746),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_706),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_720),
.B(n_747),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_746),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_747),
.B(n_707),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_723),
.Y(n_773)
);

AO21x2_ASAP7_75t_L g774 ( 
.A1(n_727),
.A2(n_712),
.B(n_717),
.Y(n_774)
);

BUFx12f_ASAP7_75t_L g775 ( 
.A(n_748),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_746),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_725),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_756),
.Y(n_778)
);

AO21x2_ASAP7_75t_L g779 ( 
.A1(n_759),
.A2(n_763),
.B(n_738),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_756),
.B(n_758),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_710),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_728),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_722),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_706),
.Y(n_784)
);

HB1xp67_ASAP7_75t_SL g785 ( 
.A(n_719),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_751),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_710),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_751),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_722),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_723),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_752),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_752),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_755),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_744),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_758),
.B(n_762),
.Y(n_795)
);

INVx3_ASAP7_75t_SL g796 ( 
.A(n_730),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_754),
.A2(n_757),
.B(n_724),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_739),
.B(n_725),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_739),
.B(n_725),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_739),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_738),
.A2(n_761),
.B(n_755),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_777),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_770),
.B(n_735),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_764),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_770),
.B(n_735),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_797),
.A2(n_709),
.B1(n_708),
.B2(n_740),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_773),
.B(n_763),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_778),
.B(n_721),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_773),
.B(n_763),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_802),
.B(n_714),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_775),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_778),
.B(n_728),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_769),
.Y(n_814)
);

AO21x2_ASAP7_75t_L g815 ( 
.A1(n_767),
.A2(n_724),
.B(n_716),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_769),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_802),
.B(n_714),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_784),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_777),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_784),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_764),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_790),
.B(n_760),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_795),
.B(n_781),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_800),
.B(n_761),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_800),
.B(n_714),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_786),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_772),
.B(n_728),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_786),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_777),
.B(n_711),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_781),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_788),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_788),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_777),
.B(n_711),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_791),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_791),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_792),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_764),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_807),
.A2(n_797),
.B1(n_795),
.B2(n_740),
.C(n_726),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_804),
.B(n_787),
.Y(n_839)
);

OAI221xp5_ASAP7_75t_L g840 ( 
.A1(n_809),
.A2(n_780),
.B1(n_715),
.B2(n_732),
.C(n_765),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_823),
.B(n_772),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_823),
.B(n_780),
.Y(n_842)
);

NAND4xp25_ASAP7_75t_L g843 ( 
.A(n_804),
.B(n_787),
.C(n_798),
.D(n_799),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_SL g844 ( 
.A1(n_806),
.A2(n_775),
.B1(n_729),
.B2(n_774),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_806),
.B(n_777),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_813),
.B(n_766),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_827),
.B(n_768),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_830),
.B(n_802),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_814),
.B(n_798),
.C(n_799),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_811),
.B(n_771),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_824),
.B(n_776),
.Y(n_851)
);

AOI221xp5_ASAP7_75t_L g852 ( 
.A1(n_808),
.A2(n_794),
.B1(n_731),
.B2(n_734),
.C(n_733),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_824),
.B(n_782),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_814),
.B(n_793),
.C(n_792),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_SL g855 ( 
.A1(n_808),
.A2(n_732),
.B(n_737),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_816),
.B(n_793),
.C(n_733),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_810),
.B(n_789),
.Y(n_857)
);

OA211x2_ASAP7_75t_L g858 ( 
.A1(n_812),
.A2(n_785),
.B(n_796),
.C(n_775),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_830),
.B(n_789),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_810),
.B(n_789),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_830),
.B(n_734),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_811),
.A2(n_737),
.B(n_718),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_811),
.A2(n_737),
.B(n_743),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_816),
.A2(n_774),
.B1(n_729),
.B2(n_731),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_825),
.B(n_789),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_857),
.B(n_822),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_860),
.B(n_822),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_845),
.B(n_865),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_842),
.B(n_841),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_839),
.B(n_803),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_852),
.B(n_826),
.C(n_828),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_859),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_854),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_851),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_842),
.B(n_828),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_862),
.B(n_803),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_856),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_849),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_853),
.B(n_803),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_846),
.B(n_803),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_863),
.B(n_817),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_850),
.B(n_825),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_847),
.Y(n_884)
);

NAND2x1p5_ASAP7_75t_L g885 ( 
.A(n_871),
.B(n_850),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_874),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_874),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_869),
.B(n_843),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_871),
.B(n_844),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_880),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_871),
.B(n_855),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_882),
.B(n_817),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_873),
.B(n_819),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_878),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_866),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_886),
.A2(n_838),
.B1(n_840),
.B2(n_872),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_888),
.B(n_895),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_887),
.B(n_879),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_890),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_891),
.B(n_889),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_895),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_890),
.B(n_879),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_885),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_893),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_893),
.Y(n_906)
);

INVx3_ASAP7_75t_SL g907 ( 
.A(n_897),
.Y(n_907)
);

INVx3_ASAP7_75t_SL g908 ( 
.A(n_901),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_905),
.B(n_891),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_906),
.B(n_889),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_903),
.B(n_884),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_911),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_907),
.B(n_896),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_910),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_907),
.B(n_896),
.Y(n_915)
);

OAI222xp33_ASAP7_75t_L g916 ( 
.A1(n_913),
.A2(n_899),
.B1(n_903),
.B2(n_909),
.C1(n_900),
.C2(n_904),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_914),
.B(n_908),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_912),
.B(n_898),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_915),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_913),
.B(n_902),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_919),
.B(n_885),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_917),
.B(n_892),
.Y(n_922)
);

XOR2x2_ASAP7_75t_L g923 ( 
.A(n_920),
.B(n_892),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_L g924 ( 
.A(n_918),
.B(n_916),
.C(n_736),
.Y(n_924)
);

AOI221xp5_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_876),
.B1(n_875),
.B2(n_864),
.C(n_877),
.Y(n_925)
);

OAI221xp5_ASAP7_75t_L g926 ( 
.A1(n_919),
.A2(n_873),
.B1(n_864),
.B2(n_883),
.C(n_861),
.Y(n_926)
);

AOI221xp5_ASAP7_75t_L g927 ( 
.A1(n_916),
.A2(n_877),
.B1(n_892),
.B2(n_861),
.C(n_882),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_919),
.B(n_873),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_L g929 ( 
.A(n_924),
.B(n_730),
.C(n_741),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_SL g930 ( 
.A(n_927),
.B(n_730),
.C(n_858),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_928),
.B(n_921),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_923),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_922),
.A2(n_877),
.B1(n_882),
.B2(n_881),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_926),
.Y(n_934)
);

NAND4xp25_ASAP7_75t_L g935 ( 
.A(n_931),
.B(n_925),
.C(n_719),
.D(n_730),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_SL g936 ( 
.A(n_929),
.B(n_742),
.C(n_741),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_932),
.B(n_870),
.Y(n_937)
);

NOR2x1p5_ASAP7_75t_L g938 ( 
.A(n_934),
.B(n_719),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_933),
.B(n_819),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_930),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_938),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_940),
.A2(n_870),
.B1(n_745),
.B2(n_811),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_935),
.A2(n_817),
.B1(n_774),
.B2(n_819),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_937),
.A2(n_796),
.B1(n_742),
.B2(n_745),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_939),
.A2(n_867),
.B1(n_819),
.B2(n_818),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_941),
.B(n_936),
.C(n_742),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_942),
.B(n_868),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_943),
.B(n_868),
.Y(n_948)
);

AND3x4_ASAP7_75t_L g949 ( 
.A(n_944),
.B(n_817),
.C(n_745),
.Y(n_949)
);

XOR2x2_ASAP7_75t_L g950 ( 
.A(n_946),
.B(n_945),
.Y(n_950)
);

XOR2xp5_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_801),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_949),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_947),
.B1(n_796),
.B2(n_819),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_950),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_SL g955 ( 
.A(n_954),
.B(n_951),
.C(n_836),
.Y(n_955)
);

NAND5xp2_ASAP7_75t_L g956 ( 
.A(n_953),
.B(n_801),
.C(n_836),
.D(n_831),
.E(n_835),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_955),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_957),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_959),
.A2(n_956),
.B(n_835),
.Y(n_960)
);

AOI32xp33_ASAP7_75t_L g961 ( 
.A1(n_958),
.A2(n_729),
.A3(n_834),
.B1(n_818),
.B2(n_820),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_960),
.A2(n_779),
.B(n_834),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_961),
.Y(n_963)
);

AOI322xp5_ASAP7_75t_L g964 ( 
.A1(n_963),
.A2(n_729),
.A3(n_831),
.B1(n_832),
.B2(n_826),
.C1(n_820),
.C2(n_829),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_962),
.A2(n_832),
.B1(n_815),
.B2(n_774),
.Y(n_965)
);

AOI221xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_783),
.B1(n_837),
.B2(n_821),
.C(n_805),
.Y(n_966)
);

AOI211xp5_ASAP7_75t_L g967 ( 
.A1(n_966),
.A2(n_964),
.B(n_829),
.C(n_833),
.Y(n_967)
);


endmodule