module fake_jpeg_14790_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_24),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_22),
.B1(n_30),
.B2(n_19),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_22),
.B1(n_30),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_63),
.B1(n_29),
.B2(n_21),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_62),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_0),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_20),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_27),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_27),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_18),
.B1(n_32),
.B2(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_20),
.Y(n_71)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_82),
.B1(n_80),
.B2(n_75),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_47),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_53),
.B1(n_56),
.B2(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_36),
.B(n_23),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_59),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_53),
.B1(n_29),
.B2(n_55),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_104),
.B1(n_113),
.B2(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_97),
.B1(n_77),
.B2(n_72),
.Y(n_127)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_99),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_25),
.C(n_60),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_52),
.B1(n_56),
.B2(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_112),
.B1(n_82),
.B2(n_65),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_83),
.B1(n_70),
.B2(n_66),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_64),
.B1(n_61),
.B2(n_49),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_111),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_31),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_25),
.B1(n_17),
.B2(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_25),
.B1(n_17),
.B2(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_123),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_131),
.B1(n_103),
.B2(n_25),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_78),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_93),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_137),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_132),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_72),
.B1(n_77),
.B2(n_83),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_100),
.B1(n_111),
.B2(n_96),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_81),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_81),
.B(n_86),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_100),
.C(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_132),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_69),
.C(n_88),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_1),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_69),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_157),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_144),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_166),
.B1(n_138),
.B2(n_129),
.Y(n_175)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_101),
.B1(n_112),
.B2(n_111),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_119),
.B(n_89),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_95),
.B1(n_106),
.B2(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_23),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_68),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_88),
.B1(n_23),
.B2(n_31),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_114),
.B(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_9),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_131),
.B1(n_122),
.B2(n_5),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_114),
.C(n_125),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_179),
.C(n_182),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_175),
.B(n_162),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_172),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_181),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_139),
.C(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_142),
.B1(n_153),
.B2(n_157),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_121),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_118),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_187),
.C(n_149),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_118),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_178),
.A2(n_166),
.B1(n_152),
.B2(n_153),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_198),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_173),
.B1(n_189),
.B2(n_175),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_190),
.B1(n_164),
.B2(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_148),
.B1(n_151),
.B2(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_148),
.B(n_143),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_140),
.B1(n_141),
.B2(n_119),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_179),
.C(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_169),
.C(n_158),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_213),
.C(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_199),
.C(n_209),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_225),
.B1(n_226),
.B2(n_194),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_161),
.C(n_141),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_89),
.C(n_1),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_197),
.B1(n_192),
.B2(n_212),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_231),
.C(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_198),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_208),
.B(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_205),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_202),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_208),
.B(n_196),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_192),
.B(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_222),
.B1(n_215),
.B2(n_216),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_237),
.B1(n_229),
.B2(n_230),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_7),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_8),
.B(n_10),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_237),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_248),
.B1(n_232),
.B2(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_5),
.C(n_6),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_7),
.C(n_8),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_252),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_255),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_231),
.B1(n_235),
.B2(n_9),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_241),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_8),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_262),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_242),
.A3(n_240),
.B1(n_247),
.B2(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_261),
.Y(n_264)
);

OAI221xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_246),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_251),
.C(n_250),
.Y(n_266)
);

AOI321xp33_ASAP7_75t_SL g267 ( 
.A1(n_264),
.A2(n_253),
.A3(n_255),
.B1(n_15),
.B2(n_12),
.C(n_13),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_12),
.B(n_15),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_268),
.C(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_15),
.Y(n_272)
);


endmodule