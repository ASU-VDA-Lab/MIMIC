module fake_jpeg_29524_n_517 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_55),
.Y(n_132)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_74),
.Y(n_169)
);

CKINVDCx9p33_ASAP7_75t_R g75 ( 
.A(n_17),
.Y(n_75)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_2),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_17),
.B(n_33),
.CON(n_78),
.SN(n_78)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_95),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_81),
.Y(n_121)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_21),
.B(n_5),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_17),
.B(n_6),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_21),
.B(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_24),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_107),
.B1(n_103),
.B2(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_120),
.A2(n_128),
.B1(n_137),
.B2(n_139),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_58),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_31),
.B1(n_49),
.B2(n_45),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_59),
.Y(n_130)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_60),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_133),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_31),
.B1(n_49),
.B2(n_45),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_78),
.B1(n_71),
.B2(n_54),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_35),
.B(n_38),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_146),
.A2(n_23),
.B1(n_53),
.B2(n_52),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_67),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_147),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_77),
.A2(n_28),
.B1(n_52),
.B2(n_50),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_23),
.B1(n_50),
.B2(n_53),
.Y(n_190)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_172),
.Y(n_252)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_176),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_102),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_179),
.Y(n_265)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_66),
.B1(n_79),
.B2(n_72),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_181),
.A2(n_221),
.B1(n_132),
.B2(n_121),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_42),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_187),
.Y(n_227)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_111),
.A2(n_79),
.A3(n_96),
.B1(n_44),
.B2(n_41),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_194),
.Y(n_230)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_190),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_82),
.B1(n_63),
.B2(n_65),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_210),
.B1(n_212),
.B2(n_121),
.Y(n_226)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_35),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_38),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_39),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_39),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_122),
.A2(n_26),
.B1(n_52),
.B2(n_50),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_74),
.B1(n_69),
.B2(n_91),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_80),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_83),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_207),
.Y(n_254)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_211),
.Y(n_259)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_168),
.A2(n_158),
.B1(n_146),
.B2(n_116),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_97),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_99),
.B1(n_93),
.B2(n_89),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_214),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_217),
.Y(n_262)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_129),
.B(n_96),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_223),
.B1(n_224),
.B2(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_135),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_131),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_129),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_115),
.Y(n_246)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_226),
.A2(n_249),
.B1(n_183),
.B2(n_209),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_237),
.A2(n_183),
.B1(n_28),
.B2(n_53),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_118),
.B1(n_133),
.B2(n_130),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_132),
.B1(n_202),
.B2(n_234),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_134),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_134),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_140),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_218),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_157),
.C(n_161),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_156),
.C(n_154),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_200),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_272),
.Y(n_302)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_274),
.A2(n_280),
.B(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_191),
.B1(n_204),
.B2(n_181),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_277),
.A2(n_279),
.B1(n_284),
.B2(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_187),
.B1(n_179),
.B2(n_189),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_202),
.B(n_212),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_238),
.A2(n_180),
.B1(n_221),
.B2(n_207),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_246),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_123),
.B1(n_124),
.B2(n_140),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_250),
.A2(n_123),
.B1(n_124),
.B2(n_169),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_213),
.B(n_29),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_259),
.B(n_254),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_292),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_226),
.A2(n_177),
.B1(n_216),
.B2(n_199),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_231),
.B1(n_252),
.B2(n_261),
.Y(n_331)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_262),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_244),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_297),
.B1(n_32),
.B2(n_29),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_253),
.B(n_22),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_295),
.B(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_34),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_256),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_263),
.B1(n_264),
.B2(n_240),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_265),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_243),
.A2(n_184),
.B1(n_34),
.B2(n_32),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_310),
.B1(n_331),
.B2(n_280),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

XOR2x1_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_227),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_322),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_307),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_309),
.A2(n_231),
.B(n_297),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_275),
.A2(n_227),
.B1(n_259),
.B2(n_254),
.Y(n_310)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_230),
.C(n_235),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_269),
.C(n_282),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_318),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_292),
.B(n_241),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_316),
.B(n_296),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_272),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_317),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_230),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_241),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_277),
.B1(n_285),
.B2(n_295),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_326),
.A2(n_289),
.B1(n_281),
.B2(n_268),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_287),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_327),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_286),
.A2(n_235),
.B1(n_265),
.B2(n_251),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_333),
.C(n_337),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_279),
.C(n_273),
.Y(n_337)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_312),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_287),
.B(n_274),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_354),
.B(n_328),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_318),
.B(n_288),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_344),
.B(n_345),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_316),
.B(n_252),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_284),
.B1(n_298),
.B2(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_352),
.Y(n_368)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_304),
.B1(n_310),
.B2(n_305),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_355),
.B1(n_356),
.B2(n_303),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_327),
.A2(n_289),
.B(n_278),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_326),
.A2(n_308),
.B1(n_301),
.B2(n_314),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_308),
.A2(n_299),
.B1(n_283),
.B2(n_291),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_297),
.B1(n_290),
.B2(n_271),
.Y(n_357)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_243),
.B1(n_242),
.B2(n_255),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_358),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_302),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_359),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_361),
.B(n_309),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_335),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_380),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_311),
.B(n_360),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_379),
.B1(n_384),
.B2(n_387),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_321),
.C(n_329),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_381),
.C(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_329),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_339),
.A2(n_360),
.B(n_352),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_303),
.C(n_306),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_306),
.B1(n_323),
.B2(n_307),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_356),
.B1(n_359),
.B2(n_340),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_323),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_347),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_335),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_348),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_354),
.B1(n_342),
.B2(n_343),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_368),
.B1(n_319),
.B2(n_317),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_364),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_396),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_385),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_338),
.B(n_347),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_418),
.B(n_365),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_383),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_377),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_399),
.B(n_402),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_401),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_361),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_391),
.B(n_350),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_350),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_403),
.A2(n_408),
.B1(n_414),
.B2(n_376),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_371),
.A2(n_346),
.B1(n_357),
.B2(n_354),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_406),
.A2(n_369),
.B1(n_362),
.B2(n_387),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_363),
.Y(n_408)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_312),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_413),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_302),
.Y(n_413)
);

A2O1A1O1Ixp25_ASAP7_75t_L g418 ( 
.A1(n_379),
.A2(n_343),
.B(n_313),
.C(n_348),
.D(n_320),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_381),
.C(n_374),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_423),
.C(n_425),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_380),
.B(n_370),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_427),
.B(n_423),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_422),
.A2(n_440),
.B1(n_416),
.B2(n_415),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_384),
.C(n_372),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_424),
.A2(n_404),
.B1(n_231),
.B2(n_247),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_413),
.C(n_392),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_388),
.C(n_368),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_426),
.B(n_428),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_394),
.C(n_412),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_431),
.Y(n_443)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_430),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_375),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_417),
.A2(n_365),
.B1(n_373),
.B2(n_315),
.Y(n_433)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_320),
.C(n_325),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_407),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_330),
.B1(n_242),
.B2(n_255),
.Y(n_438)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_393),
.A2(n_330),
.B1(n_255),
.B2(n_258),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_405),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_243),
.B1(n_236),
.B2(n_247),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_418),
.Y(n_444)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_421),
.A2(n_409),
.B(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_434),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_447),
.B(n_453),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_451),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_422),
.A2(n_415),
.B1(n_407),
.B2(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_452),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_428),
.A2(n_404),
.B1(n_410),
.B2(n_236),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_435),
.Y(n_454)
);

OAI321xp33_ASAP7_75t_L g463 ( 
.A1(n_454),
.A2(n_432),
.A3(n_228),
.B1(n_229),
.B2(n_245),
.C(n_261),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_426),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_431),
.A2(n_429),
.B1(n_440),
.B2(n_436),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_458),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_419),
.C(n_425),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_461),
.C(n_473),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_432),
.C(n_420),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_437),
.B(n_420),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_236),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_468),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_457),
.A2(n_232),
.B1(n_261),
.B2(n_229),
.Y(n_465)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_465),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_232),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_229),
.B1(n_228),
.B2(n_192),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_470),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_455),
.A2(n_229),
.B1(n_228),
.B2(n_192),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_229),
.C(n_8),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_472),
.C(n_471),
.Y(n_496)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_478),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_459),
.B(n_456),
.CI(n_443),
.CON(n_479),
.SN(n_479)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_443),
.C(n_448),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_484),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_450),
.C(n_452),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_444),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_475),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_467),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_487),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_466),
.B(n_7),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_7),
.C(n_8),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_8),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_476),
.Y(n_503)
);

BUFx12f_ASAP7_75t_SL g492 ( 
.A(n_479),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_492),
.A2(n_494),
.B(n_480),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_477),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_498),
.Y(n_500)
);

OAI321xp33_ASAP7_75t_L g494 ( 
.A1(n_482),
.A2(n_471),
.A3(n_466),
.B1(n_472),
.B2(n_473),
.C(n_12),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_56),
.C(n_9),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_490),
.B(n_495),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_491),
.B(n_484),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_502),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_476),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_505),
.C(n_8),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_481),
.B1(n_485),
.B2(n_483),
.C(n_488),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_L g509 ( 
.A1(n_504),
.A2(n_9),
.B(n_10),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_506),
.A2(n_509),
.B(n_500),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_10),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_511),
.C(n_508),
.Y(n_512)
);

AOI322xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_16),
.C2(n_509),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_11),
.B(n_12),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_11),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_12),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_13),
.C(n_366),
.Y(n_517)
);


endmodule