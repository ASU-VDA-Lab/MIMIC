module fake_netlist_1_401_n_835 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_835);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_835;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_58), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_33), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_48), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_80), .Y(n_106) );
BUFx2_ASAP7_75t_SL g107 ( .A(n_18), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_84), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_52), .Y(n_109) );
OR2x2_ASAP7_75t_L g110 ( .A(n_50), .B(n_42), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_37), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_11), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_62), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_45), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_31), .Y(n_119) );
NOR2xp67_ASAP7_75t_L g120 ( .A(n_4), .B(n_22), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_85), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_46), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_36), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_4), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_19), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_32), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_43), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_53), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_23), .B(n_49), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_88), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_38), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_8), .Y(n_136) );
BUFx10_ASAP7_75t_L g137 ( .A(n_9), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_56), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_115), .B(n_0), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_105), .B(n_0), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
CKINVDCx8_ASAP7_75t_R g145 ( .A(n_119), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_112), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_108), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_113), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_114), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_114), .B(n_1), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
BUFx12f_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_110), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_116), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_125), .B(n_3), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
BUFx8_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_145), .A2(n_125), .B1(n_109), .B2(n_111), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_161), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_161), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_142), .B(n_117), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_124), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_146), .B(n_102), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_146), .B(n_102), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_148), .B(n_131), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_162), .B(n_104), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_162), .B(n_104), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_162), .B(n_106), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_148), .A2(n_107), .B1(n_132), .B2(n_138), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_157), .B(n_137), .Y(n_188) );
NAND2xp33_ASAP7_75t_R g189 ( .A(n_150), .B(n_106), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_157), .B(n_120), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_154), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_137), .B1(n_129), .B2(n_128), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_152), .B(n_127), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_160), .B(n_127), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_158), .B(n_128), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_155), .B(n_129), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_145), .B(n_133), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_153), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_155), .B(n_126), .Y(n_202) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_141), .B(n_133), .C(n_134), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_197), .B(n_153), .Y(n_206) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_184), .B(n_134), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_197), .B(n_153), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_203), .B(n_140), .Y(n_209) );
NOR2xp67_ASAP7_75t_L g210 ( .A(n_185), .B(n_20), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_188), .B(n_121), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_188), .B(n_123), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_184), .B(n_135), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_164), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_185), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_195), .B(n_135), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_181), .A2(n_149), .B1(n_130), .B2(n_147), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_192), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_198), .A2(n_159), .B(n_147), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_172), .B(n_21), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_194), .B(n_143), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
NOR2xp67_ASAP7_75t_L g228 ( .A(n_174), .B(n_24), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_190), .B(n_5), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_199), .B(n_61), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_181), .A2(n_159), .B1(n_147), .B2(n_144), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_181), .B(n_5), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_193), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_181), .A2(n_147), .B1(n_144), .B2(n_143), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_163), .B(n_6), .C(n_7), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_170), .B(n_159), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_171), .B(n_159), .Y(n_241) );
INVx8_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_193), .B(n_6), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_182), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_196), .B(n_159), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_182), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_166), .B(n_147), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_200), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_169), .B(n_144), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_176), .Y(n_252) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_173), .A2(n_144), .B1(n_143), .B2(n_10), .C(n_11), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_177), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_206), .B(n_175), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_178), .B(n_179), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_207), .B(n_248), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_221), .A2(n_178), .B(n_180), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_248), .B(n_190), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_211), .B(n_190), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_213), .B(n_177), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_219), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_225), .A2(n_178), .B(n_202), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_225), .A2(n_178), .B(n_204), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_234), .A2(n_204), .B(n_205), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_207), .B(n_200), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_219), .B(n_7), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_209), .B(n_8), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_208), .B(n_10), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_207), .B(n_12), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_252), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_216), .A2(n_205), .B(n_201), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_233), .A2(n_201), .B(n_191), .C(n_187), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_222), .A2(n_191), .B(n_187), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_231), .B(n_144), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_214), .B(n_12), .Y(n_280) );
INVx11_ASAP7_75t_L g281 ( .A(n_214), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_243), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_229), .B(n_13), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
NOR2xp33_ASAP7_75t_R g285 ( .A(n_249), .B(n_13), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_242), .B(n_14), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_251), .B(n_14), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_216), .A2(n_183), .B(n_186), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_242), .B(n_15), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_242), .B(n_15), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_242), .B(n_16), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_214), .B(n_16), .Y(n_293) );
BUFx10_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_282), .A2(n_231), .B(n_235), .C(n_233), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_265), .A2(n_241), .B(n_226), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_277), .A2(n_210), .B(n_228), .Y(n_297) );
AOI211x1_ASAP7_75t_L g298 ( .A1(n_270), .A2(n_243), .B(n_251), .C(n_250), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_264), .A2(n_245), .B(n_240), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_269), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_279), .A2(n_220), .B(n_210), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_280), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_281), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_288), .A2(n_228), .B(n_224), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_284), .A2(n_224), .B(n_229), .Y(n_309) );
O2A1O1Ixp5_ASAP7_75t_L g310 ( .A1(n_278), .A2(n_230), .B(n_247), .C(n_229), .Y(n_310) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_255), .A2(n_232), .B(n_249), .Y(n_311) );
AO32x2_ASAP7_75t_L g312 ( .A1(n_292), .A2(n_238), .A3(n_253), .B1(n_217), .B2(n_227), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_256), .A2(n_246), .B(n_244), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_258), .A2(n_246), .B(n_244), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_285), .B(n_227), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_275), .A2(n_239), .B(n_237), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
AO32x2_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_227), .A3(n_17), .B1(n_18), .B2(n_239), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_236), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_300), .B(n_262), .Y(n_320) );
OAI21x1_ASAP7_75t_SL g321 ( .A1(n_309), .A2(n_272), .B(n_268), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_309), .A2(n_257), .B(n_274), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_297), .A2(n_287), .B(n_266), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_295), .A2(n_261), .B(n_260), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_319), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_302), .B(n_283), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
AO31x2_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_286), .A3(n_291), .B(n_290), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_297), .A2(n_271), .B(n_276), .Y(n_333) );
HB1xp67_ASAP7_75t_SL g334 ( .A(n_307), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_317), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_301), .A2(n_273), .B(n_276), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_301), .A2(n_263), .B(n_259), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_303), .B(n_262), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_293), .B(n_255), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_319), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_303), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_298), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_308), .A2(n_236), .B(n_212), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_329), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_325), .B(n_318), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_339), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_325), .B(n_294), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_327), .B(n_318), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_327), .B(n_318), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_326), .A2(n_310), .B(n_299), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_343), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_346), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_342), .B(n_304), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_343), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_344), .Y(n_361) );
INVx4_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_328), .B(n_307), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_344), .B(n_294), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_321), .A2(n_316), .B(n_314), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_339), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_339), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_326), .B(n_294), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_333), .A2(n_316), .B(n_313), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_335), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_328), .B(n_267), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_332), .B(n_294), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_320), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_320), .Y(n_389) );
INVxp33_ASAP7_75t_L g390 ( .A(n_334), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_340), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_357), .B(n_328), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_353), .B(n_338), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_357), .B(n_331), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_385), .B(n_332), .Y(n_395) );
OR2x6_ASAP7_75t_L g396 ( .A(n_385), .B(n_340), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_332), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_360), .B(n_332), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_376), .A2(n_321), .B(n_315), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_348), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_356), .A2(n_337), .B(n_333), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_360), .B(n_332), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_353), .B(n_338), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_347), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_348), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_361), .B(n_332), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_347), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_354), .B(n_338), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_349), .B(n_387), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_354), .B(n_338), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_376), .A2(n_285), .B1(n_291), .B2(n_290), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_349), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_356), .A2(n_337), .B(n_322), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_351), .Y(n_415) );
OR2x2_ASAP7_75t_SL g416 ( .A(n_352), .B(n_338), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_370), .B(n_340), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_379), .A2(n_289), .B1(n_286), .B2(n_311), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_370), .B(n_318), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_361), .B(n_332), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_349), .B(n_342), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_382), .B(n_318), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_371), .B(n_289), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_364), .B(n_334), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_351), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_355), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_351), .B(n_342), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_368), .A2(n_333), .B(n_345), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_363), .B(n_312), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_363), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_362), .B(n_304), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_367), .B(n_312), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_358), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_367), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_367), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_350), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_390), .A2(n_322), .B1(n_273), .B2(n_304), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_350), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_372), .B(n_312), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_366), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_366), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_372), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_373), .B(n_17), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_373), .B(n_312), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_349), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_373), .B(n_324), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_374), .B(n_312), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_374), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_378), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_378), .B(n_324), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_378), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_380), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_380), .B(n_324), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_358), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_362), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_380), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_383), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_383), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_383), .B(n_345), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_365), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_365), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_381), .B(n_345), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_400), .B(n_391), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_460), .B(n_391), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_436), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_404), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_439), .B(n_387), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_400), .B(n_381), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_405), .B(n_362), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_424), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_405), .B(n_362), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_394), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_397), .B(n_389), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_393), .B(n_389), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_410), .B(n_349), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_442), .B(n_388), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_393), .B(n_388), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_403), .B(n_368), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_459), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_465), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_403), .B(n_368), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_409), .B(n_368), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_404), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_426), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_426), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_407), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_407), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_409), .B(n_349), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_408), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g500 ( .A(n_460), .B(n_359), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_397), .B(n_386), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_411), .B(n_386), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_423), .B(n_386), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_392), .B(n_398), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_408), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_415), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_411), .B(n_375), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_436), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_428), .B(n_375), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_402), .B(n_375), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_406), .B(n_369), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_395), .B(n_369), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_413), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_395), .B(n_369), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_420), .B(n_359), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_453), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_419), .B(n_359), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_454), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_419), .B(n_359), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_415), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_432), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_466), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_429), .B(n_377), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_454), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_410), .B(n_25), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_429), .B(n_377), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_422), .B(n_377), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_456), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_410), .B(n_377), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_456), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_432), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_467), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_467), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_422), .B(n_26), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_457), .B(n_27), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_433), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_417), .B(n_28), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_417), .B(n_29), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_461), .B(n_30), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_433), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g544 ( .A(n_450), .B(n_34), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_461), .B(n_35), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_431), .B(n_39), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_462), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_431), .B(n_41), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_435), .B(n_44), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_462), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_466), .B(n_47), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_435), .B(n_51), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_443), .B(n_54), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_418), .A2(n_237), .B1(n_212), .B2(n_223), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_446), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_463), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_447), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_437), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_443), .B(n_55), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_449), .B(n_57), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_437), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_438), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_438), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_441), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_449), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_448), .B(n_59), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_441), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_452), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_421), .B(n_60), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_471), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_500), .B(n_396), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_473), .Y(n_572) );
AND2x4_ASAP7_75t_SL g573 ( .A(n_509), .B(n_421), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_502), .B(n_396), .Y(n_574) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_509), .B(n_476), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_502), .B(n_396), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_475), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_396), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_508), .B(n_421), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_514), .B(n_455), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_471), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_516), .B(n_455), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_498), .B(n_451), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_498), .B(n_451), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_493), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_477), .Y(n_586) );
BUFx3_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_488), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_510), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_482), .B(n_448), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_488), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_527), .B(n_452), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_468), .B(n_458), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_470), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_469), .B(n_458), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_493), .Y(n_596) );
AND2x4_ASAP7_75t_SL g597 ( .A(n_479), .B(n_413), .Y(n_597) );
NOR2xp67_ASAP7_75t_L g598 ( .A(n_489), .B(n_450), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_482), .B(n_413), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_501), .B(n_464), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_531), .B(n_413), .Y(n_601) );
NOR2x1p5_ASAP7_75t_SL g602 ( .A(n_537), .B(n_416), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_486), .B(n_413), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_468), .B(n_414), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_544), .B(n_464), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_486), .B(n_440), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_517), .B(n_416), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_485), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_496), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_496), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_480), .B(n_401), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_474), .B(n_401), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_490), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_487), .B(n_401), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_497), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_487), .B(n_430), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_491), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_491), .B(n_430), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_533), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_555), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_492), .B(n_399), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_556), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_497), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_492), .B(n_430), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_499), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_539), .B(n_412), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_542), .B(n_434), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_499), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_494), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_527), .B(n_434), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_481), .B(n_63), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_495), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_512), .B(n_64), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_503), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_513), .B(n_66), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_67), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_518), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_505), .B(n_68), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_527), .B(n_69), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_520), .B(n_526), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_533), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_521), .B(n_70), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_530), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_506), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_534), .B(n_72), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_535), .B(n_73), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_524), .B(n_74), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_532), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_506), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_541), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_524), .B(n_75), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_547), .B(n_77), .Y(n_652) );
NOR2xp33_ASAP7_75t_SL g653 ( .A(n_478), .B(n_78), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_483), .B(n_79), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_478), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_507), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_483), .B(n_565), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_507), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_483), .B(n_82), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_550), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_522), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_504), .B(n_83), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_504), .B(n_89), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_564), .B(n_90), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_522), .Y(n_665) );
AOI21xp5_ASAP7_75t_SL g666 ( .A1(n_539), .A2(n_91), .B(n_92), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_564), .B(n_94), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_511), .B(n_95), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_472), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_529), .B(n_96), .Y(n_670) );
OAI32xp33_ASAP7_75t_L g671 ( .A1(n_655), .A2(n_545), .A3(n_540), .B1(n_551), .B2(n_569), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_611), .B(n_568), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_572), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_588), .Y(n_674) );
NAND2xp33_ASAP7_75t_SL g675 ( .A(n_594), .B(n_540), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_591), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_617), .B(n_528), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_626), .A2(n_557), .B1(n_484), .B2(n_554), .C(n_536), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_604), .B(n_563), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_619), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_608), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_613), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_589), .B(n_525), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_657), .B(n_562), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_620), .Y(n_686) );
BUFx3_ASAP7_75t_L g687 ( .A(n_587), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_622), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_626), .A2(n_553), .B1(n_548), .B2(n_549), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_640), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_669), .B(n_561), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_590), .B(n_538), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_640), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_630), .A2(n_554), .B1(n_559), .B2(n_546), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_587), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_604), .B(n_538), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_577), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_586), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_616), .B(n_523), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_641), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_616), .B(n_523), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_629), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_618), .B(n_543), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_632), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_593), .B(n_543), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_583), .B(n_567), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_618), .B(n_558), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_634), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_584), .B(n_579), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_637), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_624), .B(n_558), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_621), .B(n_612), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_643), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_648), .Y(n_714) );
AND2x4_ASAP7_75t_SL g715 ( .A(n_571), .B(n_560), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_574), .B(n_567), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_576), .B(n_515), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_624), .B(n_552), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_614), .B(n_552), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_593), .B(n_549), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_578), .B(n_515), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_580), .B(n_559), .Y(n_722) );
AOI22xp5_ASAP7_75t_SL g723 ( .A1(n_571), .A2(n_560), .B1(n_553), .B2(n_548), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_599), .B(n_515), .Y(n_724) );
NOR2xp67_ASAP7_75t_SL g725 ( .A(n_666), .B(n_546), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_614), .B(n_515), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_607), .B(n_566), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_650), .B(n_560), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_603), .B(n_97), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_602), .A2(n_183), .B(n_186), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_641), .Y(n_731) );
AND2x4_ASAP7_75t_L g732 ( .A(n_575), .B(n_98), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_582), .B(n_99), .Y(n_733) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_598), .B(n_100), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_660), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_575), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_595), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_600), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_570), .Y(n_739) );
INVx1_ASAP7_75t_SL g740 ( .A(n_573), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_606), .B(n_186), .Y(n_741) );
INVx2_ASAP7_75t_SL g742 ( .A(n_736), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_679), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_679), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_675), .A2(n_653), .B1(n_595), .B2(n_601), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_687), .B(n_627), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_689), .A2(n_630), .B1(n_592), .B2(n_639), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_696), .B(n_644), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_694), .A2(n_727), .B1(n_725), .B2(n_678), .Y(n_749) );
OR4x1_ASAP7_75t_L g750 ( .A(n_690), .B(n_573), .C(n_639), .D(n_597), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_737), .B(n_601), .Y(n_751) );
CKINVDCx14_ASAP7_75t_R g752 ( .A(n_683), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_680), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_684), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g755 ( .A(n_694), .B(n_663), .C(n_662), .D(n_638), .Y(n_755) );
AO22x1_ASAP7_75t_L g756 ( .A1(n_740), .A2(n_645), .B1(n_654), .B2(n_659), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_696), .B(n_644), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_700), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_726), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_693), .Y(n_760) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_715), .A2(n_592), .B(n_605), .Y(n_761) );
INVxp67_ASAP7_75t_L g762 ( .A(n_674), .Y(n_762) );
O2A1O1Ixp5_ASAP7_75t_SL g763 ( .A1(n_676), .A2(n_673), .B(n_681), .C(n_682), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_691), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_723), .A2(n_631), .B1(n_646), .B2(n_597), .Y(n_765) );
AOI222xp33_ASAP7_75t_L g766 ( .A1(n_719), .A2(n_638), .B1(n_605), .B2(n_636), .C1(n_642), .C2(n_670), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_719), .A2(n_601), .B1(n_635), .B2(n_633), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_686), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_718), .A2(n_670), .B1(n_668), .B2(n_625), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_677), .B(n_623), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_738), .B(n_651), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_730), .A2(n_647), .B1(n_664), .B2(n_667), .C(n_652), .Y(n_772) );
OAI21xp33_ASAP7_75t_L g773 ( .A1(n_712), .A2(n_610), .B(n_661), .Y(n_773) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_741), .A2(n_652), .B(n_665), .Y(n_774) );
NOR2xp67_ASAP7_75t_L g775 ( .A(n_734), .B(n_610), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_732), .A2(n_609), .B(n_661), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_706), .B(n_609), .Y(n_777) );
OR2x6_ASAP7_75t_L g778 ( .A(n_732), .B(n_596), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g779 ( .A1(n_695), .A2(n_596), .B1(n_658), .B2(n_656), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_731), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_688), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_756), .A2(n_671), .B(n_701), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_749), .A2(n_718), .B1(n_701), .B2(n_703), .C(n_707), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_761), .A2(n_707), .B(n_711), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_748), .B(n_705), .Y(n_785) );
INVx3_ASAP7_75t_L g786 ( .A(n_778), .Y(n_786) );
OAI211xp5_ASAP7_75t_L g787 ( .A1(n_752), .A2(n_745), .B(n_755), .C(n_766), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_764), .A2(n_697), .B1(n_735), .B2(n_710), .C(n_698), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_746), .A2(n_742), .B(n_767), .C(n_769), .Y(n_789) );
O2A1O1Ixp5_ASAP7_75t_L g790 ( .A1(n_747), .A2(n_702), .B(n_704), .C(n_708), .Y(n_790) );
OAI221xp5_ASAP7_75t_SL g791 ( .A1(n_778), .A2(n_722), .B1(n_720), .B2(n_733), .C(n_728), .Y(n_791) );
AOI322xp5_ASAP7_75t_L g792 ( .A1(n_771), .A2(n_709), .A3(n_692), .B1(n_685), .B2(n_714), .C1(n_713), .C2(n_716), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g793 ( .A1(n_773), .A2(n_672), .B(n_699), .Y(n_793) );
AOI21xp33_ASAP7_75t_SL g794 ( .A1(n_765), .A2(n_728), .B(n_726), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_743), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_751), .A2(n_717), .B1(n_721), .B2(n_724), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_744), .A2(n_729), .B1(n_711), .B2(n_703), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_763), .A2(n_699), .B(n_672), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_753), .B(n_739), .Y(n_799) );
AOI21xp33_ASAP7_75t_SL g800 ( .A1(n_778), .A2(n_615), .B(n_658), .Y(n_800) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_762), .A2(n_585), .B1(n_656), .B2(n_649), .C(n_628), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_775), .A2(n_585), .B1(n_649), .B2(n_628), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_760), .B(n_570), .Y(n_803) );
NAND2xp33_ASAP7_75t_L g804 ( .A(n_786), .B(n_750), .Y(n_804) );
NOR3xp33_ASAP7_75t_L g805 ( .A(n_787), .B(n_772), .C(n_758), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_789), .A2(n_754), .B1(n_768), .B2(n_781), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_786), .B(n_770), .Y(n_807) );
NAND4xp25_ASAP7_75t_L g808 ( .A(n_790), .B(n_775), .C(n_776), .D(n_774), .Y(n_808) );
NAND3xp33_ASAP7_75t_SL g809 ( .A(n_782), .B(n_780), .C(n_757), .Y(n_809) );
AOI211xp5_ASAP7_75t_L g810 ( .A1(n_794), .A2(n_779), .B(n_759), .C(n_777), .Y(n_810) );
OAI21xp33_ASAP7_75t_L g811 ( .A1(n_783), .A2(n_581), .B(n_625), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_799), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g813 ( .A1(n_791), .A2(n_665), .B(n_623), .C(n_615), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_784), .A2(n_581), .B(n_186), .Y(n_814) );
OAI211xp5_ASAP7_75t_L g815 ( .A1(n_805), .A2(n_792), .B(n_798), .C(n_800), .Y(n_815) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_809), .B(n_788), .C(n_801), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_804), .A2(n_793), .B(n_795), .Y(n_817) );
OAI22xp33_ASAP7_75t_SL g818 ( .A1(n_806), .A2(n_802), .B1(n_803), .B2(n_785), .Y(n_818) );
NAND4xp25_ASAP7_75t_L g819 ( .A(n_813), .B(n_797), .C(n_796), .D(n_803), .Y(n_819) );
NOR2xp33_ASAP7_75t_SL g820 ( .A(n_808), .B(n_186), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_815), .B(n_812), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_816), .B(n_811), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_819), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_823), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_822), .Y(n_825) );
NAND4xp75_ASAP7_75t_L g826 ( .A(n_825), .B(n_821), .C(n_817), .D(n_820), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_824), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_827), .Y(n_828) );
AO22x2_ASAP7_75t_L g829 ( .A1(n_826), .A2(n_818), .B1(n_814), .B2(n_807), .Y(n_829) );
NAND2x1p5_ASAP7_75t_L g830 ( .A(n_828), .B(n_810), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_830), .B(n_829), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_831), .A2(n_215), .B(n_218), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_832), .B(n_215), .Y(n_833) );
OR2x6_ASAP7_75t_L g834 ( .A(n_833), .B(n_218), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_834), .A2(n_223), .B1(n_227), .B2(n_825), .Y(n_835) );
endmodule