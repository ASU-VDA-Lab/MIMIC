module real_jpeg_23691_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_188;
wire n_139;
wire n_33;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_70),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_70),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_12),
.B1(n_85),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_95),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_95),
.Y(n_194)
);

INVx8_ASAP7_75t_SL g81 ( 
.A(n_5),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_87),
.B(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_6),
.B(n_78),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_26),
.C(n_27),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_68),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_6),
.A2(n_42),
.B1(n_188),
.B2(n_194),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_72),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_72),
.Y(n_178)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_115)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_116),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_53),
.B1(n_96),
.B2(n_97),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_22),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_24),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_24),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_24),
.B(n_91),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_25),
.B(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_32),
.B1(n_63),
.B2(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_31),
.B(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_32),
.A2(n_64),
.A3(n_66),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_32),
.B(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_56),
.B(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_36),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_36),
.A2(n_148),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_36),
.A2(n_147),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_36),
.A2(n_146),
.B1(n_147),
.B2(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_49),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_42),
.A2(n_49),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_42),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_42),
.A2(n_185),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_43),
.B(n_50),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_43),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_74),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_71),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_69),
.B1(n_73),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_68),
.B1(n_130),
.B2(n_139),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_66),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_80),
.B(n_90),
.C(n_111),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_65),
.B(n_91),
.CON(n_139),
.SN(n_139)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_79),
.C(n_92),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_86),
.B2(n_93),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_78),
.B1(n_94),
.B2(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_91),
.B(n_124),
.Y(n_199)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_122),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_117),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_120),
.B(n_122),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_209),
.B(n_213),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_162),
.B(n_208),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_149),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_136),
.B(n_149),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.C(n_145),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_137),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_145),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_157),
.C(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_203),
.B(n_207),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_181),
.B(n_202),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_169),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_190),
.B(n_201),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_189),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_200),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);


endmodule