module fake_jpeg_24473_n_305 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_19),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_34),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_25),
.B1(n_40),
.B2(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_26),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_29),
.C(n_31),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_76),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_31),
.B1(n_29),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_57),
.B1(n_54),
.B2(n_53),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_73),
.B(n_18),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_44),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_86),
.B1(n_28),
.B2(n_27),
.Y(n_119)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_19),
.B1(n_33),
.B2(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_51),
.B1(n_57),
.B2(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_107),
.B1(n_110),
.B2(n_114),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_97),
.Y(n_128)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_117),
.C(n_91),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_105),
.B(n_26),
.Y(n_149)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_49),
.B1(n_46),
.B2(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_118),
.Y(n_144)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_46),
.B1(n_54),
.B2(n_61),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_61),
.B1(n_45),
.B2(n_52),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_119),
.B1(n_81),
.B2(n_77),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_82),
.C(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_47),
.B(n_19),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_92),
.B(n_80),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_70),
.B1(n_82),
.B2(n_77),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_127),
.B1(n_142),
.B2(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_136),
.B(n_26),
.Y(n_176)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_75),
.B(n_94),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_139),
.C(n_147),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_86),
.B(n_84),
.C(n_42),
.D(n_43),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_143),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_61),
.B1(n_87),
.B2(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_74),
.B1(n_28),
.B2(n_27),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_43),
.B(n_42),
.C(n_26),
.D(n_17),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_78),
.B1(n_76),
.B2(n_28),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_120),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_106),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_112),
.B1(n_106),
.B2(n_109),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_152),
.B(n_157),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_175),
.B(n_177),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_115),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_136),
.C(n_142),
.Y(n_182)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_107),
.B1(n_95),
.B2(n_98),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_170),
.B1(n_180),
.B2(n_179),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_98),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_172),
.B(n_174),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_98),
.C(n_15),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_15),
.B(n_16),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_113),
.B1(n_97),
.B2(n_101),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_111),
.B(n_30),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_124),
.B(n_27),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_180),
.B(n_125),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_17),
.B(n_2),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_123),
.A2(n_97),
.B1(n_113),
.B2(n_85),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_85),
.B1(n_63),
.B2(n_3),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_185),
.C(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_147),
.C(n_139),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_140),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_192),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_126),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_199),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_175),
.B(n_164),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_133),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_63),
.B(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_150),
.C(n_130),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_134),
.C(n_132),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_133),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_203),
.C(n_177),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_179),
.B1(n_173),
.B2(n_171),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_43),
.C(n_42),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_162),
.C(n_158),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_178),
.B(n_17),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_170),
.B1(n_163),
.B2(n_161),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_212),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_172),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_225),
.C(n_230),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_165),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_194),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_166),
.B1(n_173),
.B2(n_155),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_223),
.B1(n_229),
.B2(n_187),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_152),
.B(n_168),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_227),
.B(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_183),
.B1(n_184),
.B2(n_202),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_226),
.C(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_192),
.B1(n_196),
.B2(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_228),
.Y(n_245)
);

OAI322xp33_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_168),
.A3(n_156),
.B1(n_151),
.B2(n_162),
.C1(n_16),
.C2(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_168),
.C(n_63),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_1),
.CI(n_2),
.CON(n_228),
.SN(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_16),
.B(n_14),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_188),
.B1(n_186),
.B2(n_198),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_246),
.B1(n_226),
.B2(n_214),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_204),
.B(n_195),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_241),
.B(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_243),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_228),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_184),
.B(n_205),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_209),
.C(n_213),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_259),
.C(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_260),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_209),
.C(n_213),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.C(n_263),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_211),
.C(n_217),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_210),
.C(n_228),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_4),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_13),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_4),
.Y(n_263)
);

OAI321xp33_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_237),
.A3(n_245),
.B1(n_235),
.B2(n_231),
.C(n_244),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_264),
.A2(n_235),
.B(n_233),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_259),
.B(n_258),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_240),
.B1(n_245),
.B2(n_242),
.C(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI31xp67_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_233),
.A3(n_246),
.B(n_242),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_232),
.C(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_6),
.C(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_254),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_275),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_232),
.B1(n_6),
.B2(n_7),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_5),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_263),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_10),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_286),
.B(n_269),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_10),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_9),
.C(n_10),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_12),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_8),
.B(n_9),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_274),
.C(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.C(n_294),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_269),
.B(n_274),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_279),
.B(n_278),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_299),
.C(n_295),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_287),
.A2(n_286),
.B(n_11),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_12),
.C(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_293),
.B(n_12),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_303),
.Y(n_305)
);


endmodule