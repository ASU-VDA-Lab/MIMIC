module fake_netlist_1_8245_n_1283 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1283);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1283;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_265;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_258;
wire n_253;
wire n_266;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_257;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_252;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_251;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_267;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_270;
wire n_1178;
wire n_259;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_260;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_264;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_255;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_256;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_262;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_263;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_261;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_119), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_32), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_219), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_46), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_128), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_126), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_149), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_27), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_94), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_196), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_67), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_144), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_171), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_220), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_58), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_165), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_20), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_17), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_8), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_34), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_92), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_24), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_24), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_123), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_13), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_206), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_84), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_217), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_193), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_117), .Y(n_284) );
BUFx10_ASAP7_75t_L g285 ( .A(n_155), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_139), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_191), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_98), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_109), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_117), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_166), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_135), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_33), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_197), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_225), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_26), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_8), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_62), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_158), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_224), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_141), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_242), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_29), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_138), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_56), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_207), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_66), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_40), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_3), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_151), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_198), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_143), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_77), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_244), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_98), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_162), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_202), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_161), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_215), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_212), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_209), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_28), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_194), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_250), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_164), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_116), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g328 ( .A(n_186), .B(n_190), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_66), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_175), .Y(n_330) );
BUFx10_ASAP7_75t_L g331 ( .A(n_181), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_14), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_142), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_44), .Y(n_334) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_243), .B(n_203), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_238), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_178), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_55), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_237), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_195), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_167), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_20), .Y(n_342) );
BUFx10_ASAP7_75t_L g343 ( .A(n_184), .Y(n_343) );
BUFx10_ASAP7_75t_L g344 ( .A(n_160), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_137), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_200), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_6), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_187), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_15), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_28), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_11), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_218), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_132), .Y(n_353) );
BUFx10_ASAP7_75t_L g354 ( .A(n_227), .Y(n_354) );
BUFx10_ASAP7_75t_L g355 ( .A(n_71), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_240), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_192), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_31), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_234), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_32), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_210), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_31), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_119), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_216), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_182), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_204), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_67), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_163), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_96), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_65), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_44), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_150), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_241), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_214), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_131), .Y(n_375) );
BUFx8_ASAP7_75t_SL g376 ( .A(n_74), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_92), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_3), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_223), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_51), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_145), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_248), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_112), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_157), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_82), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_232), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_213), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_172), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_39), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_156), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_136), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_90), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_99), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_41), .Y(n_394) );
OAI22x1_ASAP7_75t_SL g395 ( .A1(n_297), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_338), .B(n_0), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_253), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_270), .B(n_2), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_377), .B(n_4), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_283), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_285), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_285), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_253), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_312), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_253), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_285), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_254), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_292), .B(n_4), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_253), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_259), .B(n_5), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_259), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_362), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_349), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_277), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_286), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_277), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_277), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_270), .B(n_7), .Y(n_419) );
OAI22x1_ASAP7_75t_R g420 ( .A1(n_297), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_286), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_308), .B(n_9), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_278), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_385), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_299), .B(n_10), .Y(n_425) );
INVx5_ASAP7_75t_L g426 ( .A(n_278), .Y(n_426) );
CKINVDCx8_ASAP7_75t_R g427 ( .A(n_391), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_374), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_256), .A2(n_125), .B(n_124), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_278), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_361), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_281), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_281), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_281), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_281), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_404), .B(n_304), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_397), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_404), .B(n_336), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_411), .Y(n_440) );
AOI21x1_ASAP7_75t_L g441 ( .A1(n_409), .A2(n_287), .B(n_256), .Y(n_441) );
AOI21x1_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_305), .B(n_287), .Y(n_442) );
INVxp33_ASAP7_75t_L g443 ( .A(n_399), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_411), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_400), .B(n_401), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
BUFx6f_ASAP7_75t_SL g450 ( .A(n_400), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_401), .B(n_331), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_401), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_398), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_398), .Y(n_455) );
AND3x2_ASAP7_75t_L g456 ( .A(n_420), .B(n_268), .C(n_376), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_397), .Y(n_458) );
INVx11_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_398), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_419), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_402), .Y(n_465) );
OA22x2_ASAP7_75t_L g466 ( .A1(n_413), .A2(n_261), .B1(n_267), .B2(n_258), .Y(n_466) );
AO22x2_ASAP7_75t_L g467 ( .A1(n_413), .A2(n_326), .B1(n_348), .B2(n_313), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
CKINVDCx6p67_ASAP7_75t_R g469 ( .A(n_399), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_422), .B(n_313), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_402), .B(n_326), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_403), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_406), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
NOR2x1p5_ASAP7_75t_L g476 ( .A(n_428), .B(n_308), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_406), .B(n_343), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_399), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_478), .B(n_406), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_475), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_471), .B(n_427), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_478), .B(n_396), .C(n_408), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_471), .B(n_422), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_460), .B(n_416), .Y(n_485) );
BUFx8_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_454), .A2(n_425), .B(n_396), .C(n_421), .Y(n_487) );
OR2x6_ASAP7_75t_L g488 ( .A(n_467), .B(n_420), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_467), .B(n_395), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_447), .B(n_416), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_447), .B(n_421), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_455), .B(n_252), .C(n_251), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_452), .B(n_383), .C(n_289), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_439), .B(n_343), .Y(n_496) );
INVx8_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_443), .A2(n_271), .B1(n_273), .B2(n_272), .C(n_269), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_469), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_461), .B(n_344), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_475), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_469), .B(n_355), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_477), .B(n_450), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_462), .B(n_344), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_467), .B(n_355), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_462), .B(n_354), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_472), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_460), .B(n_432), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_460), .B(n_432), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_460), .B(n_432), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_476), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_474), .B(n_354), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_467), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_463), .B(n_464), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_464), .B(n_429), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_474), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_449), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_449), .B(n_303), .C(n_265), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_476), .B(n_306), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_468), .B(n_255), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_466), .B(n_355), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_451), .B(n_407), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_466), .B(n_314), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_451), .B(n_274), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_468), .B(n_429), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_470), .B(n_429), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_470), .B(n_429), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_441), .B(n_257), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_442), .B(n_407), .Y(n_536) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_438), .Y(n_537) );
NOR2x1p5_ASAP7_75t_L g538 ( .A(n_456), .B(n_376), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_438), .B(n_429), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_444), .B(n_334), .C(n_329), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_444), .B(n_412), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_459), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_444), .B(n_414), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_445), .B(n_414), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_448), .B(n_424), .Y(n_545) );
AO221x1_ASAP7_75t_L g546 ( .A1(n_457), .A2(n_395), .B1(n_319), .B2(n_359), .C(n_353), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_457), .B(n_263), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_458), .B(n_424), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_458), .B(n_431), .Y(n_549) );
OR2x6_ASAP7_75t_L g550 ( .A(n_473), .B(n_275), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_515), .A2(n_517), .B1(n_484), .B2(n_518), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_498), .A2(n_284), .B(n_288), .C(n_279), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_484), .A2(n_518), .B1(n_488), .B2(n_524), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_492), .B(n_342), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_480), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
BUFx12f_ASAP7_75t_L g557 ( .A(n_538), .Y(n_557) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_497), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_502), .B(n_319), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_499), .B(n_324), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_483), .B(n_350), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_480), .B(n_358), .Y(n_562) );
BUFx6f_ASAP7_75t_SL g563 ( .A(n_488), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_523), .B(n_324), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_531), .A2(n_534), .B(n_532), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_521), .Y(n_566) );
AOI33xp33_ASAP7_75t_L g567 ( .A1(n_526), .A2(n_431), .A3(n_309), .B1(n_296), .B2(n_316), .B3(n_298), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
AO21x1_ASAP7_75t_L g569 ( .A1(n_532), .A2(n_264), .B(n_262), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_497), .B(n_353), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_497), .B(n_359), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_539), .A2(n_276), .B(n_266), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_479), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_507), .B(n_522), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_495), .B(n_370), .C(n_367), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g577 ( .A1(n_482), .A2(n_293), .B(n_347), .C(n_327), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_489), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_486), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_539), .A2(n_282), .B(n_280), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_488), .A2(n_310), .B1(n_369), .B2(n_351), .Y(n_581) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_536), .A2(n_373), .B(n_348), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_481), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_503), .B(n_368), .Y(n_584) );
AOI33xp33_ASAP7_75t_L g585 ( .A1(n_528), .A2(n_380), .A3(n_363), .B1(n_394), .B2(n_378), .B3(n_360), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_505), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_504), .B(n_368), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_485), .A2(n_315), .B(n_294), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_485), .A2(n_318), .B(n_317), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_490), .A2(n_389), .B1(n_393), .B2(n_371), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_513), .B(n_290), .Y(n_592) );
AOI21x1_ASAP7_75t_L g593 ( .A1(n_535), .A2(n_335), .B(n_328), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_542), .B(n_310), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_490), .A2(n_351), .B1(n_369), .B2(n_332), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_529), .B(n_392), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_510), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_514), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_511), .A2(n_322), .B(n_321), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_500), .B(n_506), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_520), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_323), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_511), .A2(n_333), .B(n_330), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_496), .B(n_508), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_512), .A2(n_357), .B(n_352), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_491), .A2(n_366), .B(n_365), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_493), .A2(n_375), .B(n_372), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_494), .B(n_260), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_525), .A2(n_381), .B(n_379), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_541), .A2(n_384), .B(n_382), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_516), .B(n_291), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_490), .A2(n_390), .B(n_430), .C(n_410), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_541), .A2(n_323), .B1(n_430), .B2(n_410), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_540), .A2(n_346), .B(n_325), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_547), .B(n_295), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_546), .A2(n_323), .B1(n_301), .B2(n_302), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_545), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_548), .B(n_12), .Y(n_621) );
BUFx12f_ASAP7_75t_L g622 ( .A(n_537), .Y(n_622) );
BUFx4f_ASAP7_75t_L g623 ( .A(n_537), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_549), .A2(n_346), .B(n_325), .Y(n_624) );
BUFx8_ASAP7_75t_L g625 ( .A(n_502), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_497), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_519), .A2(n_426), .B(n_433), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_492), .B(n_12), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_492), .B(n_300), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_519), .A2(n_436), .B(n_434), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_492), .B(n_307), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_492), .B(n_311), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_499), .B(n_13), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_519), .A2(n_426), .B(n_434), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_509), .Y(n_635) );
BUFx3_ASAP7_75t_L g636 ( .A(n_486), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_492), .B(n_320), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_492), .B(n_337), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_492), .B(n_339), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_492), .B(n_340), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_509), .B(n_341), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_509), .B(n_345), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_492), .B(n_356), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_492), .B(n_14), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_509), .B(n_364), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_509), .B(n_387), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_492), .B(n_388), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_492), .B(n_15), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_492), .B(n_16), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_530), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_492), .B(n_16), .Y(n_651) );
INVx3_ASAP7_75t_L g652 ( .A(n_497), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_492), .B(n_17), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_497), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_492), .B(n_18), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_499), .B(n_18), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_492), .B(n_19), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_519), .A2(n_386), .B(n_403), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_498), .A2(n_23), .B(n_21), .C(n_22), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_492), .B(n_21), .Y(n_660) );
INVx3_ASAP7_75t_L g661 ( .A(n_497), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_492), .B(n_22), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_519), .A2(n_386), .B(n_403), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_492), .B(n_23), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_492), .B(n_25), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_SL g666 ( .A1(n_487), .A2(n_129), .B(n_130), .C(n_127), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_565), .A2(n_415), .B(n_405), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_626), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_567), .B(n_29), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_564), .B(n_30), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_620), .A2(n_415), .B1(n_417), .B2(n_405), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_555), .B(n_30), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_574), .Y(n_673) );
INVx5_ASAP7_75t_L g674 ( .A(n_626), .Y(n_674) );
OAI21x1_ASAP7_75t_L g675 ( .A1(n_582), .A2(n_417), .B(n_415), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_595), .B(n_33), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_625), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_596), .B(n_34), .Y(n_678) );
AO21x1_ASAP7_75t_L g679 ( .A1(n_553), .A2(n_417), .B(n_415), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_573), .A2(n_423), .B(n_418), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_630), .A2(n_435), .B(n_423), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_580), .A2(n_423), .B(n_418), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_580), .A2(n_423), .B(n_418), .Y(n_683) );
AOI21x1_ASAP7_75t_L g684 ( .A1(n_593), .A2(n_569), .B(n_658), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_558), .B(n_35), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_585), .B(n_35), .Y(n_686) );
AOI21xp5_ASAP7_75t_SL g687 ( .A1(n_553), .A2(n_423), .B(n_418), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_633), .Y(n_688) );
INVx5_ASAP7_75t_L g689 ( .A(n_622), .Y(n_689) );
OAI21x1_ASAP7_75t_L g690 ( .A1(n_663), .A2(n_435), .B(n_423), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_636), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_578), .Y(n_692) );
BUFx4f_ASAP7_75t_SL g693 ( .A(n_557), .Y(n_693) );
AOI21xp5_ASAP7_75t_SL g694 ( .A1(n_633), .A2(n_435), .B(n_133), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_558), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_654), .B(n_36), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_559), .B(n_37), .Y(n_697) );
AOI21xp5_ASAP7_75t_SL g698 ( .A1(n_656), .A2(n_435), .B(n_134), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_595), .B(n_37), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_635), .B(n_38), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_594), .B(n_38), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_652), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_586), .Y(n_703) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_554), .A2(n_39), .B(n_40), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_560), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_552), .B(n_42), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_551), .A2(n_47), .B1(n_45), .B2(n_46), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_581), .A2(n_48), .B1(n_45), .B2(n_47), .Y(n_708) );
AOI21xp5_ASAP7_75t_SL g709 ( .A1(n_656), .A2(n_146), .B(n_140), .Y(n_709) );
NAND2x1p5_ASAP7_75t_L g710 ( .A(n_654), .B(n_48), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_597), .A2(n_148), .B(n_147), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_652), .B(n_49), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_594), .B(n_49), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_629), .A2(n_50), .B(n_51), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_627), .A2(n_153), .B(n_152), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_615), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_623), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_628), .B(n_50), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_643), .A2(n_52), .B(n_53), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_584), .B(n_52), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_634), .A2(n_159), .B(n_154), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_644), .B(n_53), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_649), .B(n_54), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_570), .B(n_55), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_572), .B(n_57), .Y(n_725) );
OR2x6_ASAP7_75t_L g726 ( .A(n_568), .B(n_57), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_587), .B(n_58), .Y(n_727) );
OAI21xp33_ASAP7_75t_SL g728 ( .A1(n_611), .A2(n_59), .B(n_60), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_661), .B(n_59), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_604), .B(n_60), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_600), .B(n_61), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_575), .B(n_61), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_616), .Y(n_733) );
INVx3_ASAP7_75t_L g734 ( .A(n_623), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_592), .B(n_62), .Y(n_735) );
OA21x2_ASAP7_75t_L g736 ( .A1(n_624), .A2(n_169), .B(n_168), .Y(n_736) );
OAI22x1_ASAP7_75t_L g737 ( .A1(n_588), .A2(n_655), .B1(n_662), .B2(n_648), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_665), .B(n_63), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_631), .B(n_64), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_556), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_589), .A2(n_174), .B(n_173), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_561), .A2(n_64), .B(n_65), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_590), .A2(n_177), .B(n_176), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_551), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_563), .A2(n_68), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_625), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_599), .A2(n_189), .B(n_249), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_566), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_605), .B(n_73), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g750 ( .A(n_563), .B(n_73), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_632), .B(n_74), .Y(n_751) );
INVx3_ASAP7_75t_SL g752 ( .A(n_602), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_659), .A2(n_75), .B(n_76), .C(n_77), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_603), .A2(n_199), .B(n_247), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_562), .B(n_75), .Y(n_755) );
AND2x6_ASAP7_75t_L g756 ( .A(n_571), .B(n_76), .Y(n_756) );
AOI221x1_ASAP7_75t_L g757 ( .A1(n_617), .A2(n_78), .B1(n_79), .B2(n_80), .C(n_81), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_606), .A2(n_188), .B(n_246), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_641), .B(n_78), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_641), .B(n_79), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_642), .B(n_80), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_607), .A2(n_185), .B(n_239), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_608), .A2(n_183), .B(n_236), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_637), .B(n_82), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_576), .B(n_83), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_642), .B(n_83), .Y(n_766) );
BUFx5_ASAP7_75t_L g767 ( .A(n_621), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_651), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_645), .B(n_85), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_645), .B(n_646), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_646), .B(n_86), .Y(n_771) );
NAND2xp33_ASAP7_75t_L g772 ( .A(n_653), .B(n_179), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_650), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_583), .Y(n_774) );
OA22x2_ASAP7_75t_L g775 ( .A1(n_657), .A2(n_664), .B1(n_660), .B2(n_639), .Y(n_775) );
AO21x1_ASAP7_75t_L g776 ( .A1(n_613), .A2(n_180), .B(n_235), .Y(n_776) );
AOI221xp5_ASAP7_75t_SL g777 ( .A1(n_577), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_638), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_640), .B(n_88), .Y(n_779) );
AOI21x1_ASAP7_75t_L g780 ( .A1(n_614), .A2(n_205), .B(n_233), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_647), .B(n_89), .Y(n_781) );
OAI21x1_ASAP7_75t_SL g782 ( .A1(n_591), .A2(n_91), .B(n_93), .Y(n_782) );
INVx5_ASAP7_75t_L g783 ( .A(n_598), .Y(n_783) );
AO21x1_ASAP7_75t_L g784 ( .A1(n_610), .A2(n_208), .B(n_231), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_609), .B(n_94), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_612), .A2(n_95), .B(n_97), .C(n_99), .Y(n_786) );
AO31x2_ASAP7_75t_L g787 ( .A1(n_666), .A2(n_97), .A3(n_100), .B(n_101), .Y(n_787) );
OAI21xp5_ASAP7_75t_SL g788 ( .A1(n_619), .A2(n_100), .B(n_101), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_601), .B(n_102), .Y(n_789) );
O2A1O1Ixp5_ASAP7_75t_L g790 ( .A1(n_618), .A2(n_211), .B(n_229), .C(n_228), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_601), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_596), .B(n_102), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_565), .A2(n_222), .B(n_221), .Y(n_793) );
OR2x6_ASAP7_75t_L g794 ( .A(n_579), .B(n_103), .Y(n_794) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_558), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_567), .B(n_103), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_567), .B(n_104), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_659), .A2(n_104), .B(n_105), .C(n_106), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_574), .Y(n_799) );
AO31x2_ASAP7_75t_L g800 ( .A1(n_569), .A2(n_105), .A3(n_106), .B(n_107), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_558), .B(n_107), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_626), .B(n_108), .Y(n_802) );
OAI22x1_ASAP7_75t_L g803 ( .A1(n_633), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_567), .B(n_110), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_596), .B(n_111), .Y(n_805) );
NOR2xp67_ASAP7_75t_SL g806 ( .A(n_626), .B(n_112), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_567), .B(n_113), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g808 ( .A1(n_595), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_574), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_574), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_558), .B(n_114), .Y(n_811) );
NOR2x1_ASAP7_75t_SL g812 ( .A(n_674), .B(n_115), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_716), .B(n_118), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_716), .B(n_120), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_733), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_676), .A2(n_121), .B1(n_122), .B2(n_699), .Y(n_816) );
INVx1_ASAP7_75t_SL g817 ( .A(n_689), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_733), .Y(n_818) );
AO21x2_ASAP7_75t_L g819 ( .A1(n_679), .A2(n_683), .B(n_682), .Y(n_819) );
INVx2_ASAP7_75t_SL g820 ( .A(n_689), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_689), .Y(n_821) );
NOR2xp67_ASAP7_75t_L g822 ( .A(n_674), .B(n_746), .Y(n_822) );
BUFx2_ASAP7_75t_L g823 ( .A(n_677), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_681), .A2(n_684), .B(n_690), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_713), .B(n_778), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_673), .B(n_692), .Y(n_826) );
AO21x2_ASAP7_75t_L g827 ( .A1(n_680), .A2(n_687), .B(n_776), .Y(n_827) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_802), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_695), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_802), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_688), .B(n_692), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_703), .Y(n_832) );
AO21x2_ASAP7_75t_L g833 ( .A1(n_741), .A2(n_747), .B(n_743), .Y(n_833) );
INVx2_ASAP7_75t_SL g834 ( .A(n_695), .Y(n_834) );
INVx1_ASAP7_75t_SL g835 ( .A(n_696), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_703), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_790), .A2(n_780), .B(n_793), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_799), .B(n_809), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_775), .A2(n_772), .B(n_737), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_701), .B(n_678), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_672), .A2(n_760), .B(n_759), .Y(n_841) );
INVx1_ASAP7_75t_SL g842 ( .A(n_696), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_693), .Y(n_843) );
AO21x2_ASAP7_75t_L g844 ( .A1(n_754), .A2(n_758), .B(n_763), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_799), .B(n_809), .Y(n_845) );
OA21x2_ASAP7_75t_L g846 ( .A1(n_757), .A2(n_777), .B(n_762), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_715), .A2(n_721), .B(n_736), .Y(n_847) );
NAND2x1_ASAP7_75t_L g848 ( .A(n_702), .B(n_756), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_810), .B(n_748), .Y(n_849) );
INVx4_ASAP7_75t_L g850 ( .A(n_717), .Y(n_850) );
BUFx2_ASAP7_75t_L g851 ( .A(n_726), .Y(n_851) );
OAI22xp33_ASAP7_75t_SL g852 ( .A1(n_750), .A2(n_726), .B1(n_685), .B2(n_710), .Y(n_852) );
BUFx2_ASAP7_75t_R g853 ( .A(n_801), .Y(n_853) );
BUFx3_ASAP7_75t_L g854 ( .A(n_668), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_810), .Y(n_855) );
AND2x4_ASAP7_75t_L g856 ( .A(n_702), .B(n_795), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_792), .B(n_805), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_730), .Y(n_858) );
BUFx3_ASAP7_75t_L g859 ( .A(n_717), .Y(n_859) );
BUFx4f_ASAP7_75t_L g860 ( .A(n_756), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_706), .A2(n_670), .B1(n_686), .B2(n_708), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_761), .A2(n_766), .B(n_771), .Y(n_862) );
OA21x2_ASAP7_75t_L g863 ( .A1(n_784), .A2(n_704), .B(n_798), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_729), .Y(n_864) );
NAND2x1p5_ASAP7_75t_L g865 ( .A(n_717), .B(n_734), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_752), .B(n_697), .Y(n_866) );
BUFx2_ASAP7_75t_L g867 ( .A(n_756), .Y(n_867) );
NOR2xp67_ASAP7_75t_L g868 ( .A(n_691), .B(n_720), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_749), .B(n_731), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_669), .Y(n_870) );
NAND2x1p5_ASAP7_75t_L g871 ( .A(n_734), .B(n_783), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_796), .A2(n_797), .B1(n_807), .B2(n_804), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g873 ( .A(n_788), .B(n_745), .C(n_808), .Y(n_873) );
AO21x2_ASAP7_75t_L g874 ( .A1(n_769), .A2(n_732), .B(n_782), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_727), .Y(n_875) );
OA21x2_ASAP7_75t_L g876 ( .A1(n_753), .A2(n_785), .B(n_755), .Y(n_876) );
AND2x6_ASAP7_75t_L g877 ( .A(n_712), .B(n_789), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_694), .A2(n_698), .B(n_773), .Y(n_878) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_751), .A2(n_723), .B(n_722), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_773), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_718), .A2(n_738), .B(n_779), .Y(n_881) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_783), .B(n_806), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_774), .Y(n_883) );
INVx2_ASAP7_75t_SL g884 ( .A(n_783), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_774), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_700), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_709), .A2(n_781), .B(n_707), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_791), .Y(n_888) );
OAI21x1_ASAP7_75t_L g889 ( .A1(n_671), .A2(n_768), .B(n_744), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_803), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_787), .Y(n_891) );
OA21x2_ASAP7_75t_L g892 ( .A1(n_786), .A2(n_714), .B(n_719), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_724), .B(n_725), .Y(n_893) );
OAI21x1_ASAP7_75t_L g894 ( .A1(n_739), .A2(n_764), .B(n_811), .Y(n_894) );
INVx5_ASAP7_75t_L g895 ( .A(n_756), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_731), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_800), .Y(n_897) );
OAI21x1_ASAP7_75t_L g898 ( .A1(n_705), .A2(n_767), .B(n_735), .Y(n_898) );
OAI21x1_ASAP7_75t_SL g899 ( .A1(n_742), .A2(n_728), .B(n_767), .Y(n_899) );
AND2x4_ASAP7_75t_L g900 ( .A(n_765), .B(n_740), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_800), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_765), .B(n_800), .Y(n_902) );
OA21x2_ASAP7_75t_L g903 ( .A1(n_767), .A2(n_675), .B(n_582), .Y(n_903) );
BUFx12f_ASAP7_75t_L g904 ( .A(n_767), .Y(n_904) );
CKINVDCx6p67_ASAP7_75t_R g905 ( .A(n_689), .Y(n_905) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_716), .Y(n_906) );
CKINVDCx6p67_ASAP7_75t_R g907 ( .A(n_689), .Y(n_907) );
NAND2x1p5_ASAP7_75t_L g908 ( .A(n_674), .B(n_558), .Y(n_908) );
AO21x2_ASAP7_75t_L g909 ( .A1(n_679), .A2(n_683), .B(n_682), .Y(n_909) );
INVx6_ASAP7_75t_L g910 ( .A(n_689), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_677), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_688), .B(n_492), .Y(n_912) );
AOI21x1_ASAP7_75t_L g913 ( .A1(n_679), .A2(n_684), .B(n_667), .Y(n_913) );
OAI21x1_ASAP7_75t_SL g914 ( .A1(n_711), .A2(n_553), .B(n_679), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_716), .B(n_492), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_716), .Y(n_916) );
O2A1O1Ixp33_ASAP7_75t_L g917 ( .A1(n_753), .A2(n_798), .B(n_786), .C(n_659), .Y(n_917) );
BUFx10_ASAP7_75t_L g918 ( .A(n_794), .Y(n_918) );
INVxp67_ASAP7_75t_L g919 ( .A(n_756), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_689), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_689), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_688), .B(n_492), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g923 ( .A1(n_770), .A2(n_565), .B(n_517), .Y(n_923) );
AND2x4_ASAP7_75t_L g924 ( .A(n_716), .B(n_733), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_689), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_716), .Y(n_926) );
AND2x4_ASAP7_75t_L g927 ( .A(n_716), .B(n_733), .Y(n_927) );
INVx3_ASAP7_75t_L g928 ( .A(n_674), .Y(n_928) );
NAND3xp33_ASAP7_75t_L g929 ( .A(n_777), .B(n_788), .C(n_757), .Y(n_929) );
AO21x2_ASAP7_75t_L g930 ( .A1(n_679), .A2(n_683), .B(n_682), .Y(n_930) );
BUFx2_ASAP7_75t_SL g931 ( .A(n_689), .Y(n_931) );
AND2x4_ASAP7_75t_L g932 ( .A(n_716), .B(n_733), .Y(n_932) );
AO21x2_ASAP7_75t_L g933 ( .A1(n_679), .A2(n_683), .B(n_682), .Y(n_933) );
NOR2xp67_ASAP7_75t_L g934 ( .A(n_689), .B(n_568), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_770), .A2(n_565), .B(n_517), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_733), .B(n_595), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_688), .A2(n_553), .B1(n_529), .B2(n_488), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_716), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_688), .B(n_492), .Y(n_939) );
INVx3_ASAP7_75t_L g940 ( .A(n_674), .Y(n_940) );
INVx6_ASAP7_75t_L g941 ( .A(n_689), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_688), .B(n_492), .Y(n_942) );
BUFx3_ASAP7_75t_L g943 ( .A(n_689), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_716), .Y(n_944) );
INVx3_ASAP7_75t_L g945 ( .A(n_674), .Y(n_945) );
NAND2x1p5_ASAP7_75t_L g946 ( .A(n_674), .B(n_558), .Y(n_946) );
AO21x2_ASAP7_75t_L g947 ( .A1(n_679), .A2(n_683), .B(n_682), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_716), .B(n_492), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_770), .A2(n_565), .B(n_517), .Y(n_949) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_674), .Y(n_950) );
INVx4_ASAP7_75t_L g951 ( .A(n_689), .Y(n_951) );
BUFx2_ASAP7_75t_L g952 ( .A(n_689), .Y(n_952) );
AND2x4_ASAP7_75t_SL g953 ( .A(n_925), .B(n_905), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_914), .A2(n_913), .B(n_891), .Y(n_954) );
AO21x1_ASAP7_75t_L g955 ( .A1(n_897), .A2(n_901), .B(n_839), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_832), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_880), .B(n_815), .Y(n_957) );
BUFx2_ASAP7_75t_R g958 ( .A(n_931), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_836), .Y(n_959) );
BUFx3_ASAP7_75t_L g960 ( .A(n_925), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_855), .Y(n_961) );
INVx3_ASAP7_75t_L g962 ( .A(n_904), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_815), .B(n_924), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_848), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_873), .A2(n_937), .B1(n_890), .B2(n_869), .Y(n_965) );
BUFx3_ASAP7_75t_L g966 ( .A(n_908), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_818), .Y(n_967) );
BUFx3_ASAP7_75t_L g968 ( .A(n_908), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_916), .Y(n_969) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_864), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_915), .B(n_948), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_924), .B(n_927), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_926), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_938), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_860), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_944), .Y(n_976) );
BUFx3_ASAP7_75t_L g977 ( .A(n_946), .Y(n_977) );
INVx2_ASAP7_75t_SL g978 ( .A(n_910), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_906), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_838), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_826), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_824), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_845), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_849), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_843), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_867), .B(n_919), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_924), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_927), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_927), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_814), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_936), .B(n_864), .Y(n_991) );
INVx3_ASAP7_75t_L g992 ( .A(n_860), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_814), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_816), .A2(n_895), .B1(n_919), .B2(n_814), .Y(n_994) );
INVx3_ASAP7_75t_L g995 ( .A(n_895), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_838), .Y(n_996) );
OR2x6_ASAP7_75t_L g997 ( .A(n_828), .B(n_830), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_932), .Y(n_998) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_943), .Y(n_999) );
INVx6_ASAP7_75t_L g1000 ( .A(n_950), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_943), .Y(n_1001) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_852), .A2(n_851), .B1(n_895), .B2(n_918), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_813), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_870), .B(n_902), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_946), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_872), .B(n_816), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_888), .Y(n_1007) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_910), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_895), .Y(n_1009) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_907), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_912), .B(n_922), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_893), .A2(n_896), .B1(n_861), .B2(n_857), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_843), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_821), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_831), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_872), .B(n_875), .Y(n_1016) );
BUFx12f_ASAP7_75t_L g1017 ( .A(n_918), .Y(n_1017) );
INVx1_ASAP7_75t_SL g1018 ( .A(n_817), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_858), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_923), .B(n_935), .Y(n_1020) );
INVxp67_ASAP7_75t_L g1021 ( .A(n_921), .Y(n_1021) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_828), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_812), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_952), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_928), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_928), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_840), .A2(n_866), .B1(n_942), .B2(n_912), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_940), .Y(n_1028) );
AOI21x1_ASAP7_75t_L g1029 ( .A1(n_837), .A2(n_847), .B(n_846), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_949), .B(n_886), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_830), .B(n_862), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_835), .B(n_842), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_945), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_861), .A2(n_879), .B1(n_866), .B2(n_868), .Y(n_1034) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_910), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1036 ( .A(n_900), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_822), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_825), .Y(n_1038) );
CKINVDCx6p67_ASAP7_75t_R g1039 ( .A(n_951), .Y(n_1039) );
INVx4_ASAP7_75t_L g1040 ( .A(n_941), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_929), .A2(n_853), .B1(n_941), .B2(n_882), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_900), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_881), .A2(n_877), .B1(n_823), .B2(n_894), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_841), .B(n_876), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_903), .Y(n_1045) );
BUFx2_ASAP7_75t_R g1046 ( .A(n_911), .Y(n_1046) );
AOI21xp5_ASAP7_75t_SL g1047 ( .A1(n_833), .A2(n_844), .B(n_882), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_951), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_834), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1045), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_1034), .A2(n_856), .B1(n_911), .B2(n_884), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_971), .B(n_920), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1016), .B(n_1038), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1004), .B(n_885), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_957), .B(n_963), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_957), .B(n_883), .Y(n_1056) );
INVx4_ASAP7_75t_L g1057 ( .A(n_995), .Y(n_1057) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_953), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_967), .B(n_898), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_1000), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_1006), .A2(n_877), .B1(n_899), .B2(n_892), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1044), .B(n_898), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1016), .B(n_942), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1044), .B(n_876), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1065 ( .A(n_1007), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_1006), .A2(n_877), .B1(n_892), .B2(n_894), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_991), .B(n_876), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_981), .B(n_939), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_976), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_983), .B(n_939), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_972), .B(n_846), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_984), .B(n_922), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_972), .B(n_819), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_976), .Y(n_1074) );
BUFx3_ASAP7_75t_L g1075 ( .A(n_966), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1020), .B(n_819), .Y(n_1076) );
INVxp67_ASAP7_75t_L g1077 ( .A(n_1014), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_1011), .B(n_820), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_965), .A2(n_877), .B1(n_874), .B2(n_889), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_966), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_1012), .A2(n_889), .B1(n_887), .B2(n_856), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1030), .B(n_947), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1030), .B(n_909), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_980), .B(n_909), .Y(n_1084) );
OR2x6_ASAP7_75t_SL g1085 ( .A(n_994), .B(n_934), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1027), .B(n_829), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_980), .B(n_930), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_964), .B(n_878), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1031), .B(n_933), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1015), .B(n_917), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_987), .B(n_930), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_996), .B(n_854), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_979), .Y(n_1093) );
BUFx3_ASAP7_75t_L g1094 ( .A(n_968), .Y(n_1094) );
INVx1_ASAP7_75t_SL g1095 ( .A(n_953), .Y(n_1095) );
NOR2x1p5_ASAP7_75t_L g1096 ( .A(n_995), .B(n_850), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_987), .B(n_933), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_988), .B(n_863), .Y(n_1098) );
INVx3_ASAP7_75t_L g1099 ( .A(n_995), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_988), .B(n_863), .Y(n_1100) );
INVx5_ASAP7_75t_L g1101 ( .A(n_1009), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_989), .B(n_863), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_986), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_998), .B(n_827), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1069), .Y(n_1105) );
NOR2xp67_ASAP7_75t_L g1106 ( .A(n_1057), .B(n_1037), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1085), .A2(n_1043), .B1(n_1002), .B2(n_1039), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1065), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1073), .B(n_954), .Y(n_1109) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_1085), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1053), .B(n_956), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1073), .B(n_954), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1069), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1071), .B(n_1089), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1071), .B(n_954), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1050), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1067), .B(n_1022), .Y(n_1117) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1101), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1089), .B(n_955), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1074), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1063), .B(n_959), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1055), .B(n_961), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1067), .B(n_1022), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1062), .B(n_1064), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1064), .B(n_998), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1076), .B(n_970), .Y(n_1126) );
NOR2x1_ASAP7_75t_L g1127 ( .A(n_1096), .B(n_960), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1093), .B(n_969), .Y(n_1128) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_1075), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1077), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_1051), .A2(n_1039), .B1(n_1023), .B2(n_962), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1082), .B(n_982), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1083), .B(n_982), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1134 ( .A(n_1101), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1068), .B(n_973), .Y(n_1135) );
INVx3_ASAP7_75t_L g1136 ( .A(n_1057), .Y(n_1136) );
INVx3_ASAP7_75t_L g1137 ( .A(n_1057), .Y(n_1137) );
INVx2_ASAP7_75t_SL g1138 ( .A(n_1101), .Y(n_1138) );
AOI21xp33_ASAP7_75t_L g1139 ( .A1(n_1090), .A2(n_1041), .B(n_1048), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_1086), .A2(n_990), .B1(n_993), .B2(n_1036), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1084), .B(n_974), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1070), .B(n_1032), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1078), .A2(n_1052), .B1(n_1081), .B2(n_1061), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1084), .B(n_1029), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1145 ( .A(n_1088), .B(n_1009), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_1103), .A2(n_1036), .B1(n_1042), .B2(n_997), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_1075), .A2(n_1094), .B1(n_1080), .B2(n_1103), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1072), .B(n_1032), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1054), .B(n_1003), .Y(n_1149) );
BUFx3_ASAP7_75t_L g1150 ( .A(n_1080), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1105), .Y(n_1151) );
OR2x6_ASAP7_75t_L g1152 ( .A(n_1110), .B(n_1047), .Y(n_1152) );
AND2x2_ASAP7_75t_SL g1153 ( .A(n_1110), .B(n_1059), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1105), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1124), .B(n_1087), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1113), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1113), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1120), .Y(n_1158) );
BUFx6f_ASAP7_75t_L g1159 ( .A(n_1118), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1124), .B(n_1087), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_1145), .B(n_1088), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1120), .Y(n_1162) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_1145), .B(n_1088), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1114), .B(n_1104), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1126), .B(n_1059), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1109), .B(n_1091), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1116), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1109), .B(n_1091), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1112), .B(n_1097), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1141), .B(n_1121), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1112), .B(n_1097), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1108), .Y(n_1172) );
OR2x6_ASAP7_75t_L g1173 ( .A(n_1136), .B(n_1047), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1130), .B(n_1010), .Y(n_1174) );
AND2x4_ASAP7_75t_SL g1175 ( .A(n_1136), .B(n_1099), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1115), .B(n_1098), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1115), .B(n_1098), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1178 ( .A(n_1145), .B(n_1088), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1125), .B(n_1100), .Y(n_1179) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1144), .B(n_1102), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_1129), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1122), .B(n_1056), .Y(n_1182) );
INVxp67_ASAP7_75t_SL g1183 ( .A(n_1106), .Y(n_1183) );
INVxp67_ASAP7_75t_SL g1184 ( .A(n_1136), .Y(n_1184) );
NAND2xp5_ASAP7_75t_SL g1185 ( .A(n_1153), .B(n_1137), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1180), .B(n_1119), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1172), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1151), .Y(n_1188) );
NAND2x1_ASAP7_75t_L g1189 ( .A(n_1152), .B(n_1137), .Y(n_1189) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1167), .Y(n_1190) );
AND2x4_ASAP7_75t_L g1191 ( .A(n_1161), .B(n_1137), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1151), .Y(n_1192) );
NAND4xp25_ASAP7_75t_L g1193 ( .A(n_1174), .B(n_1143), .C(n_1107), .D(n_1139), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1170), .B(n_1117), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1155), .B(n_1117), .Y(n_1195) );
OAI22x1_ASAP7_75t_L g1196 ( .A1(n_1183), .A2(n_1127), .B1(n_1138), .B2(n_1118), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1155), .B(n_1123), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1180), .B(n_1132), .Y(n_1198) );
AOI32xp33_ASAP7_75t_L g1199 ( .A1(n_1181), .A2(n_1095), .A3(n_1058), .B1(n_1131), .B2(n_1147), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1154), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1160), .B(n_1133), .Y(n_1201) );
NOR2x1_ASAP7_75t_L g1202 ( .A(n_1152), .B(n_1129), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1154), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1156), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1166), .B(n_1111), .Y(n_1205) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_1153), .A2(n_1140), .B1(n_1142), .B2(n_1148), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1156), .Y(n_1207) );
INVx1_ASAP7_75t_SL g1208 ( .A(n_1175), .Y(n_1208) );
AND4x1_ASAP7_75t_L g1209 ( .A(n_1153), .B(n_958), .C(n_1046), .D(n_1066), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1195), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_1206), .A2(n_1184), .B1(n_1152), .B2(n_1165), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1199), .A2(n_1152), .B1(n_1165), .B2(n_1150), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1195), .B(n_1176), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1197), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1197), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1203), .Y(n_1216) );
AOI21xp33_ASAP7_75t_SL g1217 ( .A1(n_1185), .A2(n_1152), .B(n_985), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1190), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_1185), .A2(n_1150), .B1(n_1173), .B2(n_1134), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1203), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1188), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1192), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1200), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1204), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1193), .A2(n_1182), .B1(n_1135), .B2(n_1164), .C(n_1177), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1207), .B(n_1168), .Y(n_1226) );
INVx1_ASAP7_75t_SL g1227 ( .A(n_1208), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1187), .Y(n_1228) );
INVx1_ASAP7_75t_SL g1229 ( .A(n_1194), .Y(n_1229) );
AOI21xp5_ASAP7_75t_L g1230 ( .A1(n_1212), .A2(n_1189), .B(n_1196), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1226), .Y(n_1231) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_1225), .A2(n_1205), .B1(n_1186), .B2(n_1149), .C(n_1196), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1226), .Y(n_1233) );
OAI21xp5_ASAP7_75t_SL g1234 ( .A1(n_1217), .A2(n_1202), .B(n_1209), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1216), .Y(n_1235) );
AOI22xp5_ASAP7_75t_L g1236 ( .A1(n_1211), .A2(n_1191), .B1(n_1198), .B2(n_1163), .Y(n_1236) );
AOI22xp5_ASAP7_75t_L g1237 ( .A1(n_1227), .A2(n_1161), .B1(n_1178), .B2(n_1163), .Y(n_1237) );
NOR3xp33_ASAP7_75t_L g1238 ( .A(n_1219), .B(n_1018), .C(n_1021), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_1229), .A2(n_1178), .B1(n_1163), .B2(n_1161), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1210), .B(n_1201), .Y(n_1240) );
O2A1O1Ixp33_ASAP7_75t_L g1241 ( .A1(n_1228), .A2(n_1024), .B(n_999), .C(n_1001), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1220), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1221), .Y(n_1243) );
AOI22x1_ASAP7_75t_L g1244 ( .A1(n_1230), .A2(n_985), .B1(n_1017), .B2(n_1096), .Y(n_1244) );
NAND3xp33_ASAP7_75t_SL g1245 ( .A(n_1232), .B(n_1013), .C(n_1213), .Y(n_1245) );
NAND3xp33_ASAP7_75t_L g1246 ( .A(n_1232), .B(n_1223), .C(n_1222), .Y(n_1246) );
NAND4xp25_ASAP7_75t_L g1247 ( .A(n_1234), .B(n_1079), .C(n_1094), .D(n_1146), .Y(n_1247) );
NAND3xp33_ASAP7_75t_L g1248 ( .A(n_1236), .B(n_1224), .C(n_1215), .Y(n_1248) );
NAND3xp33_ASAP7_75t_L g1249 ( .A(n_1238), .B(n_1214), .C(n_1218), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_1231), .A2(n_1128), .B1(n_1157), .B2(n_1158), .C(n_1162), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1233), .B(n_1017), .Y(n_1251) );
OAI21xp5_ASAP7_75t_L g1252 ( .A1(n_1245), .A2(n_1241), .B(n_1237), .Y(n_1252) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_1244), .A2(n_1239), .B1(n_1243), .B2(n_1242), .C(n_1235), .Y(n_1253) );
OAI21xp5_ASAP7_75t_L g1254 ( .A1(n_1246), .A2(n_1240), .B(n_1013), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1250), .B(n_1169), .Y(n_1255) );
NOR4xp25_ASAP7_75t_L g1256 ( .A(n_1254), .B(n_1251), .C(n_1248), .D(n_1249), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1255), .Y(n_1257) );
OAI21x1_ASAP7_75t_SL g1258 ( .A1(n_1252), .A2(n_1040), .B(n_1247), .Y(n_1258) );
NOR2x1_ASAP7_75t_L g1259 ( .A(n_1253), .B(n_968), .Y(n_1259) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_1259), .B(n_1179), .Y(n_1260) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_1257), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1258), .Y(n_1262) );
NAND3xp33_ASAP7_75t_L g1263 ( .A(n_1256), .B(n_850), .C(n_1025), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1261), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1263), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_1262), .A2(n_978), .B1(n_1035), .B2(n_1008), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_1264), .A2(n_1260), .B1(n_1159), .B2(n_1040), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1265), .B(n_1190), .Y(n_1268) );
OAI22x1_ASAP7_75t_L g1269 ( .A1(n_1266), .A2(n_978), .B1(n_1008), .B2(n_1035), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1268), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_1267), .A2(n_1159), .B1(n_977), .B2(n_1005), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1269), .B(n_1171), .Y(n_1272) );
AOI21xp33_ASAP7_75t_L g1273 ( .A1(n_1270), .A2(n_1028), .B(n_1026), .Y(n_1273) );
AO22x1_ASAP7_75t_L g1274 ( .A1(n_1272), .A2(n_1005), .B1(n_977), .B2(n_859), .Y(n_1274) );
AOI21xp5_ASAP7_75t_L g1275 ( .A1(n_1274), .A2(n_1271), .B(n_871), .Y(n_1275) );
AO21x2_ASAP7_75t_L g1276 ( .A1(n_1273), .A2(n_1033), .B(n_1049), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1275), .B(n_1019), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1276), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1279 ( .A1(n_1278), .A2(n_865), .B(n_975), .Y(n_1279) );
AOI22xp5_ASAP7_75t_L g1280 ( .A1(n_1277), .A2(n_992), .B1(n_1000), .B2(n_1009), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1279), .B(n_1280), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1281), .Y(n_1282) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_1282), .A2(n_1092), .B(n_1060), .Y(n_1283) );
endmodule