module fake_jpeg_27480_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_19),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_33),
.C(n_19),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_31),
.B1(n_32),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_65),
.B1(n_23),
.B2(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_31),
.B1(n_26),
.B2(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_24),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_38),
.B1(n_27),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_79),
.B1(n_50),
.B2(n_33),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_33),
.B1(n_27),
.B2(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_81),
.B1(n_54),
.B2(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_33),
.B1(n_28),
.B2(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_33),
.B1(n_55),
.B2(n_51),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_97),
.B1(n_100),
.B2(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_34),
.C(n_35),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_99),
.B1(n_45),
.B2(n_15),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_95),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_35),
.C(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_36),
.B1(n_37),
.B2(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_105),
.B1(n_84),
.B2(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_66),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_66),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_15),
.B1(n_23),
.B2(n_30),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_66),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_82),
.B1(n_60),
.B2(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_72),
.B1(n_62),
.B2(n_67),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_12),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_97),
.B1(n_93),
.B2(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_72),
.B1(n_62),
.B2(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_131),
.Y(n_144)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_128),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_131),
.B(n_109),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_135),
.B1(n_84),
.B2(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_39),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

OAI21x1_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_39),
.B(n_35),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_39),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_107),
.C(n_84),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_30),
.B(n_25),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_18),
.B(n_17),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_45),
.B1(n_35),
.B2(n_25),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_100),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_140),
.B1(n_150),
.B2(n_156),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_141),
.B(n_153),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_121),
.B1(n_129),
.B2(n_126),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_88),
.C(n_103),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_152),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_165),
.B1(n_16),
.B2(n_29),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_106),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_148),
.B(n_159),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_87),
.B1(n_85),
.B2(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_133),
.B(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_39),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_35),
.B(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_167),
.B(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_22),
.B1(n_16),
.B2(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_162),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_114),
.A2(n_22),
.B1(n_16),
.B2(n_29),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_29),
.B1(n_18),
.B2(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_18),
.B(n_17),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_116),
.A3(n_113),
.B1(n_136),
.B2(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_180),
.B(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_184),
.B1(n_187),
.B2(n_6),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_183),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_155),
.Y(n_183)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_29),
.B1(n_14),
.B2(n_13),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_29),
.C(n_14),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_149),
.C(n_168),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_156),
.B1(n_161),
.B2(n_138),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_13),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_186),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_203),
.B(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_163),
.B1(n_164),
.B2(n_145),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_206),
.B1(n_217),
.B2(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_147),
.B1(n_152),
.B2(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_146),
.B1(n_166),
.B2(n_6),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_12),
.C(n_4),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_211),
.C(n_180),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_12),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_191),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_3),
.C(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_3),
.B(n_6),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_224),
.B1(n_235),
.B2(n_197),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_175),
.B1(n_170),
.B2(n_185),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_169),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_209),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_172),
.B1(n_173),
.B2(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_218),
.C(n_198),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_244),
.C(n_235),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_204),
.B1(n_213),
.B2(n_172),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_234),
.B1(n_228),
.B2(n_182),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_213),
.C(n_200),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_227),
.B1(n_234),
.B2(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_173),
.B1(n_206),
.B2(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_171),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

XNOR2x2_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_215),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_225),
.B(n_199),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_247),
.C(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_230),
.C(n_220),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_260),
.C(n_262),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_238),
.B(n_191),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_224),
.C(n_226),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_217),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_223),
.C(n_194),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_264),
.B1(n_182),
.B2(n_193),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_249),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_267),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_270),
.C(n_258),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_250),
.B1(n_252),
.B2(n_228),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_262),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_214),
.B(n_208),
.C(n_211),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_263),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_219),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_270),
.C(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_253),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_286),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_278),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_290),
.B(n_289),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_283),
.B(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_280),
.B1(n_176),
.B2(n_10),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_11),
.B(n_8),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_9),
.B(n_11),
.C(n_238),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_9),
.Y(n_296)
);


endmodule