module fake_jpeg_13873_n_97 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_15),
.B(n_27),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_33),
.B1(n_45),
.B2(n_40),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_51),
.B1(n_34),
.B2(n_50),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_30),
.B(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_70),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_41),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_42),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_21),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_17),
.B(n_25),
.C(n_8),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_38),
.B1(n_4),
.B2(n_6),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_34),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_51),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_88),
.A3(n_81),
.B1(n_28),
.B2(n_9),
.C1(n_11),
.C2(n_14),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_75),
.B(n_18),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_77),
.A3(n_74),
.B1(n_79),
.B2(n_76),
.C1(n_82),
.C2(n_84),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_23),
.Y(n_97)
);


endmodule