module fake_jpeg_9829_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_27),
.B1(n_32),
.B2(n_18),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_59),
.B(n_63),
.C(n_21),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_61),
.B1(n_62),
.B2(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_55),
.B1(n_28),
.B2(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_27),
.B1(n_32),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_0),
.Y(n_96)
);

OR2x4_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_33),
.B1(n_24),
.B2(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_25),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_94),
.B1(n_53),
.B2(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_79),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_40),
.A3(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_77),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_29),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_80),
.B(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_96),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_40),
.A3(n_34),
.B1(n_31),
.B2(n_25),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_63),
.B(n_44),
.Y(n_113)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_95),
.B1(n_58),
.B2(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_31),
.B1(n_25),
.B2(n_10),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_98),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

AOI21x1_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_55),
.B(n_46),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_121),
.B(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_89),
.B1(n_92),
.B2(n_53),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_67),
.C(n_69),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_52),
.C(n_51),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_124),
.Y(n_148)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_130),
.C(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_100),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_116),
.B(n_101),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_118),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_149),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_75),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_80),
.B1(n_95),
.B2(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_154)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_84),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_146),
.B(n_102),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_82),
.B1(n_45),
.B2(n_66),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_82),
.B1(n_49),
.B2(n_60),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_151),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_52),
.B1(n_86),
.B2(n_93),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_34),
.C(n_40),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_40),
.B(n_52),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_108),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_107),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_97),
.B1(n_117),
.B2(n_102),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_104),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_144),
.B(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_104),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.C(n_177),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_116),
.B(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_99),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_143),
.B1(n_133),
.B2(n_145),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_142),
.B1(n_110),
.B2(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_195),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_130),
.B1(n_151),
.B2(n_139),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_188),
.B1(n_194),
.B2(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_162),
.B1(n_152),
.B2(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_136),
.C(n_126),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_176),
.C(n_153),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_103),
.B1(n_135),
.B2(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_158),
.B(n_154),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_103),
.B1(n_85),
.B2(n_135),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_196),
.B(n_200),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_103),
.B1(n_85),
.B2(n_132),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_132),
.B1(n_109),
.B2(n_57),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_174),
.B1(n_156),
.B2(n_165),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_132),
.B1(n_57),
.B2(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_218),
.C(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_181),
.B(n_189),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_220),
.B(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_177),
.C(n_157),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_224),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_187),
.B1(n_202),
.B2(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_229),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_181),
.A2(n_174),
.B(n_57),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_0),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_232),
.A2(n_239),
.B1(n_247),
.B2(n_206),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_180),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_237),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_202),
.B1(n_191),
.B2(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_203),
.B1(n_184),
.B2(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_197),
.C(n_184),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_197),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_217),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_57),
.C(n_2),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_8),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_215),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_0),
.C(n_2),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_260),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_231),
.B(n_210),
.Y(n_261)
);

OAI321xp33_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_263),
.A3(n_264),
.B1(n_243),
.B2(n_209),
.C(n_207),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_268),
.C(n_250),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_220),
.B(n_216),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_251),
.B1(n_248),
.B2(n_208),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_265),
.A2(n_234),
.B1(n_233),
.B2(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_206),
.B1(n_247),
.B2(n_228),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_245),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_217),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_227),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_227),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_275),
.C(n_282),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_235),
.C(n_237),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_232),
.B1(n_239),
.B2(n_248),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_281),
.Y(n_289)
);

AO221x1_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_229),
.B1(n_225),
.B2(n_231),
.C(n_211),
.Y(n_278)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_280),
.B(n_14),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_253),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_9),
.B(n_13),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_10),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_297),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_259),
.B(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_7),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_272),
.C(n_276),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_281),
.C(n_283),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_304),
.B(n_14),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_6),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_296),
.B(n_298),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_7),
.B(n_11),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_4),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_287),
.B1(n_291),
.B2(n_286),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_312),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_287),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_315),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_2),
.B(n_3),
.Y(n_312)
);

AOI31xp67_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_4),
.A3(n_5),
.B(n_306),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_307),
.B(n_300),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_309),
.B(n_5),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_4),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_5),
.B(n_320),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_317),
.C(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_323),
.Y(n_326)
);


endmodule