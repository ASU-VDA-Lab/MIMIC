module fake_jpeg_20832_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_0),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_67),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_70),
.B1(n_63),
.B2(n_55),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_62),
.B1(n_73),
.B2(n_53),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_90),
.Y(n_105)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_70),
.B1(n_75),
.B2(n_52),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_99),
.B1(n_61),
.B2(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_60),
.C(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_69),
.C(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_48),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_59),
.B1(n_68),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_122),
.B1(n_113),
.B2(n_115),
.Y(n_128)
);

INVx5_ASAP7_75t_SL g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_0),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_109),
.C(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_128),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_51),
.B(n_49),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_132),
.B(n_131),
.Y(n_139)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_1),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_1),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_142),
.A3(n_127),
.B1(n_135),
.B2(n_132),
.C1(n_123),
.C2(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_126),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_25),
.B(n_42),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_17),
.C(n_39),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_148),
.C(n_149),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_145),
.C(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_16),
.C(n_36),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_13),
.B(n_35),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_12),
.A3(n_34),
.B1(n_32),
.B2(n_30),
.C1(n_27),
.C2(n_9),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_23),
.B1(n_47),
.B2(n_7),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_2),
.Y(n_161)
);


endmodule