module fake_jpeg_18968_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_8),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_31),
.B1(n_25),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_61),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_31),
.B1(n_25),
.B2(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_34),
.Y(n_65)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_31),
.B1(n_19),
.B2(n_24),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_52),
.B1(n_61),
.B2(n_51),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_89),
.B1(n_49),
.B2(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_38),
.C(n_37),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_38),
.B1(n_37),
.B2(n_16),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_81),
.B1(n_48),
.B2(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_24),
.B1(n_30),
.B2(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_56),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_98),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_109),
.B1(n_81),
.B2(n_71),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_39),
.B(n_56),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_107),
.B(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_55),
.B1(n_46),
.B2(n_59),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_55),
.B1(n_46),
.B2(n_49),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_39),
.B(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_46),
.B1(n_53),
.B2(n_48),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_48),
.B1(n_88),
.B2(n_30),
.Y(n_141)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_119),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_96),
.B(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_122),
.B(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_68),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_69),
.B(n_82),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_73),
.C(n_87),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_101),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_132),
.B1(n_137),
.B2(n_141),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_69),
.B(n_106),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_133),
.B(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_71),
.B1(n_75),
.B2(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_136),
.B1(n_127),
.B2(n_139),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_78),
.B1(n_66),
.B2(n_65),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_39),
.B(n_56),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_139),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_67),
.B1(n_53),
.B2(n_48),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_67),
.B1(n_11),
.B2(n_15),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_88),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_100),
.B(n_95),
.C(n_114),
.D(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_153),
.B1(n_161),
.B2(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_100),
.B1(n_95),
.B2(n_97),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_125),
.C(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_92),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_93),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_120),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_98),
.B1(n_88),
.B2(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_92),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_113),
.B1(n_112),
.B2(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_178),
.C(n_148),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_140),
.A3(n_128),
.B1(n_134),
.B2(n_124),
.C1(n_122),
.C2(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_193),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_134),
.C(n_120),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_165),
.B1(n_164),
.B2(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_186),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_112),
.B1(n_26),
.B2(n_21),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_186),
.B(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_26),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_172),
.B1(n_169),
.B2(n_161),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_21),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_143),
.B(n_8),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_148),
.B(n_153),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_205),
.C(n_208),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_146),
.C(n_147),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_146),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_150),
.C(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_155),
.B1(n_167),
.B2(n_21),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_181),
.A2(n_173),
.B1(n_191),
.B2(n_175),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_205),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_191),
.B(n_174),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_220),
.B(n_224),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_167),
.B(n_180),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_180),
.B(n_175),
.Y(n_224)
);

NAND4xp25_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_187),
.C(n_183),
.D(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_223),
.C(n_218),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_200),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_196),
.B1(n_194),
.B2(n_189),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_221),
.B1(n_226),
.B2(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_199),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_240),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_206),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_195),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_209),
.B(n_201),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_243),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_188),
.B(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_230),
.B(n_220),
.C(n_219),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_241),
.B(n_215),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_187),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_231),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_253),
.B1(n_247),
.B2(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_257),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_260),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_261),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_235),
.B(n_237),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_7),
.B(n_13),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_239),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_249),
.C(n_250),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_266),
.C(n_5),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_263),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_6),
.A3(n_12),
.B1(n_10),
.B2(n_3),
.C1(n_4),
.C2(n_14),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_259),
.B(n_8),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_6),
.A3(n_12),
.B1(n_11),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_267),
.A3(n_6),
.B1(n_9),
.B2(n_14),
.C1(n_2),
.C2(n_1),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_0),
.A3(n_14),
.B1(n_269),
.B2(n_229),
.C(n_63),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_274),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);


endmodule