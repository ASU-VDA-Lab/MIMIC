module fake_jpeg_30631_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_23),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_8),
.B1(n_12),
.B2(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_31),
.B1(n_16),
.B2(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_19),
.B1(n_14),
.B2(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_10),
.B1(n_16),
.B2(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_1),
.B(n_3),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_26),
.C(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_50)
);

NAND4xp25_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_40),
.C(n_3),
.D(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_26),
.C(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.Y(n_52)
);


endmodule