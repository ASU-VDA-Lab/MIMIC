module fake_jpeg_21970_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_28),
.B1(n_24),
.B2(n_39),
.Y(n_44)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_26),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_63),
.B1(n_37),
.B2(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_64),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_62),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_13),
.Y(n_56)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_10),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_37),
.B1(n_39),
.B2(n_28),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_88),
.B1(n_39),
.B2(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_77),
.B1(n_26),
.B2(n_25),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_84),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_82),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_17),
.B1(n_41),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_59),
.B1(n_62),
.B2(n_51),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_41),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_17),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_17),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_37),
.B1(n_39),
.B2(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_37),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_58),
.C(n_17),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_98),
.Y(n_123)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_93),
.A2(n_100),
.B1(n_48),
.B2(n_89),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_102),
.Y(n_135)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_24),
.Y(n_140)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_114),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_39),
.B1(n_55),
.B2(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_55),
.B1(n_53),
.B2(n_24),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_113),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_49),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_76),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_81),
.B(n_91),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_132),
.B(n_143),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_125),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_90),
.B1(n_78),
.B2(n_45),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_128),
.B1(n_134),
.B2(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_142),
.Y(n_161)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_138),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_81),
.A3(n_83),
.B1(n_109),
.B2(n_113),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_42),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_79),
.B(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_42),
.B1(n_49),
.B2(n_36),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_80),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_75),
.B(n_52),
.C(n_35),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_80),
.C(n_58),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_159),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_147),
.B(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_99),
.B1(n_42),
.B2(n_108),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_115),
.B1(n_112),
.B2(n_104),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_132),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_32),
.B1(n_112),
.B2(n_58),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_96),
.C(n_13),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_119),
.C(n_13),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_78),
.B1(n_85),
.B2(n_86),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_32),
.B1(n_74),
.B2(n_95),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_26),
.B(n_96),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_171),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_96),
.C(n_35),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_36),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_136),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_35),
.B1(n_16),
.B2(n_31),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_129),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_124),
.B1(n_144),
.B2(n_122),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_123),
.B1(n_135),
.B2(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_16),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_162),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_173),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_175),
.B(n_178),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_179),
.B(n_42),
.C(n_35),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_182),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_131),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_123),
.B(n_135),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_186),
.B(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_134),
.B(n_129),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_156),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_152),
.A2(n_165),
.B(n_153),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_163),
.B1(n_149),
.B2(n_42),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_96),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_149),
.B(n_167),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_27),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_0),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_159),
.C(n_145),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_217),
.C(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_155),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_160),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_214),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_222),
.B(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_29),
.B1(n_21),
.B2(n_15),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_47),
.C(n_46),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_35),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_181),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_47),
.C(n_46),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_15),
.B(n_31),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_30),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_240),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_183),
.B1(n_179),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_226),
.A2(n_244),
.B1(n_246),
.B2(n_22),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_177),
.B1(n_182),
.B2(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_189),
.C(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_243),
.C(n_208),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_189),
.B(n_176),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_223),
.B1(n_222),
.B2(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_198),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_174),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_36),
.C(n_30),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_201),
.B1(n_214),
.B2(n_209),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_252),
.B(n_228),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_217),
.C(n_202),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_205),
.B(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_226),
.B1(n_230),
.B2(n_237),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_223),
.B(n_218),
.C(n_23),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.C(n_231),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_235),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_30),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_21),
.B1(n_15),
.B2(n_22),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_266),
.B1(n_22),
.B2(n_23),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_36),
.C(n_23),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_263),
.C(n_265),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_30),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_21),
.C(n_30),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_230),
.B1(n_244),
.B2(n_243),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_278),
.B1(n_263),
.B2(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_281),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_10),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_11),
.Y(n_284)
);

BUFx12_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_246),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_36),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_36),
.B1(n_23),
.B2(n_19),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_12),
.C(n_11),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_280),
.Y(n_296)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_277),
.C(n_282),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.C(n_277),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_2),
.B(n_3),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_262),
.C(n_255),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_295),
.B1(n_1),
.B2(n_2),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_27),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_12),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_280),
.B1(n_282),
.B2(n_275),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_12),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_310),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_276),
.B1(n_22),
.B2(n_23),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_19),
.C(n_22),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_305),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_307),
.B(n_308),
.C(n_309),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_287),
.B(n_286),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_2),
.B(n_3),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_283),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_27),
.Y(n_310)
);

AOI21x1_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_298),
.B(n_3),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_314),
.B(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_27),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_27),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_310),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_300),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_309),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_5),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_3),
.C(n_4),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_4),
.B(n_5),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.C(n_322),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_327),
.B1(n_7),
.B2(n_8),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_7),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_7),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_9),
.Y(n_335)
);


endmodule