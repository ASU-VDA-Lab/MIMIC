module fake_jpeg_26050_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_49),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_0),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_37),
.B1(n_38),
.B2(n_17),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_4),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_10),
.B(n_11),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_75),
.B1(n_16),
.B2(n_18),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_8),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_14),
.C(n_15),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_9),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_82),
.C(n_84),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_83),
.C(n_19),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_88),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_75),
.B1(n_72),
.B2(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_85),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_34),
.Y(n_102)
);


endmodule