module fake_jpeg_6931_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_46),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_43),
.B(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_60),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_26),
.B1(n_37),
.B2(n_25),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_62),
.A2(n_65),
.B1(n_82),
.B2(n_83),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_70),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_26),
.B1(n_37),
.B2(n_25),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_31),
.B(n_29),
.C(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_68),
.B(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_31),
.B1(n_29),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_69),
.A2(n_92),
.B1(n_96),
.B2(n_5),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_75),
.Y(n_131)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_86),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_16),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_16),
.B1(n_32),
.B2(n_19),
.Y(n_92)
);

NAND2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_36),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_100),
.B1(n_104),
.B2(n_20),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_23),
.B1(n_22),
.B2(n_35),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_40),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_20),
.Y(n_106)
);

OR2x2_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_6),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_61),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_23),
.C(n_20),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_115),
.C(n_74),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_20),
.C(n_1),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_126),
.B(n_132),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_6),
.B(n_12),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_0),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_138),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_137),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_5),
.B1(n_12),
.B2(n_9),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_13),
.B1(n_4),
.B2(n_3),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_0),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_0),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_85),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_97),
.B1(n_76),
.B2(n_87),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_98),
.C(n_84),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_140),
.C(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_95),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_151),
.Y(n_190)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_81),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_159),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_65),
.B1(n_62),
.B2(n_104),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_171),
.B1(n_72),
.B2(n_109),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_2),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_110),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_71),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_165),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_167),
.Y(n_216)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_138),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_77),
.B(n_73),
.Y(n_195)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_128),
.B(n_97),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_128),
.B(n_76),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_188),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_114),
.B1(n_136),
.B2(n_85),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_180),
.B(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_136),
.B1(n_87),
.B2(n_72),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_181),
.A2(n_196),
.B1(n_161),
.B2(n_157),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_78),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_201),
.B(n_195),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_91),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_151),
.C(n_170),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_202),
.B1(n_205),
.B2(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_197),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_151),
.B(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_109),
.B1(n_135),
.B2(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_204),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_77),
.B(n_125),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_213),
.B(n_147),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_135),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_214),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_117),
.B(n_162),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_117),
.B1(n_172),
.B2(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_155),
.B1(n_146),
.B2(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_184),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_146),
.A2(n_177),
.B1(n_163),
.B2(n_169),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_163),
.B(n_165),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_160),
.Y(n_214)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_150),
.B1(n_147),
.B2(n_167),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_233),
.B1(n_187),
.B2(n_193),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_219),
.A2(n_225),
.B(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_222),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_219),
.C(n_215),
.Y(n_246)
);

NAND2x1_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_183),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_234),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_161),
.B1(n_166),
.B2(n_210),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_197),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_239),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_190),
.B(n_207),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_206),
.B(n_191),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_193),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_203),
.B1(n_192),
.B2(n_199),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_237),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_244),
.B1(n_245),
.B2(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_189),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_239),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

NOR4xp25_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_189),
.C(n_182),
.D(n_213),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_231),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_228),
.B(n_238),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_182),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_189),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_238),
.B(n_187),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_179),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_247),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_217),
.B1(n_218),
.B2(n_227),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_257),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_256),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_238),
.B1(n_223),
.B2(n_194),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_276),
.B(n_250),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_242),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_224),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_221),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_186),
.B1(n_208),
.B2(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_297),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_300),
.B(n_259),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_290),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_186),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_278),
.B(n_267),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_255),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_268),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_277),
.B(n_254),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_259),
.B(n_260),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_249),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_304),
.B(n_307),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_285),
.B(n_248),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.C(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_249),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_270),
.B1(n_275),
.B2(n_299),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_314),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_321),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_283),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

OAI321xp33_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_264),
.A3(n_265),
.B1(n_269),
.B2(n_296),
.C(n_284),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_281),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_308),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_309),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_313),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_330),
.B(n_326),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_319),
.C(n_311),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_290),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_322),
.C(n_318),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);


endmodule