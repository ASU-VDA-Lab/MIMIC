module real_jpeg_18141_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_31;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_11),
.C(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.C(n_39),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_5),
.C(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.C(n_41),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_7),
.B(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_35),
.C(n_42),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.C(n_40),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_20),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_19),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp67_ASAP7_75t_R g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_18),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_31),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule