module fake_jpeg_6307_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_39),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_18),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_43),
.B1(n_44),
.B2(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_68),
.B1(n_44),
.B2(n_36),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_37),
.B1(n_44),
.B2(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_26),
.B1(n_21),
.B2(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_60),
.B1(n_65),
.B2(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_61),
.Y(n_74)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx12f_ASAP7_75t_SL g67 ( 
.A(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_31),
.B1(n_30),
.B2(n_18),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_31),
.B1(n_38),
.B2(n_30),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_85),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_41),
.B1(n_31),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_63),
.B1(n_55),
.B2(n_66),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_86),
.B1(n_63),
.B2(n_53),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_38),
.C(n_42),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_87),
.C(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_51),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_38),
.B1(n_26),
.B2(n_21),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_38),
.C(n_42),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_21),
.B1(n_26),
.B2(n_29),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_101),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_71),
.B1(n_77),
.B2(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_62),
.B1(n_45),
.B2(n_53),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_87),
.B1(n_71),
.B2(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_22),
.B(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_108),
.C(n_79),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_62),
.B1(n_54),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_19),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_107),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_52),
.B1(n_48),
.B2(n_19),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_19),
.B1(n_27),
.B2(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_34),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_46),
.C(n_50),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_91),
.C(n_84),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_112),
.B1(n_108),
.B2(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_70),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_70),
.B1(n_82),
.B2(n_75),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_24),
.B1(n_77),
.B2(n_22),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_115),
.B1(n_114),
.B2(n_94),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_133),
.B1(n_100),
.B2(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_33),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_29),
.B1(n_24),
.B2(n_46),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_113),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_104),
.B1(n_111),
.B2(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_33),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_95),
.B(n_0),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_10),
.B(n_11),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_84),
.B(n_91),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_159),
.B1(n_162),
.B2(n_133),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_100),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_138),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_129),
.B1(n_126),
.B2(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_154),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_103),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_160),
.C(n_164),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_143),
.B1(n_164),
.B2(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_22),
.B1(n_32),
.B2(n_25),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_32),
.B1(n_25),
.B2(n_84),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_93),
.B1(n_25),
.B2(n_28),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_127),
.B(n_126),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_120),
.C(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_25),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_136),
.C(n_140),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_142),
.B(n_137),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_173),
.B1(n_186),
.B2(n_165),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_127),
.B1(n_122),
.B2(n_139),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_183),
.B1(n_162),
.B2(n_145),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_160),
.C(n_146),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_140),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_153),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_136),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_131),
.B(n_2),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_131),
.B1(n_134),
.B2(n_3),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_146),
.C(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_149),
.C(n_156),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_169),
.B1(n_163),
.B2(n_159),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_201),
.B(n_179),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_215),
.B1(n_173),
.B2(n_186),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_145),
.B1(n_166),
.B2(n_3),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_209),
.B1(n_177),
.B2(n_189),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_16),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_185),
.C(n_180),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_212),
.C(n_184),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_1),
.C(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_9),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_222),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_201),
.B1(n_200),
.B2(n_178),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_170),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_176),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_209),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_177),
.C(n_174),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_174),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_206),
.Y(n_227)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_224),
.C(n_212),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_210),
.B(n_205),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_197),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_231),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_179),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_181),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_187),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_216),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_243),
.B(n_233),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_195),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_248),
.Y(n_260)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_218),
.B(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_181),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_210),
.B(n_214),
.Y(n_243)
);

OAI22x1_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_224),
.C(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_255),
.B(n_259),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_231),
.CI(n_243),
.CON(n_254),
.SN(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_220),
.B(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_244),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_265),
.C(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_244),
.B1(n_247),
.B2(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_245),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_251),
.B(n_254),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_252),
.B1(n_256),
.B2(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_274),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_275),
.B(n_266),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_259),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_267),
.A2(n_249),
.B(n_254),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_269),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_7),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_258),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_265),
.B(n_262),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_270),
.B(n_6),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_284),
.B(n_8),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_9),
.B(n_11),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_13),
.C(n_14),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_14),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_289),
.B(n_15),
.C(n_281),
.Y(n_290)
);


endmodule