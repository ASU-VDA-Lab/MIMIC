module fake_jpeg_22336_n_236 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_25),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_43),
.B(n_23),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_25),
.B1(n_21),
.B2(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_72),
.B1(n_70),
.B2(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_17),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_73),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_22),
.B1(n_24),
.B2(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_23),
.B1(n_15),
.B2(n_20),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_26),
.B(n_14),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_52),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_50),
.C(n_36),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_69),
.B1(n_60),
.B2(n_63),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_94),
.B(n_81),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_55),
.B1(n_51),
.B2(n_40),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_98),
.B1(n_77),
.B2(n_78),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_27),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_8),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_103),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_108),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_76),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_113),
.B(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_80),
.B1(n_84),
.B2(n_91),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_76),
.Y(n_113)
);

HB1xp67_ASAP7_75t_SL g114 ( 
.A(n_94),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_52),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_37),
.B(n_35),
.C(n_38),
.D(n_14),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_89),
.C(n_98),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_85),
.B1(n_60),
.B2(n_100),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_121),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_95),
.A3(n_87),
.B1(n_14),
.B2(n_19),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_11),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_10),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_88),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_137),
.B1(n_111),
.B2(n_113),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_118),
.B1(n_119),
.B2(n_108),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_80),
.C(n_92),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_133),
.C(n_134),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_93),
.C(n_99),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_102),
.C(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_103),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_95),
.B1(n_44),
.B2(n_47),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_95),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_35),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_120),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_116),
.C(n_110),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_105),
.C(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_104),
.C(n_101),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_152),
.C(n_28),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_160),
.B1(n_137),
.B2(n_139),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_128),
.C(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_159),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_47),
.B1(n_71),
.B2(n_49),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_10),
.B(n_1),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_11),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_149),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_105),
.B(n_65),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_126),
.B(n_105),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_141),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

XNOR2x2_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_138),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_47),
.C(n_49),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_19),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_144),
.C(n_148),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_188),
.C(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_152),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_191),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_156),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_145),
.C(n_158),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_181),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_171),
.B1(n_175),
.B2(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_173),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_3),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_176),
.B1(n_172),
.B2(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.C(n_12),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_203),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_160),
.B1(n_147),
.B2(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_170),
.C(n_19),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_190),
.B1(n_188),
.B2(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_209),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_6),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_0),
.B(n_2),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_207),
.B(n_3),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_200),
.B(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_210),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_204),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_209),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_214),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_222),
.C(n_210),
.Y(n_231)
);

AO221x1_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_232),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_223),
.B1(n_6),
.B2(n_7),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_7),
.B(n_9),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_12),
.Y(n_236)
);


endmodule