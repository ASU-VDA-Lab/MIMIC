module fake_ibex_1092_n_2705 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_482, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2705);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2705;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1806;
wire n_1599;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2612;
wire n_2193;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_950;
wire n_512;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2669;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2704;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_1506;
wire n_559;

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_469),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_429),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_36),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_293),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_43),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_200),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_139),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_273),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_298),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_403),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_167),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_75),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_371),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_406),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_278),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_285),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_30),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_306),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_415),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_422),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_54),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_61),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_211),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_247),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_326),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_447),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_199),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_382),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_116),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_360),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_412),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_21),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_300),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_129),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_128),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_178),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_80),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_203),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_432),
.Y(n_532)
);

INVx4_ASAP7_75t_R g533 ( 
.A(n_311),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_38),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_411),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_369),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_473),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_56),
.Y(n_538)
);

BUFx5_ASAP7_75t_L g539 ( 
.A(n_206),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_11),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_437),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_297),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_329),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_299),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_446),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_149),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_223),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_29),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_398),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_384),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_367),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_472),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_374),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_238),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_251),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_400),
.Y(n_557)
);

BUFx5_ASAP7_75t_L g558 ( 
.A(n_163),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_22),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_89),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_140),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_79),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_30),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_66),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_125),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_356),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_200),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_466),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_186),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_237),
.B(n_55),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_99),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_95),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_413),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_78),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_46),
.Y(n_575)
);

BUFx5_ASAP7_75t_L g576 ( 
.A(n_279),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_370),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_286),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_229),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_346),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_322),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_205),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_59),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_183),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_315),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_338),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_167),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_121),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_18),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_450),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_1),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_393),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_247),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_84),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_56),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_362),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_119),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_372),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_140),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_45),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_227),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_282),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_170),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_452),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_18),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_21),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_82),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_368),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_3),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_197),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_486),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_347),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_153),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_103),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_339),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_203),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_425),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_137),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_378),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_81),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_409),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_27),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_442),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_333),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_232),
.Y(n_627)
);

BUFx5_ASAP7_75t_L g628 ( 
.A(n_126),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_468),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_31),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_65),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_459),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_454),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_292),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_444),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_104),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_182),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_33),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_379),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_354),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_228),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_419),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_390),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_262),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_158),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_489),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_389),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_352),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_73),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_202),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_228),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_154),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_349),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_291),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_149),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_332),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_64),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_479),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_418),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_336),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_253),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_106),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_399),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_222),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_63),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_276),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_302),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_244),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_314),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_42),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_467),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_77),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_60),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_301),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_305),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_180),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_490),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_475),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_51),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_33),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_202),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_22),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_32),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_383),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_5),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_407),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_269),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_100),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_73),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_387),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_232),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_483),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_122),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_462),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_39),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_45),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_132),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_68),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_317),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_227),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_82),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_11),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_252),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_53),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_263),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_52),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_394),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_359),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_357),
.B(n_481),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_434),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_144),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_355),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_266),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_28),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_48),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_49),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_328),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_132),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_25),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_348),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_219),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_144),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_122),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_151),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_138),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_451),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_190),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_169),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_482),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_256),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_1),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_337),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_430),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_121),
.B(n_15),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_221),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_27),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_381),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_105),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_420),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_480),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_74),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_195),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_426),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_164),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_31),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_295),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_55),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_340),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_212),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_364),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_376),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_95),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_465),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_36),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_170),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_287),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_445),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_231),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_351),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_308),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_455),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_13),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_120),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_470),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_107),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_198),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_41),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_161),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_280),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_221),
.Y(n_770)
);

BUFx2_ASAP7_75t_SL g771 ( 
.A(n_448),
.Y(n_771)
);

CKINVDCx14_ASAP7_75t_R g772 ( 
.A(n_98),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_294),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_401),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_363),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_290),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_463),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_212),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_66),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_119),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_178),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_46),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_153),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_90),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_142),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_488),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_146),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_57),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_189),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_135),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_90),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_307),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_240),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_175),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_182),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_152),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_190),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_80),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

CKINVDCx11_ASAP7_75t_R g800 ( 
.A(n_509),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_772),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_639),
.A2(n_255),
.B(n_254),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_510),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_710),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_510),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_510),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_504),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_510),
.Y(n_808)
);

BUFx12f_ASAP7_75t_L g809 ( 
.A(n_543),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_505),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_674),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_710),
.A2(n_258),
.B(n_257),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_710),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_543),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_622),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_539),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_539),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_539),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_672),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_622),
.B(n_652),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_543),
.Y(n_821)
);

OAI22x1_ASAP7_75t_SL g822 ( 
.A1(n_509),
.A2(n_3),
.B1(n_0),
.B2(n_2),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_587),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_772),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_610),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_763),
.B(n_0),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_539),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_763),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_523),
.B(n_259),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_572),
.Y(n_831)
);

BUFx8_ASAP7_75t_SL g832 ( 
.A(n_547),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_610),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_539),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_610),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_789),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_546),
.A2(n_627),
.B1(n_784),
.B2(n_715),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_610),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_618),
.B(n_2),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_539),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_655),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_587),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_797),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_514),
.B(n_4),
.Y(n_844)
);

OA21x2_ASAP7_75t_L g845 ( 
.A1(n_639),
.A2(n_261),
.B(n_260),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_705),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_566),
.B(n_4),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_568),
.B(n_6),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_673),
.B(n_6),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_539),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_587),
.Y(n_851)
);

BUFx8_ASAP7_75t_SL g852 ( 
.A(n_547),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_514),
.B(n_7),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_523),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_586),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_702),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_672),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_705),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_617),
.B(n_7),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_643),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_615),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_747),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_672),
.B(n_8),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_615),
.B(n_264),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_700),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_626),
.B(n_9),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_705),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_558),
.Y(n_869)
);

BUFx8_ASAP7_75t_SL g870 ( 
.A(n_592),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_700),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_558),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_586),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_658),
.B(n_10),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_558),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_642),
.A2(n_267),
.B(n_265),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_558),
.B(n_12),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_643),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_625),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_643),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_625),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_496),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_497),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_558),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_642),
.B(n_13),
.Y(n_885)
);

XOR2xp5_ASAP7_75t_L g886 ( 
.A(n_592),
.B(n_630),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_729),
.B(n_14),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_593),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_558),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_628),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_729),
.B(n_707),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_628),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_630),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_707),
.B(n_14),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_502),
.Y(n_895)
);

OAI22x1_ASAP7_75t_SL g896 ( 
.A1(n_651),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_717),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_717),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_700),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_856),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_856),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_873),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_873),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_888),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_888),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_893),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_832),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_893),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_816),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_820),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_832),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_816),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_852),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_852),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_844),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_844),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_831),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_801),
.B(n_593),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_870),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_870),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_SL g921 ( 
.A1(n_863),
.A2(n_516),
.B1(n_517),
.B2(n_515),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_801),
.B(n_606),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_841),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_809),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_R g925 ( 
.A(n_824),
.B(n_606),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_817),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_824),
.B(n_809),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_841),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_820),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_799),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_800),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_814),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_814),
.B(n_654),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_882),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_812),
.A2(n_500),
.B(n_493),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_818),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_886),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_800),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_883),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_895),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_851),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_880),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_880),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_836),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_803),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_844),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_854),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_843),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_854),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_818),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_837),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_839),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_894),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_894),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_857),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_821),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_821),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_820),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_849),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_823),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_864),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_827),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_823),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_823),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_823),
.B(n_508),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_828),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_830),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_842),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_819),
.B(n_858),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_842),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_842),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_827),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_827),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_842),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_861),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_861),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_861),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_861),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_878),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_878),
.B(n_570),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_878),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_813),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_858),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_866),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_760),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_887),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_871),
.B(n_794),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_871),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_899),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_899),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_822),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_896),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_807),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_815),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_810),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_887),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_811),
.Y(n_1000)
);

OR2x2_ASAP7_75t_SL g1001 ( 
.A(n_862),
.B(n_494),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_804),
.B(n_760),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_803),
.Y(n_1003)
);

XOR2xp5_ASAP7_75t_L g1004 ( 
.A(n_887),
.B(n_654),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_855),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_855),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_879),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_879),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_881),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_881),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_891),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_847),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_834),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_804),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_830),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_826),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_840),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_829),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_847),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_891),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_804),
.B(n_760),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_848),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_860),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_891),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_840),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_850),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_R g1027 ( 
.A(n_830),
.B(n_663),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_867),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_804),
.B(n_513),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_850),
.B(n_628),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_884),
.Y(n_1032)
);

NOR2x1p5_ASAP7_75t_L g1033 ( 
.A(n_874),
.B(n_560),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_885),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_869),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_869),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_877),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_872),
.B(n_628),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_892),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_865),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_830),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_802),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_830),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_872),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_889),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_890),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_802),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_898),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_803),
.B(n_525),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_803),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_805),
.B(n_663),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_805),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_802),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_805),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_845),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_805),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_845),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_845),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_806),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_876),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_898),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_876),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_876),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_806),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_806),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_806),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_R g1067 ( 
.A(n_808),
.B(n_527),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_808),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_808),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_808),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_825),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_825),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_825),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_825),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_833),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_833),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_975),
.B(n_628),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_976),
.B(n_628),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_965),
.B(n_492),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1047),
.A2(n_526),
.B(n_524),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_915),
.B(n_628),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_930),
.B(n_528),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_916),
.B(n_649),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_945),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_947),
.B(n_649),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_910),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_949),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_957),
.B(n_529),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_934),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_929),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_929),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_961),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1015),
.B(n_495),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_948),
.B(n_649),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1005),
.B(n_499),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_1053),
.A2(n_537),
.B(n_536),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_950),
.B(n_649),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_988),
.B(n_591),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1020),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_985),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_990),
.B(n_614),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1076),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1034),
.B(n_501),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_924),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1009),
.B(n_506),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_987),
.B(n_635),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1037),
.A2(n_1000),
.B1(n_1033),
.B2(n_1019),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_1041),
.B(n_576),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_991),
.B(n_792),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_932),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_992),
.B(n_507),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_993),
.B(n_511),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_940),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_921),
.B(n_594),
.C(n_565),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1024),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1012),
.B(n_512),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_1043),
.B(n_576),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_924),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1022),
.B(n_518),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1010),
.B(n_521),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_941),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1045),
.B(n_532),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_L g1125 ( 
.A(n_953),
.B(n_693),
.C(n_676),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1031),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_1027),
.B(n_576),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_997),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_934),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_951),
.B(n_649),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_970),
.B(n_535),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_972),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1038),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_989),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1002),
.B(n_541),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1021),
.B(n_545),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_935),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_970),
.B(n_550),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_1001),
.B(n_696),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1016),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1028),
.B(n_552),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1040),
.B(n_557),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1027),
.B(n_578),
.Y(n_1143)
);

BUFx8_ASAP7_75t_L g1144 ( 
.A(n_983),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1018),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_955),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_956),
.B(n_579),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_972),
.B(n_581),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1055),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_999),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_960),
.B(n_582),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_999),
.B(n_600),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_983),
.B(n_675),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_SL g1154 ( 
.A(n_983),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_958),
.B(n_959),
.Y(n_1155)
);

AOI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_996),
.A2(n_520),
.B1(n_522),
.B2(n_503),
.C(n_498),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1057),
.A2(n_544),
.B(n_542),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_927),
.B(n_619),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_623),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1049),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_918),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_L g1162 ( 
.A(n_923),
.B(n_770),
.C(n_538),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1051),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_964),
.A2(n_670),
.B1(n_745),
.B2(n_651),
.Y(n_1164)
);

INVx8_ASAP7_75t_L g1165 ( 
.A(n_1008),
.Y(n_1165)
);

CKINVDCx8_ASAP7_75t_R g1166 ( 
.A(n_907),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_L g1167 ( 
.A(n_1067),
.B(n_540),
.C(n_534),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_971),
.B(n_629),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_998),
.A2(n_531),
.B1(n_569),
.B2(n_562),
.C(n_530),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1014),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_963),
.B(n_966),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1029),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_968),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1004),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_967),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_973),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_974),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_1046),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_918),
.A2(n_595),
.B1(n_596),
.B2(n_588),
.C(n_585),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_978),
.B(n_632),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_979),
.B(n_633),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_980),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_936),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_981),
.B(n_634),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_982),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_936),
.Y(n_1186)
);

XOR2x2_ASAP7_75t_L g1187 ( 
.A(n_906),
.B(n_734),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_909),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_984),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_977),
.B(n_942),
.Y(n_1190)
);

AO221x1_ASAP7_75t_L g1191 ( 
.A1(n_922),
.A2(n_699),
.B1(n_748),
.B2(n_739),
.C(n_675),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_943),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_909),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_944),
.B(n_554),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_912),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1062),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1030),
.B(n_640),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1032),
.B(n_644),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_912),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_954),
.B(n_646),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_962),
.B(n_647),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1063),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1050),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1044),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_928),
.B(n_559),
.C(n_555),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1051),
.B(n_648),
.Y(n_1206)
);

AND2x6_ASAP7_75t_SL g1207 ( 
.A(n_938),
.B(n_599),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1039),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1052),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1042),
.B(n_1060),
.C(n_933),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_922),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_926),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_926),
.B(n_656),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_933),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_901),
.B(n_659),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_902),
.B(n_660),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_903),
.B(n_661),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_937),
.B(n_952),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_937),
.B(n_666),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_1054),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_925),
.B(n_667),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_952),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_925),
.B(n_669),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_911),
.Y(n_1224)
);

BUFx5_ASAP7_75t_L g1225 ( 
.A(n_1064),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_1074),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_904),
.B(n_671),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_969),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_969),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1013),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1013),
.B(n_678),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1017),
.B(n_649),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1025),
.B(n_649),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1074),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1025),
.B(n_684),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_905),
.B(n_686),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1026),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_931),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1026),
.B(n_687),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1056),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1035),
.B(n_690),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1058),
.B(n_692),
.Y(n_1242)
);

NOR3xp33_ASAP7_75t_L g1243 ( 
.A(n_994),
.B(n_563),
.C(n_561),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1036),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1036),
.Y(n_1245)
);

AND2x6_ASAP7_75t_SL g1246 ( 
.A(n_908),
.B(n_601),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1068),
.B(n_551),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_995),
.B(n_567),
.C(n_564),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1070),
.B(n_553),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1075),
.B(n_694),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1069),
.B(n_708),
.Y(n_1251)
);

AOI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_939),
.A2(n_608),
.B1(n_611),
.B2(n_607),
.C(n_602),
.Y(n_1252)
);

NOR2x1p5_ASAP7_75t_L g1253 ( 
.A(n_913),
.B(n_571),
.Y(n_1253)
);

BUFx5_ASAP7_75t_L g1254 ( 
.A(n_1065),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1071),
.Y(n_1255)
);

BUFx5_ASAP7_75t_L g1256 ( 
.A(n_1066),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1073),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1072),
.B(n_556),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1048),
.B(n_573),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1048),
.B(n_577),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1061),
.B(n_580),
.C(n_574),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1061),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_914),
.B(n_712),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_919),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_946),
.B(n_597),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_946),
.B(n_598),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_946),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_920),
.B(n_713),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_917),
.B(n_583),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1003),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1059),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1003),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1003),
.B(n_720),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1003),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1059),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1059),
.B(n_589),
.C(n_584),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1059),
.B(n_604),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_945),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_986),
.B(n_726),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_965),
.B(n_730),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1011),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1011),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_965),
.B(n_732),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_975),
.B(n_613),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_910),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_975),
.B(n_621),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1012),
.B(n_605),
.C(n_590),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_988),
.B(n_699),
.Y(n_1288)
);

AO221x1_ASAP7_75t_L g1289 ( 
.A1(n_935),
.A2(n_750),
.B1(n_748),
.B2(n_739),
.C(n_745),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1012),
.B(n_637),
.C(n_609),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_975),
.B(n_653),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_986),
.B(n_733),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_SL g1293 ( 
.A(n_983),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_965),
.B(n_737),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_986),
.B(n_740),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_921),
.B(n_645),
.C(n_638),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1011),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1012),
.B(n_664),
.C(n_657),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1011),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_910),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_975),
.B(n_743),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_910),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_975),
.B(n_757),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1011),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_965),
.B(n_746),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_910),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_975),
.B(n_769),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_986),
.B(n_751),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_965),
.B(n_753),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_986),
.B(n_756),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_986),
.B(n_761),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_910),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1150),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1208),
.B(n_750),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1082),
.B(n_665),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1128),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1140),
.B(n_679),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1145),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1100),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1087),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1134),
.B(n_612),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1165),
.B(n_771),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1137),
.B(n_548),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1117),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1146),
.B(n_519),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1224),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1166),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1090),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1091),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1115),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1165),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1092),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1126),
.B(n_549),
.Y(n_1334)
);

NOR2x2_ASAP7_75t_L g1335 ( 
.A(n_1164),
.B(n_670),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_L g1336 ( 
.A(n_1084),
.B(n_681),
.C(n_680),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1123),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1144),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1144),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1203),
.Y(n_1340)
);

O2A1O1Ixp5_ASAP7_75t_L g1341 ( 
.A1(n_1183),
.A2(n_775),
.B(n_786),
.C(n_709),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1105),
.B(n_616),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1089),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1193),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1186),
.A2(n_1218),
.B(n_1080),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1101),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1129),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1234),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1161),
.B(n_677),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1234),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1278),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1086),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1132),
.B(n_773),
.Y(n_1353)
);

INVx8_ASAP7_75t_L g1354 ( 
.A(n_1154),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1203),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1246),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1102),
.B(n_1133),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1112),
.B(n_682),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1288),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1099),
.B(n_688),
.Y(n_1360)
);

INVx5_ASAP7_75t_L g1361 ( 
.A(n_1203),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1209),
.B(n_1240),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1088),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1093),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1285),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1279),
.B(n_689),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1300),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_SL g1368 ( 
.A1(n_1118),
.A2(n_620),
.B(n_631),
.C(n_624),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1302),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1292),
.B(n_695),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1209),
.B(n_774),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1306),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1312),
.Y(n_1373)
);

AND3x1_ASAP7_75t_L g1374 ( 
.A(n_1243),
.B(n_788),
.C(n_785),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1149),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1160),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1077),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1209),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1077),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1296),
.A2(n_788),
.B1(n_785),
.B2(n_636),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1295),
.B(n_697),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1078),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1109),
.B(n_575),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1308),
.B(n_698),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1311),
.B(n_701),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_L g1386 ( 
.A(n_1149),
.B(n_759),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1310),
.B(n_703),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1121),
.B(n_704),
.Y(n_1388)
);

AND3x2_ASAP7_75t_SL g1389 ( 
.A(n_1207),
.B(n_1191),
.C(n_1289),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1240),
.B(n_776),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1220),
.B(n_641),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1204),
.B(n_716),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1116),
.A2(n_650),
.B1(n_668),
.B2(n_662),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1078),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1153),
.A2(n_719),
.B1(n_721),
.B2(n_718),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1080),
.B(n_1284),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1288),
.A2(n_724),
.B1(n_725),
.B2(n_722),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1081),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1240),
.B(n_777),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1284),
.B(n_727),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1192),
.B(n_16),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1286),
.B(n_731),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1081),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1220),
.B(n_683),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1174),
.A2(n_741),
.B1(n_742),
.B2(n_738),
.Y(n_1405)
);

NOR3xp33_ASAP7_75t_SL g1406 ( 
.A(n_1190),
.B(n_752),
.C(n_749),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1141),
.B(n_754),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1104),
.B(n_755),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1083),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1083),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1226),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1085),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1238),
.B(n_17),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1120),
.B(n_1175),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1264),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1178),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1210),
.A2(n_685),
.B1(n_706),
.B2(n_691),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1179),
.A2(n_768),
.B1(n_778),
.B2(n_765),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1286),
.B(n_779),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1154),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1291),
.B(n_781),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1139),
.A2(n_783),
.B1(n_787),
.B2(n_782),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1085),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1095),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1095),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1211),
.A2(n_791),
.B1(n_795),
.B2(n_790),
.Y(n_1426)
);

CKINVDCx14_ASAP7_75t_R g1427 ( 
.A(n_1269),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1182),
.B(n_714),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1291),
.B(n_796),
.Y(n_1429)
);

BUFx4f_ASAP7_75t_L g1430 ( 
.A(n_1176),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1098),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1205),
.A2(n_1159),
.B1(n_1108),
.B2(n_1111),
.Y(n_1432)
);

BUFx4f_ASAP7_75t_L g1433 ( 
.A(n_1177),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1098),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1130),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1079),
.B(n_723),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1281),
.B(n_1282),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1247),
.A2(n_728),
.B1(n_736),
.B2(n_735),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1130),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1103),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1194),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1178),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1163),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1301),
.B(n_744),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1200),
.B(n_766),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1196),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1253),
.B(n_1106),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1297),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1301),
.B(n_767),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1232),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1201),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1170),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1303),
.B(n_780),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1299),
.B(n_603),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1232),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1233),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1303),
.A2(n_764),
.B(n_717),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1293),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1178),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1185),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1202),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1233),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1307),
.A2(n_764),
.B(n_717),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1293),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1304),
.B(n_793),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1258),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1307),
.B(n_798),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1168),
.Y(n_1468)
);

NOR2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1287),
.B(n_1290),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1124),
.B(n_603),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1258),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1222),
.B(n_576),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1237),
.B(n_1244),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1125),
.B(n_19),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1259),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1259),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1215),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1216),
.B(n_19),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1147),
.A2(n_762),
.B1(n_764),
.B2(n_833),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1298),
.A2(n_762),
.B1(n_764),
.B2(n_24),
.Y(n_1480)
);

O2A1O1Ixp5_ASAP7_75t_L g1481 ( 
.A1(n_1242),
.A2(n_533),
.B(n_762),
.C(n_270),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1217),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1188),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1189),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1135),
.B(n_833),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1255),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1173),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1260),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1172),
.B(n_20),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1260),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1151),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1097),
.B(n_20),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1113),
.B(n_1114),
.Y(n_1493)
);

AND3x2_ASAP7_75t_SL g1494 ( 
.A(n_1187),
.B(n_23),
.C(n_24),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1257),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1249),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1156),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1249),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1227),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1136),
.B(n_835),
.Y(n_1500)
);

AND2x6_ASAP7_75t_SL g1501 ( 
.A(n_1236),
.B(n_23),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1197),
.B(n_25),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1195),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1157),
.B(n_26),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1280),
.B(n_26),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1152),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1169),
.A2(n_838),
.B1(n_846),
.B2(n_835),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1283),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1276),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1294),
.B(n_28),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1305),
.B(n_29),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1265),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_R g1513 ( 
.A(n_1127),
.B(n_32),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1263),
.Y(n_1514)
);

NAND2xp33_ASAP7_75t_SL g1515 ( 
.A(n_1094),
.B(n_835),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1265),
.Y(n_1516)
);

INVx5_ASAP7_75t_L g1517 ( 
.A(n_1199),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1309),
.B(n_34),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1157),
.B(n_1212),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1155),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1213),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1198),
.B(n_35),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1266),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1268),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1142),
.B(n_37),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1266),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1277),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1162),
.A2(n_838),
.B1(n_846),
.B2(n_835),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1181),
.Y(n_1529)
);

AND2x6_ASAP7_75t_SL g1530 ( 
.A(n_1171),
.B(n_37),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1167),
.B(n_838),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1252),
.A2(n_846),
.B1(n_853),
.B2(n_838),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1221),
.B(n_39),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1214),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1228),
.B(n_40),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1223),
.B(n_40),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1143),
.A2(n_853),
.B1(n_859),
.B2(n_846),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1277),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1229),
.B(n_41),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1230),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1219),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_L g1542 ( 
.A(n_1245),
.B(n_853),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1261),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1231),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1158),
.Y(n_1545)
);

AND2x6_ASAP7_75t_L g1546 ( 
.A(n_1273),
.B(n_853),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1235),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1206),
.A2(n_868),
.B1(n_897),
.B2(n_859),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1131),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1148),
.A2(n_48),
.B(n_44),
.C(n_47),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1096),
.B(n_1107),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1110),
.A2(n_897),
.B(n_868),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1239),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1138),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1241),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1122),
.A2(n_897),
.B1(n_898),
.B2(n_868),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1180),
.B(n_44),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1250),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1225),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1251),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1184),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1225),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1248),
.A2(n_1119),
.B1(n_1256),
.B2(n_1254),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1254),
.B(n_49),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1254),
.B(n_50),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1254),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1254),
.B(n_50),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1256),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1271),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1256),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1262),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1571)
);

INVx5_ASAP7_75t_L g1572 ( 
.A(n_1275),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1267),
.A2(n_58),
.B1(n_54),
.B2(n_57),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1270),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1317),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1497),
.B(n_58),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1351),
.Y(n_1577)
);

O2A1O1Ixp5_ASAP7_75t_SL g1578 ( 
.A1(n_1362),
.A2(n_1274),
.B(n_1272),
.C(n_271),
.Y(n_1578)
);

AOI22x1_ASAP7_75t_L g1579 ( 
.A1(n_1457),
.A2(n_272),
.B1(n_274),
.B2(n_268),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1376),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1345),
.A2(n_277),
.B(n_275),
.Y(n_1581)
);

AND2x2_ASAP7_75t_SL g1582 ( 
.A(n_1386),
.B(n_59),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1557),
.A2(n_283),
.B(n_284),
.C(n_281),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1319),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1496),
.B(n_62),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1363),
.B(n_67),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1396),
.A2(n_289),
.B(n_288),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1315),
.B(n_69),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1498),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_SL g1590 ( 
.A(n_1328),
.B(n_70),
.C(n_71),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1340),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1374),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1400),
.B(n_76),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1321),
.B(n_1391),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1375),
.B(n_296),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1357),
.A2(n_79),
.B(n_76),
.C(n_78),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1346),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1400),
.B(n_81),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1402),
.B(n_83),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1489),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1600)
);

A2O1A1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1506),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1402),
.B(n_86),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1440),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1466),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1491),
.A2(n_92),
.B(n_88),
.C(n_91),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1471),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1338),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1475),
.A2(n_96),
.B1(n_93),
.B2(n_94),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1339),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1377),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1320),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1325),
.B(n_97),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1340),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_SL g1614 ( 
.A(n_1323),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1489),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1391),
.B(n_101),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1561),
.B(n_102),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1315),
.B(n_102),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1510),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1438),
.B(n_108),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1404),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1452),
.B(n_109),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1507),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1350),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_1327),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1392),
.B(n_110),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1473),
.A2(n_304),
.B(n_303),
.Y(n_1627)
);

INVx5_ASAP7_75t_L g1628 ( 
.A(n_1354),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1329),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1392),
.B(n_111),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1447),
.B(n_112),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1507),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1324),
.B(n_115),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1379),
.A2(n_310),
.B(n_309),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1520),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1355),
.B(n_115),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1476),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1331),
.B(n_117),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1322),
.B(n_118),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1337),
.B(n_1326),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1534),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1322),
.B(n_120),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1465),
.B(n_123),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1422),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1382),
.A2(n_1398),
.B(n_1394),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1465),
.B(n_124),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1355),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1488),
.A2(n_129),
.B1(n_126),
.B2(n_127),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1419),
.B(n_127),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1540),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1403),
.A2(n_133),
.B(n_130),
.C(n_131),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1330),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1446),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1421),
.B(n_130),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1333),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1313),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1429),
.B(n_131),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1490),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_L g1659 ( 
.A(n_1356),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1326),
.B(n_134),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1409),
.A2(n_1412),
.B(n_1410),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1467),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1446),
.B(n_312),
.Y(n_1663)
);

CKINVDCx11_ASAP7_75t_R g1664 ( 
.A(n_1323),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1467),
.B(n_136),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1447),
.B(n_139),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_L g1667 ( 
.A(n_1451),
.B(n_141),
.C(n_142),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1352),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1423),
.A2(n_145),
.B1(n_141),
.B2(n_143),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1445),
.B(n_143),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1361),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1361),
.Y(n_1672)
);

CKINVDCx10_ASAP7_75t_R g1673 ( 
.A(n_1323),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1364),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1424),
.A2(n_316),
.B(n_313),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1425),
.A2(n_319),
.B(n_318),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1432),
.B(n_145),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1361),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1411),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1510),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1469),
.B(n_147),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1378),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1517),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1431),
.A2(n_321),
.B(n_320),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1434),
.A2(n_324),
.B(n_323),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1474),
.A2(n_148),
.B(n_150),
.C(n_151),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_R g1687 ( 
.A(n_1415),
.B(n_150),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1359),
.B(n_1441),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1435),
.A2(n_327),
.B(n_325),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1348),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1517),
.B(n_155),
.Y(n_1691)
);

NOR2x1_ASAP7_75t_L g1692 ( 
.A(n_1447),
.B(n_155),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1349),
.B(n_156),
.C(n_157),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1365),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1334),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1341),
.B(n_156),
.C(n_157),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1483),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1334),
.B(n_158),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1468),
.B(n_159),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1439),
.A2(n_160),
.B(n_161),
.C(n_162),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1502),
.A2(n_160),
.B(n_162),
.C(n_163),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1522),
.A2(n_164),
.B(n_165),
.C(n_166),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1367),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1369),
.Y(n_1704)
);

NAND2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1314),
.B(n_1332),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1450),
.A2(n_331),
.B(n_330),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1455),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1335),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1426),
.B(n_171),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1443),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1460),
.B(n_171),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1372),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1373),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1483),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1422),
.A2(n_1405),
.B1(n_1380),
.B2(n_1518),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1397),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1483),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1559),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1395),
.B(n_173),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1477),
.B(n_174),
.C(n_175),
.Y(n_1720)
);

OR2x6_ASAP7_75t_L g1721 ( 
.A(n_1354),
.B(n_176),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1354),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1430),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1559),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1444),
.B(n_176),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_SL g1726 ( 
.A(n_1513),
.B(n_177),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1456),
.A2(n_335),
.B(n_334),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1358),
.B(n_177),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1462),
.A2(n_342),
.B(n_341),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1521),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1481),
.A2(n_344),
.B(n_343),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1436),
.A2(n_179),
.B1(n_181),
.B2(n_183),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1485),
.A2(n_1500),
.B(n_1461),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1383),
.B(n_1508),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1316),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1318),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1512),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1393),
.B(n_187),
.C(n_188),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_R g1739 ( 
.A(n_1343),
.B(n_188),
.Y(n_1739)
);

AO21x1_ASAP7_75t_L g1740 ( 
.A1(n_1492),
.A2(n_350),
.B(n_345),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1428),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1418),
.B(n_189),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1427),
.B(n_191),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1449),
.A2(n_1453),
.B(n_1550),
.C(n_1360),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1533),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1536),
.A2(n_192),
.B(n_193),
.C(n_194),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1541),
.B(n_194),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1342),
.B(n_195),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1420),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1493),
.B(n_196),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1342),
.Y(n_1751)
);

OR2x6_ASAP7_75t_SL g1752 ( 
.A(n_1458),
.B(n_196),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1428),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1503),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1487),
.Y(n_1755)
);

OAI21x1_ASAP7_75t_L g1756 ( 
.A1(n_1463),
.A2(n_358),
.B(n_353),
.Y(n_1756)
);

O2A1O1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1525),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1544),
.B(n_201),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1414),
.B(n_201),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1516),
.A2(n_388),
.B(n_487),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1523),
.A2(n_386),
.B(n_485),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1414),
.B(n_204),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1484),
.B(n_204),
.Y(n_1763)
);

AO21x1_ASAP7_75t_L g1764 ( 
.A1(n_1504),
.A2(n_391),
.B(n_484),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1503),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1433),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1374),
.B(n_207),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1464),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1478),
.B(n_208),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1526),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1527),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_R g1772 ( 
.A(n_1347),
.B(n_209),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1406),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1538),
.A2(n_395),
.B(n_478),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1417),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_SL g1776 ( 
.A(n_1499),
.B(n_213),
.C(n_214),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1388),
.B(n_215),
.Y(n_1777)
);

INVx8_ASAP7_75t_L g1778 ( 
.A(n_1549),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1552),
.A2(n_397),
.B(n_477),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1574),
.A2(n_396),
.B(n_476),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_SL g1781 ( 
.A(n_1568),
.B(n_361),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1408),
.A2(n_215),
.B(n_216),
.C(n_217),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1472),
.A2(n_402),
.B(n_474),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1413),
.B(n_1401),
.Y(n_1784)
);

INVx6_ASAP7_75t_L g1785 ( 
.A(n_1487),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1407),
.B(n_216),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1336),
.B(n_217),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1486),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1482),
.B(n_218),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1495),
.B(n_218),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1535),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1505),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_1792)
);

AO21x1_ASAP7_75t_L g1793 ( 
.A1(n_1504),
.A2(n_404),
.B(n_471),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1539),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1549),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1558),
.B(n_220),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1366),
.A2(n_223),
.B(n_224),
.C(n_225),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1560),
.B(n_224),
.Y(n_1798)
);

INVx4_ASAP7_75t_L g1799 ( 
.A(n_1448),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1511),
.B(n_225),
.Y(n_1800)
);

AND2x2_ASAP7_75t_SL g1801 ( 
.A(n_1389),
.B(n_226),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1448),
.B(n_226),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1529),
.B(n_1437),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1543),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1573),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1370),
.B(n_230),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1381),
.B(n_233),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1570),
.Y(n_1808)
);

CKINVDCx20_ASAP7_75t_R g1809 ( 
.A(n_1514),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1563),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1564),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1480),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1384),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1547),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1501),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1344),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1385),
.B(n_241),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1553),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1524),
.B(n_241),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1387),
.B(n_242),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1545),
.B(n_242),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1555),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1416),
.A2(n_1459),
.B(n_1442),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1532),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1551),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1825)
);

AOI21x1_ASAP7_75t_L g1826 ( 
.A1(n_1531),
.A2(n_417),
.B(n_464),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1565),
.A2(n_245),
.B(n_246),
.C(n_248),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1562),
.A2(n_416),
.B(n_461),
.Y(n_1828)
);

CKINVDCx16_ASAP7_75t_R g1829 ( 
.A(n_1480),
.Y(n_1829)
);

BUFx4f_ASAP7_75t_L g1830 ( 
.A(n_1549),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1566),
.A2(n_414),
.B(n_460),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1371),
.B(n_246),
.Y(n_1832)
);

AOI22x1_ASAP7_75t_SL g1833 ( 
.A1(n_1494),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1571),
.B(n_249),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1554),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1390),
.B(n_252),
.Y(n_1836)
);

OAI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1528),
.A2(n_365),
.B(n_366),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1501),
.Y(n_1838)
);

BUFx8_ASAP7_75t_L g1839 ( 
.A(n_1509),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1567),
.A2(n_373),
.B1(n_375),
.B2(n_377),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1399),
.B(n_1353),
.Y(n_1841)
);

NOR3xp33_ASAP7_75t_SL g1842 ( 
.A(n_1515),
.B(n_380),
.C(n_385),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1470),
.A2(n_392),
.B(n_405),
.Y(n_1843)
);

CKINVDCx12_ASAP7_75t_R g1844 ( 
.A(n_1530),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1572),
.A2(n_408),
.B1(n_423),
.B2(n_424),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1454),
.B(n_491),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1556),
.A2(n_427),
.B(n_428),
.C(n_431),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1530),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1479),
.B(n_433),
.C(n_435),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1569),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1548),
.B(n_436),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1537),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1546),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1542),
.A2(n_449),
.B(n_453),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1546),
.Y(n_1855)
);

INVx11_ASAP7_75t_L g1856 ( 
.A(n_1546),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1354),
.B(n_457),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1374),
.A2(n_458),
.B1(n_893),
.B2(n_886),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1376),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1497),
.B(n_1376),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1321),
.B(n_1351),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1497),
.B(n_1137),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1354),
.Y(n_1863)
);

CKINVDCx12_ASAP7_75t_R g1864 ( 
.A(n_1323),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1519),
.A2(n_1345),
.B(n_1053),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1368),
.A2(n_921),
.B(n_1357),
.C(n_1497),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1497),
.B(n_1376),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1351),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1497),
.B(n_1137),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1396),
.A2(n_1058),
.B(n_1345),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1351),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1497),
.B(n_1376),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1497),
.A2(n_1496),
.B1(n_1498),
.B2(n_1396),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1497),
.A2(n_1496),
.B1(n_1498),
.B2(n_1396),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1328),
.Y(n_1875)
);

INVx3_ASAP7_75t_SL g1876 ( 
.A(n_1328),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1351),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1376),
.B(n_1561),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1497),
.B(n_1137),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1396),
.A2(n_1498),
.B1(n_1496),
.B2(n_1471),
.Y(n_1880)
);

AOI21x1_ASAP7_75t_L g1881 ( 
.A1(n_1519),
.A2(n_1504),
.B(n_1492),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1497),
.B(n_1376),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1376),
.B(n_1561),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1376),
.B(n_1561),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_SL g1885 ( 
.A(n_1432),
.B(n_901),
.C(n_900),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1580),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1744),
.A2(n_1661),
.B(n_1645),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1672),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1635),
.B(n_1577),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1880),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1859),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1672),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1878),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1625),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1881),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1873),
.B(n_1874),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1628),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1883),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1884),
.B(n_1621),
.Y(n_1899)
);

AO21x2_ASAP7_75t_L g1900 ( 
.A1(n_1731),
.A2(n_1581),
.B(n_1740),
.Y(n_1900)
);

CKINVDCx20_ASAP7_75t_R g1901 ( 
.A(n_1664),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1884),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1603),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1873),
.B(n_1874),
.Y(n_1904)
);

BUFx8_ASAP7_75t_SL g1905 ( 
.A(n_1659),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1628),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1575),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1584),
.Y(n_1908)
);

CKINVDCx8_ASAP7_75t_R g1909 ( 
.A(n_1673),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1672),
.Y(n_1910)
);

AOI22x1_ASAP7_75t_L g1911 ( 
.A1(n_1634),
.A2(n_1676),
.B1(n_1684),
.B2(n_1675),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1611),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1628),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1770),
.A2(n_1794),
.B(n_1791),
.Y(n_1914)
);

OAI21x1_ASAP7_75t_L g1915 ( 
.A1(n_1826),
.A2(n_1823),
.B(n_1779),
.Y(n_1915)
);

AO21x2_ASAP7_75t_L g1916 ( 
.A1(n_1764),
.A2(n_1793),
.B(n_1696),
.Y(n_1916)
);

BUFx2_ASAP7_75t_R g1917 ( 
.A(n_1755),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1629),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1751),
.A2(n_1617),
.B1(n_1680),
.B2(n_1619),
.Y(n_1919)
);

NAND2x1p5_ASAP7_75t_L g1920 ( 
.A(n_1591),
.B(n_1613),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_SL g1921 ( 
.A1(n_1828),
.A2(n_1680),
.B(n_1619),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1862),
.B(n_1869),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1871),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1879),
.B(n_1715),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1652),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1655),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1756),
.A2(n_1733),
.B(n_1587),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1803),
.B(n_1594),
.Y(n_1928)
);

INVx2_ASAP7_75t_SL g1929 ( 
.A(n_1673),
.Y(n_1929)
);

BUFx2_ASAP7_75t_R g1930 ( 
.A(n_1875),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1803),
.B(n_1799),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1722),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1696),
.A2(n_1783),
.B(n_1583),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1868),
.Y(n_1934)
);

AOI22x1_ASAP7_75t_L g1935 ( 
.A1(n_1685),
.A2(n_1689),
.B1(n_1727),
.B2(n_1706),
.Y(n_1935)
);

OAI21x1_ASAP7_75t_L g1936 ( 
.A1(n_1850),
.A2(n_1579),
.B(n_1627),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1860),
.B(n_1867),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1710),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1591),
.B(n_1613),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1708),
.A2(n_1858),
.B1(n_1805),
.B2(n_1582),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_SL g1941 ( 
.A1(n_1643),
.A2(n_1646),
.B(n_1642),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_SL g1942 ( 
.A1(n_1639),
.A2(n_1840),
.B(n_1732),
.Y(n_1942)
);

INVx2_ASAP7_75t_SL g1943 ( 
.A(n_1785),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1597),
.Y(n_1944)
);

INVx4_ASAP7_75t_L g1945 ( 
.A(n_1785),
.Y(n_1945)
);

AOI22x1_ASAP7_75t_L g1946 ( 
.A1(n_1729),
.A2(n_1760),
.B1(n_1774),
.B2(n_1761),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1849),
.A2(n_1842),
.B(n_1837),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1656),
.Y(n_1948)
);

AO21x2_ASAP7_75t_L g1949 ( 
.A1(n_1837),
.A2(n_1802),
.B(n_1665),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1806),
.A2(n_1817),
.B(n_1807),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1671),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1857),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1641),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_SL g1954 ( 
.A(n_1721),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1647),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1650),
.Y(n_1956)
);

BUFx12f_ASAP7_75t_L g1957 ( 
.A(n_1721),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1640),
.B(n_1730),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1694),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1678),
.Y(n_1960)
);

AO21x2_ASAP7_75t_L g1961 ( 
.A1(n_1824),
.A2(n_1598),
.B(n_1593),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1780),
.A2(n_1831),
.B(n_1784),
.Y(n_1962)
);

BUFx2_ASAP7_75t_SL g1963 ( 
.A(n_1614),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1622),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1751),
.Y(n_1965)
);

BUFx2_ASAP7_75t_SL g1966 ( 
.A(n_1614),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1622),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1854),
.A2(n_1843),
.B(n_1845),
.Y(n_1968)
);

BUFx4f_ASAP7_75t_L g1969 ( 
.A(n_1857),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1607),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1659),
.Y(n_1971)
);

INVx6_ASAP7_75t_L g1972 ( 
.A(n_1682),
.Y(n_1972)
);

AO21x2_ASAP7_75t_L g1973 ( 
.A1(n_1599),
.A2(n_1602),
.B(n_1626),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1609),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1750),
.A2(n_1866),
.B(n_1736),
.Y(n_1975)
);

AO21x2_ASAP7_75t_L g1976 ( 
.A1(n_1630),
.A2(n_1840),
.B(n_1820),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1698),
.A2(n_1654),
.B(n_1649),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1734),
.B(n_1872),
.Y(n_1978)
);

CKINVDCx16_ASAP7_75t_R g1979 ( 
.A(n_1749),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1703),
.Y(n_1980)
);

BUFx4_ASAP7_75t_SL g1981 ( 
.A(n_1721),
.Y(n_1981)
);

OR3x4_ASAP7_75t_SL g1982 ( 
.A(n_1844),
.B(n_1833),
.C(n_1864),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1683),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1704),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1877),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1683),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1624),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1754),
.A2(n_1765),
.B(n_1851),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1653),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1882),
.B(n_1885),
.Y(n_1990)
);

OR2x6_ASAP7_75t_L g1991 ( 
.A(n_1857),
.B(n_1723),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1712),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1617),
.Y(n_1993)
);

OAI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1657),
.A2(n_1660),
.B(n_1618),
.Y(n_1994)
);

AO21x2_ASAP7_75t_L g1995 ( 
.A1(n_1585),
.A2(n_1677),
.B(n_1612),
.Y(n_1995)
);

CKINVDCx8_ASAP7_75t_R g1996 ( 
.A(n_1766),
.Y(n_1996)
);

AO21x1_ASAP7_75t_L g1997 ( 
.A1(n_1726),
.A2(n_1810),
.B(n_1781),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1713),
.Y(n_1998)
);

BUFx4f_ASAP7_75t_SL g1999 ( 
.A(n_1876),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1789),
.B(n_1801),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1691),
.A2(n_1636),
.B(n_1816),
.Y(n_2001)
);

BUFx2_ASAP7_75t_L g2002 ( 
.A(n_1809),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1803),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_SL g2004 ( 
.A(n_1863),
.B(n_1773),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_SL g2005 ( 
.A1(n_1732),
.A2(n_1812),
.B(n_1666),
.Y(n_2005)
);

CKINVDCx14_ASAP7_75t_R g2006 ( 
.A(n_1687),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1679),
.Y(n_2007)
);

CKINVDCx16_ASAP7_75t_R g2008 ( 
.A(n_1739),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1768),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1711),
.Y(n_2010)
);

NAND2x1p5_ASAP7_75t_L g2011 ( 
.A(n_1682),
.B(n_1830),
.Y(n_2011)
);

BUFx8_ASAP7_75t_L g2012 ( 
.A(n_1848),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1772),
.Y(n_2013)
);

OAI21x1_ASAP7_75t_L g2014 ( 
.A1(n_1600),
.A2(n_1615),
.B(n_1668),
.Y(n_2014)
);

BUFx12f_ASAP7_75t_L g2015 ( 
.A(n_1839),
.Y(n_2015)
);

AO21x2_ASAP7_75t_L g2016 ( 
.A1(n_1827),
.A2(n_1725),
.B(n_1800),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1633),
.A2(n_1829),
.B1(n_1858),
.B2(n_1759),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1711),
.Y(n_2018)
);

BUFx2_ASAP7_75t_SL g2019 ( 
.A(n_1682),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1674),
.Y(n_2020)
);

AO21x1_ASAP7_75t_SL g2021 ( 
.A1(n_1856),
.A2(n_1812),
.B(n_1788),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1741),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_L g2023 ( 
.A1(n_1757),
.A2(n_1701),
.B(n_1702),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1752),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1596),
.A2(n_1662),
.B(n_1623),
.Y(n_2025)
);

BUFx2_ASAP7_75t_SL g2026 ( 
.A(n_1798),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1753),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1705),
.Y(n_2028)
);

AO21x2_ASAP7_75t_L g2029 ( 
.A1(n_1847),
.A2(n_1606),
.B(n_1589),
.Y(n_2029)
);

OAI21x1_ASAP7_75t_L g2030 ( 
.A1(n_1632),
.A2(n_1797),
.B(n_1782),
.Y(n_2030)
);

NAND2x1p5_ASAP7_75t_L g2031 ( 
.A(n_1830),
.B(n_1855),
.Y(n_2031)
);

NAND2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1855),
.B(n_1697),
.Y(n_2032)
);

INVx4_ASAP7_75t_L g2033 ( 
.A(n_1778),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1839),
.Y(n_2034)
);

BUFx5_ASAP7_75t_L g2035 ( 
.A(n_1835),
.Y(n_2035)
);

AO21x2_ASAP7_75t_L g2036 ( 
.A1(n_1610),
.A2(n_1700),
.B(n_1651),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1690),
.B(n_1748),
.Y(n_2037)
);

OAI21x1_ASAP7_75t_L g2038 ( 
.A1(n_1735),
.A2(n_1796),
.B(n_1790),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1777),
.A2(n_1786),
.B(n_1670),
.Y(n_2039)
);

AO21x2_ASAP7_75t_L g2040 ( 
.A1(n_1601),
.A2(n_1605),
.B(n_1746),
.Y(n_2040)
);

BUFx10_ASAP7_75t_L g2041 ( 
.A(n_1798),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1586),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1814),
.B(n_1818),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1822),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1588),
.Y(n_2045)
);

BUFx5_ASAP7_75t_L g2046 ( 
.A(n_1846),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1815),
.Y(n_2047)
);

INVx3_ASAP7_75t_L g2048 ( 
.A(n_1718),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1838),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_1861),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1811),
.A2(n_1745),
.B(n_1738),
.Y(n_2051)
);

AO21x2_ASAP7_75t_L g2052 ( 
.A1(n_1738),
.A2(n_1719),
.B(n_1716),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1688),
.B(n_1576),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1718),
.Y(n_2054)
);

CKINVDCx20_ASAP7_75t_R g2055 ( 
.A(n_1592),
.Y(n_2055)
);

OAI21x1_ASAP7_75t_L g2056 ( 
.A1(n_1616),
.A2(n_1604),
.B(n_1771),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1747),
.B(n_1758),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1819),
.B(n_1699),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1720),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_1795),
.B(n_1808),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1742),
.Y(n_2061)
);

CKINVDCx16_ASAP7_75t_R g2062 ( 
.A(n_1592),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1724),
.B(n_1808),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_1778),
.Y(n_2064)
);

INVx8_ASAP7_75t_L g2065 ( 
.A(n_1778),
.Y(n_2065)
);

OA21x2_ASAP7_75t_L g2066 ( 
.A1(n_1811),
.A2(n_1804),
.B(n_1792),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_L g2067 ( 
.A1(n_1737),
.A2(n_1669),
.B(n_1707),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1832),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1714),
.Y(n_2069)
);

INVx6_ASAP7_75t_L g2070 ( 
.A(n_1724),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_1631),
.B(n_1692),
.Y(n_2071)
);

OAI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1728),
.A2(n_1620),
.B(n_1763),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1608),
.Y(n_2073)
);

AO21x2_ASAP7_75t_L g2074 ( 
.A1(n_1667),
.A2(n_1813),
.B(n_1693),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1717),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1637),
.A2(n_1648),
.B(n_1658),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1853),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1825),
.A2(n_1686),
.B(n_1775),
.Y(n_2078)
);

OR2x6_ASAP7_75t_L g2079 ( 
.A(n_1832),
.B(n_1836),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1836),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1787),
.A2(n_1709),
.B(n_1769),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1841),
.A2(n_1762),
.B(n_1638),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1834),
.A2(n_1681),
.B1(n_1767),
.B2(n_1644),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1846),
.A2(n_1776),
.B(n_1590),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1852),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1681),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1821),
.B(n_1743),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1595),
.B(n_1663),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_1852),
.Y(n_2089)
);

OAI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_1744),
.A2(n_1695),
.B(n_1661),
.Y(n_2090)
);

OA21x2_ASAP7_75t_L g2091 ( 
.A1(n_1865),
.A2(n_1881),
.B(n_1731),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1865),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1580),
.Y(n_2093)
);

AO21x2_ASAP7_75t_L g2094 ( 
.A1(n_1881),
.A2(n_1731),
.B(n_1870),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_1577),
.Y(n_2095)
);

BUFx4_ASAP7_75t_SL g2096 ( 
.A(n_1755),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1580),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_1628),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1673),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_1865),
.A2(n_1881),
.B(n_1578),
.Y(n_2100)
);

NAND2x1p5_ASAP7_75t_L g2101 ( 
.A(n_1628),
.B(n_1340),
.Y(n_2101)
);

OA21x2_ASAP7_75t_L g2102 ( 
.A1(n_1865),
.A2(n_1881),
.B(n_1731),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1580),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1880),
.Y(n_2104)
);

BUFx10_ASAP7_75t_L g2105 ( 
.A(n_1785),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1673),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_1628),
.Y(n_2107)
);

NAND2x1p5_ASAP7_75t_L g2108 ( 
.A(n_1628),
.B(n_1340),
.Y(n_2108)
);

BUFx12f_ASAP7_75t_L g2109 ( 
.A(n_1664),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1862),
.B(n_1497),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1878),
.B(n_1883),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_1628),
.B(n_1340),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_SL g2113 ( 
.A1(n_1880),
.A2(n_1874),
.B(n_1873),
.Y(n_2113)
);

BUFx12f_ASAP7_75t_L g2114 ( 
.A(n_1664),
.Y(n_2114)
);

BUFx2_ASAP7_75t_SL g2115 ( 
.A(n_1628),
.Y(n_2115)
);

INVx6_ASAP7_75t_L g2116 ( 
.A(n_1628),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1628),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_1625),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2007),
.Y(n_2119)
);

BUFx12f_ASAP7_75t_L g2120 ( 
.A(n_2015),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1969),
.A2(n_2089),
.B1(n_1967),
.B2(n_1904),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1907),
.Y(n_2122)
);

OAI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1969),
.A2(n_2062),
.B1(n_2055),
.B2(n_2079),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1907),
.Y(n_2124)
);

OAI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_2055),
.A2(n_2079),
.B1(n_1952),
.B2(n_1919),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_2065),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_SL g2127 ( 
.A1(n_1904),
.A2(n_1954),
.B1(n_2026),
.B2(n_1957),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1953),
.Y(n_2128)
);

OAI21xp33_ASAP7_75t_L g2129 ( 
.A1(n_1940),
.A2(n_1922),
.B(n_1978),
.Y(n_2129)
);

AO21x2_ASAP7_75t_L g2130 ( 
.A1(n_1942),
.A2(n_1921),
.B(n_1887),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1965),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1956),
.Y(n_2132)
);

BUFx2_ASAP7_75t_R g2133 ( 
.A(n_1905),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1886),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1891),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1904),
.B(n_1896),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_2098),
.Y(n_2137)
);

NOR2x1_ASAP7_75t_L g2138 ( 
.A(n_1991),
.B(n_2098),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1944),
.Y(n_2139)
);

INVx4_ASAP7_75t_L g2140 ( 
.A(n_2065),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1908),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_1914),
.A2(n_2090),
.B(n_1975),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1965),
.Y(n_2143)
);

INVx4_ASAP7_75t_L g2144 ( 
.A(n_2065),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_2101),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1912),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_1964),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2020),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_2101),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1952),
.A2(n_2104),
.B1(n_1890),
.B2(n_2079),
.Y(n_2150)
);

BUFx4f_ASAP7_75t_SL g2151 ( 
.A(n_2015),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1890),
.B(n_2104),
.Y(n_2152)
);

CKINVDCx11_ASAP7_75t_R g2153 ( 
.A(n_1909),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1903),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_1937),
.B(n_1987),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1918),
.Y(n_2156)
);

INVx6_ASAP7_75t_L g2157 ( 
.A(n_2105),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1905),
.Y(n_2158)
);

BUFx8_ASAP7_75t_L g2159 ( 
.A(n_2034),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1952),
.A2(n_1940),
.B1(n_1991),
.B2(n_1993),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1948),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1925),
.Y(n_2162)
);

NAND2x1p5_ASAP7_75t_L g2163 ( 
.A(n_1897),
.B(n_1913),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1894),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1926),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_SL g2166 ( 
.A1(n_1954),
.A2(n_1957),
.B1(n_2005),
.B2(n_2113),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2093),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2097),
.Y(n_2168)
);

INVx6_ASAP7_75t_L g2169 ( 
.A(n_2105),
.Y(n_2169)
);

INVx1_ASAP7_75t_SL g2170 ( 
.A(n_1987),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2103),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_SL g2172 ( 
.A(n_1981),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_1924),
.A2(n_2110),
.B1(n_2085),
.B2(n_2061),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2110),
.A2(n_1978),
.B1(n_2021),
.B2(n_1922),
.Y(n_2174)
);

AO21x2_ASAP7_75t_L g2175 ( 
.A1(n_1916),
.A2(n_2100),
.B(n_1900),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_SL g2176 ( 
.A1(n_1997),
.A2(n_1941),
.B(n_2084),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_1915),
.A2(n_1936),
.B(n_1927),
.Y(n_2177)
);

AOI21x1_ASAP7_75t_L g2178 ( 
.A1(n_1950),
.A2(n_2092),
.B(n_1895),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_2000),
.A2(n_2073),
.B1(n_1990),
.B2(n_2083),
.Y(n_2179)
);

INVx6_ASAP7_75t_L g2180 ( 
.A(n_2033),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1959),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1980),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1990),
.A2(n_2083),
.B1(n_2053),
.B2(n_2068),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1984),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1992),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1998),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2044),
.Y(n_2187)
);

BUFx12f_ASAP7_75t_L g2188 ( 
.A(n_2034),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1961),
.B(n_1995),
.Y(n_2189)
);

CKINVDCx11_ASAP7_75t_R g2190 ( 
.A(n_1894),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2022),
.Y(n_2191)
);

INVx6_ASAP7_75t_L g2192 ( 
.A(n_2033),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_2108),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2111),
.B(n_1899),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_2118),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2053),
.A2(n_1994),
.B1(n_2086),
.B2(n_2057),
.Y(n_2196)
);

AOI21x1_ASAP7_75t_L g2197 ( 
.A1(n_1950),
.A2(n_2092),
.B(n_1895),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2027),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2043),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_2118),
.Y(n_2200)
);

AO22x1_ASAP7_75t_L g2201 ( 
.A1(n_2024),
.A2(n_2106),
.B1(n_2099),
.B2(n_1981),
.Y(n_2201)
);

AO21x2_ASAP7_75t_L g2202 ( 
.A1(n_1916),
.A2(n_1900),
.B(n_2094),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2112),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2010),
.Y(n_2204)
);

OR2x6_ASAP7_75t_L g2205 ( 
.A(n_2115),
.B(n_1963),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_1993),
.A2(n_2017),
.B1(n_2042),
.B2(n_2071),
.Y(n_2206)
);

AO21x1_ASAP7_75t_SL g2207 ( 
.A1(n_1893),
.A2(n_1902),
.B(n_1898),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2018),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2080),
.Y(n_2209)
);

OAI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_2078),
.A2(n_2025),
.B(n_2056),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_SL g2211 ( 
.A1(n_2006),
.A2(n_2112),
.B(n_1929),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1897),
.Y(n_2212)
);

BUFx2_ASAP7_75t_R g2213 ( 
.A(n_2099),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1889),
.Y(n_2214)
);

BUFx2_ASAP7_75t_SL g2215 ( 
.A(n_1901),
.Y(n_2215)
);

CKINVDCx11_ASAP7_75t_R g2216 ( 
.A(n_2109),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2096),
.Y(n_2217)
);

BUFx2_ASAP7_75t_R g2218 ( 
.A(n_2106),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1913),
.Y(n_2219)
);

INVx6_ASAP7_75t_L g2220 ( 
.A(n_1945),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_SL g2221 ( 
.A1(n_2024),
.A2(n_2006),
.B1(n_2041),
.B2(n_2008),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2045),
.Y(n_2222)
);

INVx8_ASAP7_75t_L g2223 ( 
.A(n_2109),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_SL g2224 ( 
.A(n_1971),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2117),
.Y(n_2225)
);

BUFx2_ASAP7_75t_L g2226 ( 
.A(n_2117),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2116),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1958),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2037),
.B(n_2058),
.Y(n_2229)
);

OAI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2071),
.A2(n_2042),
.B1(n_2050),
.B2(n_2059),
.Y(n_2230)
);

INVx6_ASAP7_75t_L g2231 ( 
.A(n_1945),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_1999),
.Y(n_2232)
);

BUFx8_ASAP7_75t_SL g2233 ( 
.A(n_2114),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1934),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2087),
.A2(n_2057),
.B1(n_2050),
.B2(n_2059),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1985),
.B(n_1951),
.Y(n_2236)
);

BUFx2_ASAP7_75t_SL g2237 ( 
.A(n_1901),
.Y(n_2237)
);

BUFx3_ASAP7_75t_L g2238 ( 
.A(n_1999),
.Y(n_2238)
);

OAI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2056),
.A2(n_2067),
.B(n_2030),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2041),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1920),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1920),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2039),
.A2(n_2074),
.B1(n_1977),
.B2(n_2071),
.Y(n_2243)
);

CKINVDCx8_ASAP7_75t_R g2244 ( 
.A(n_1979),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2096),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2013),
.A2(n_2082),
.B1(n_2074),
.B2(n_1928),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_2052),
.A2(n_2072),
.B1(n_1995),
.B2(n_2040),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1951),
.B(n_1960),
.Y(n_2248)
);

BUFx2_ASAP7_75t_L g2249 ( 
.A(n_1970),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1939),
.Y(n_2250)
);

BUFx2_ASAP7_75t_L g2251 ( 
.A(n_1970),
.Y(n_2251)
);

BUFx8_ASAP7_75t_SL g2252 ( 
.A(n_2114),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1960),
.B(n_1923),
.Y(n_2253)
);

NAND2x1p5_ASAP7_75t_L g2254 ( 
.A(n_1932),
.B(n_2028),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2116),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2052),
.A2(n_2040),
.B1(n_2036),
.B2(n_1973),
.Y(n_2256)
);

INVx3_ASAP7_75t_SL g2257 ( 
.A(n_2013),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_SL g2258 ( 
.A1(n_2046),
.A2(n_2003),
.B1(n_1931),
.B2(n_1966),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2095),
.B(n_1938),
.Y(n_2259)
);

CKINVDCx20_ASAP7_75t_R g2260 ( 
.A(n_2002),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1930),
.Y(n_2261)
);

INVx6_ASAP7_75t_L g2262 ( 
.A(n_1932),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2028),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2009),
.B(n_1928),
.Y(n_2264)
);

OAI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_2067),
.A2(n_2076),
.B(n_2023),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_1968),
.A2(n_1988),
.B(n_1962),
.Y(n_2266)
);

BUFx2_ASAP7_75t_R g2267 ( 
.A(n_2047),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1906),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_1974),
.Y(n_2269)
);

AOI222xp33_ASAP7_75t_L g2270 ( 
.A1(n_2012),
.A2(n_1982),
.B1(n_1928),
.B2(n_1943),
.C1(n_2047),
.C2(n_2049),
.Y(n_2270)
);

BUFx4f_ASAP7_75t_SL g2271 ( 
.A(n_2012),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2107),
.B(n_2064),
.Y(n_2272)
);

BUFx12f_ASAP7_75t_L g2273 ( 
.A(n_2049),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2136),
.B(n_1961),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2119),
.Y(n_2275)
);

INVxp67_ASAP7_75t_SL g2276 ( 
.A(n_2131),
.Y(n_2276)
);

CKINVDCx16_ASAP7_75t_R g2277 ( 
.A(n_2172),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2121),
.A2(n_2051),
.B1(n_2066),
.B2(n_2088),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_R g2279 ( 
.A(n_2172),
.B(n_1996),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2229),
.B(n_2019),
.Y(n_2280)
);

CKINVDCx16_ASAP7_75t_R g2281 ( 
.A(n_2120),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_2236),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2170),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2134),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2170),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2135),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_R g2287 ( 
.A(n_2151),
.B(n_2004),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_2159),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2228),
.B(n_1955),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2248),
.B(n_1888),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_2159),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_R g2292 ( 
.A(n_2151),
.B(n_2245),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_2126),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2173),
.B(n_1955),
.Y(n_2294)
);

OAI222xp33_ASAP7_75t_L g2295 ( 
.A1(n_2121),
.A2(n_2031),
.B1(n_1982),
.B2(n_1986),
.C1(n_1983),
.C2(n_2011),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2155),
.B(n_2136),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2141),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2129),
.A2(n_2046),
.B1(n_2066),
.B2(n_2081),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2122),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2146),
.Y(n_2300)
);

NAND2x1p5_ASAP7_75t_L g2301 ( 
.A(n_2140),
.B(n_2077),
.Y(n_2301)
);

INVx2_ASAP7_75t_SL g2302 ( 
.A(n_2205),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2123),
.A2(n_2051),
.B1(n_2066),
.B2(n_2031),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2194),
.B(n_1888),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2123),
.A2(n_2011),
.B(n_1983),
.Y(n_2305)
);

CKINVDCx16_ASAP7_75t_R g2306 ( 
.A(n_2188),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2214),
.B(n_1892),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2124),
.Y(n_2308)
);

CKINVDCx16_ASAP7_75t_R g2309 ( 
.A(n_2205),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2128),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_R g2311 ( 
.A(n_2271),
.B(n_1892),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_2153),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2156),
.Y(n_2313)
);

CKINVDCx16_ASAP7_75t_R g2314 ( 
.A(n_2205),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2253),
.B(n_1910),
.Y(n_2315)
);

CKINVDCx20_ASAP7_75t_R g2316 ( 
.A(n_2190),
.Y(n_2316)
);

CKINVDCx20_ASAP7_75t_R g2317 ( 
.A(n_2216),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_2126),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2226),
.Y(n_2319)
);

OAI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2177),
.A2(n_1968),
.B(n_2001),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2125),
.A2(n_2046),
.B1(n_2036),
.B2(n_1973),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2272),
.B(n_1972),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2173),
.B(n_2060),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_2153),
.Y(n_2324)
);

CKINVDCx16_ASAP7_75t_R g2325 ( 
.A(n_2238),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_2216),
.Y(n_2326)
);

CKINVDCx11_ASAP7_75t_R g2327 ( 
.A(n_2244),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2132),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2162),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2179),
.B(n_2060),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2165),
.Y(n_2331)
);

CKINVDCx16_ASAP7_75t_R g2332 ( 
.A(n_2215),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_2233),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2179),
.B(n_2060),
.Y(n_2334)
);

OR2x6_ASAP7_75t_L g2335 ( 
.A(n_2160),
.B(n_2032),
.Y(n_2335)
);

CKINVDCx20_ASAP7_75t_R g2336 ( 
.A(n_2252),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_R g2337 ( 
.A(n_2271),
.B(n_1917),
.Y(n_2337)
);

NAND2xp33_ASAP7_75t_R g2338 ( 
.A(n_2261),
.B(n_1917),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2196),
.B(n_2016),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2167),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2183),
.A2(n_2046),
.B1(n_2016),
.B2(n_2029),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2139),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2196),
.B(n_2035),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2222),
.B(n_2183),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2131),
.Y(n_2345)
);

NAND2x1_ASAP7_75t_L g2346 ( 
.A(n_2138),
.B(n_2176),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_2223),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2143),
.Y(n_2348)
);

OR2x6_ASAP7_75t_L g2349 ( 
.A(n_2160),
.B(n_2077),
.Y(n_2349)
);

BUFx2_ASAP7_75t_L g2350 ( 
.A(n_2145),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_2223),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2148),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2154),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2143),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_2223),
.Y(n_2355)
);

BUFx12f_ASAP7_75t_L g2356 ( 
.A(n_2232),
.Y(n_2356)
);

NAND2xp33_ASAP7_75t_R g2357 ( 
.A(n_2158),
.B(n_1930),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2168),
.Y(n_2358)
);

AOI22xp33_ASAP7_75t_L g2359 ( 
.A1(n_2125),
.A2(n_2046),
.B1(n_2029),
.B2(n_1976),
.Y(n_2359)
);

CKINVDCx6p67_ASAP7_75t_R g2360 ( 
.A(n_2232),
.Y(n_2360)
);

NOR3xp33_ASAP7_75t_SL g2361 ( 
.A(n_2211),
.B(n_1972),
.C(n_1976),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2126),
.Y(n_2362)
);

CKINVDCx16_ASAP7_75t_R g2363 ( 
.A(n_2237),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2249),
.B(n_1972),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2251),
.B(n_2063),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_2212),
.Y(n_2366)
);

AND2x4_ASAP7_75t_SL g2367 ( 
.A(n_2140),
.B(n_2144),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2273),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2259),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_2133),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2161),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2189),
.A2(n_1947),
.B(n_1933),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2181),
.Y(n_2373)
);

CKINVDCx20_ASAP7_75t_R g2374 ( 
.A(n_2260),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2149),
.Y(n_2375)
);

CKINVDCx16_ASAP7_75t_R g2376 ( 
.A(n_2217),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2133),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_2213),
.Y(n_2378)
);

OAI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2166),
.A2(n_2174),
.B1(n_2127),
.B2(n_2206),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2184),
.Y(n_2380)
);

OAI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2206),
.A2(n_2070),
.B1(n_2054),
.B2(n_2048),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2235),
.B(n_2054),
.Y(n_2382)
);

AOI22xp33_ASAP7_75t_L g2383 ( 
.A1(n_2166),
.A2(n_1949),
.B1(n_1935),
.B2(n_1911),
.Y(n_2383)
);

INVx2_ASAP7_75t_SL g2384 ( 
.A(n_2157),
.Y(n_2384)
);

NOR2x1_ASAP7_75t_SL g2385 ( 
.A(n_2207),
.B(n_2069),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2157),
.Y(n_2386)
);

INVxp67_ASAP7_75t_L g2387 ( 
.A(n_2263),
.Y(n_2387)
);

CKINVDCx8_ASAP7_75t_R g2388 ( 
.A(n_2213),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_R g2389 ( 
.A(n_2144),
.B(n_2048),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2147),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2171),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2218),
.Y(n_2392)
);

A2O1A1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2211),
.A2(n_2038),
.B(n_2014),
.C(n_1962),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2174),
.A2(n_2070),
.B1(n_2102),
.B2(n_2091),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_R g2395 ( 
.A(n_2180),
.B(n_2075),
.Y(n_2395)
);

OR2x4_ASAP7_75t_L g2396 ( 
.A(n_2241),
.B(n_1989),
.Y(n_2396)
);

CKINVDCx16_ASAP7_75t_R g2397 ( 
.A(n_2164),
.Y(n_2397)
);

AOI22xp33_ASAP7_75t_L g2398 ( 
.A1(n_2127),
.A2(n_1949),
.B1(n_1946),
.B2(n_2038),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2274),
.B(n_2130),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2296),
.B(n_2152),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2344),
.B(n_2182),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2275),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2274),
.B(n_2130),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2339),
.B(n_2256),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2341),
.B(n_2256),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2335),
.B(n_2265),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2283),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2284),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2341),
.B(n_2239),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2286),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2345),
.B(n_2150),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2379),
.A2(n_2270),
.B1(n_2150),
.B2(n_2230),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2297),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2300),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2299),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2313),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2308),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2329),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2310),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_2335),
.B(n_2265),
.Y(n_2420)
);

INVx2_ASAP7_75t_SL g2421 ( 
.A(n_2396),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2331),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2340),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2353),
.B(n_2185),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2335),
.B(n_2239),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2348),
.B(n_2247),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2285),
.B(n_2247),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2379),
.A2(n_2270),
.B1(n_2230),
.B2(n_2243),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2358),
.Y(n_2429)
);

OR2x2_ASAP7_75t_L g2430 ( 
.A(n_2354),
.B(n_2276),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2391),
.Y(n_2431)
);

AOI221xp5_ASAP7_75t_L g2432 ( 
.A1(n_2303),
.A2(n_2243),
.B1(n_2234),
.B2(n_2209),
.C(n_2204),
.Y(n_2432)
);

HB1xp67_ASAP7_75t_L g2433 ( 
.A(n_2319),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2369),
.B(n_2142),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2371),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2373),
.B(n_2186),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2320),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2328),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2390),
.Y(n_2439)
);

NOR2x1_ASAP7_75t_L g2440 ( 
.A(n_2305),
.B(n_2137),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2380),
.B(n_2142),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2342),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2352),
.Y(n_2443)
);

OR2x2_ASAP7_75t_L g2444 ( 
.A(n_2282),
.B(n_2246),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2323),
.B(n_2330),
.Y(n_2445)
);

OAI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2305),
.A2(n_2221),
.B(n_2258),
.C(n_2264),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2278),
.B(n_2210),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2397),
.B(n_2195),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2349),
.Y(n_2449)
);

INVxp33_ASAP7_75t_L g2450 ( 
.A(n_2395),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_2334),
.B(n_2187),
.Y(n_2451)
);

INVx1_ASAP7_75t_SL g2452 ( 
.A(n_2376),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2278),
.B(n_2394),
.Y(n_2453)
);

CKINVDCx20_ASAP7_75t_R g2454 ( 
.A(n_2374),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2350),
.Y(n_2455)
);

AOI21xp5_ASAP7_75t_SL g2456 ( 
.A1(n_2385),
.A2(n_2242),
.B(n_2250),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2307),
.B(n_2191),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2289),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2396),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2394),
.B(n_2202),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2343),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2359),
.B(n_2202),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2375),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2294),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_L g2465 ( 
.A(n_2309),
.B(n_2200),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2315),
.B(n_2198),
.Y(n_2466)
);

OR2x2_ASAP7_75t_L g2467 ( 
.A(n_2366),
.B(n_2147),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2303),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2290),
.B(n_2199),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2349),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2453),
.B(n_2298),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2458),
.B(n_2387),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_2449),
.B(n_2361),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2453),
.B(n_2321),
.Y(n_2474)
);

BUFx2_ASAP7_75t_SL g2475 ( 
.A(n_2421),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2451),
.B(n_2382),
.Y(n_2476)
);

HB1xp67_ASAP7_75t_L g2477 ( 
.A(n_2433),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2451),
.B(n_2365),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2449),
.B(n_2470),
.Y(n_2479)
);

OR2x2_ASAP7_75t_L g2480 ( 
.A(n_2434),
.B(n_2314),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2438),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2399),
.B(n_2175),
.Y(n_2482)
);

NAND2x1p5_ASAP7_75t_L g2483 ( 
.A(n_2440),
.B(n_2302),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2439),
.B(n_2280),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2400),
.B(n_2364),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2407),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2415),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2415),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2399),
.B(n_2175),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2449),
.B(n_2266),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2403),
.B(n_2178),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2417),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2417),
.Y(n_2493)
);

INVxp67_ASAP7_75t_SL g2494 ( 
.A(n_2430),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2403),
.B(n_2197),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2419),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2400),
.B(n_2264),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2464),
.B(n_2372),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2430),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2421),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2445),
.B(n_2208),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2435),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2450),
.B(n_2277),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2442),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2437),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2443),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2499),
.B(n_2464),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2487),
.Y(n_2508)
);

INVxp67_ASAP7_75t_SL g2509 ( 
.A(n_2477),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2494),
.B(n_2434),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2487),
.Y(n_2511)
);

OR2x2_ASAP7_75t_L g2512 ( 
.A(n_2482),
.B(n_2445),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2482),
.B(n_2447),
.Y(n_2513)
);

NOR2x1p5_ASAP7_75t_L g2514 ( 
.A(n_2473),
.B(n_2470),
.Y(n_2514)
);

BUFx2_ASAP7_75t_L g2515 ( 
.A(n_2500),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2492),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2489),
.B(n_2426),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2488),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2474),
.B(n_2427),
.Y(n_2519)
);

NOR2xp67_ASAP7_75t_L g2520 ( 
.A(n_2473),
.B(n_2378),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2486),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2489),
.B(n_2447),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2488),
.Y(n_2523)
);

INVxp67_ASAP7_75t_L g2524 ( 
.A(n_2480),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2474),
.B(n_2427),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2471),
.B(n_2468),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2493),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2471),
.B(n_2468),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2476),
.B(n_2404),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2490),
.B(n_2470),
.Y(n_2530)
);

OAI221xp5_ASAP7_75t_L g2531 ( 
.A1(n_2480),
.A2(n_2428),
.B1(n_2412),
.B2(n_2446),
.C(n_2483),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2493),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2492),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2478),
.B(n_2426),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2485),
.B(n_2461),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2483),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2491),
.B(n_2404),
.Y(n_2537)
);

OAI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2483),
.A2(n_2456),
.B(n_2450),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2491),
.B(n_2460),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2496),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2496),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2495),
.B(n_2460),
.Y(n_2542)
);

OR2x2_ASAP7_75t_L g2543 ( 
.A(n_2517),
.B(n_2497),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2526),
.B(n_2495),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2517),
.B(n_2501),
.Y(n_2545)
);

OAI32xp33_ASAP7_75t_L g2546 ( 
.A1(n_2538),
.A2(n_2452),
.A3(n_2363),
.B1(n_2332),
.B2(n_2463),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2512),
.B(n_2484),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2521),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2515),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2526),
.B(n_2498),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2528),
.B(n_2513),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2515),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2512),
.B(n_2472),
.Y(n_2553)
);

AOI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2531),
.A2(n_2503),
.B1(n_2473),
.B2(n_2479),
.Y(n_2554)
);

NAND4xp75_ASAP7_75t_L g2555 ( 
.A(n_2520),
.B(n_2465),
.C(n_2448),
.D(n_2432),
.Y(n_2555)
);

NAND2x2_ASAP7_75t_L g2556 ( 
.A(n_2514),
.B(n_2388),
.Y(n_2556)
);

OAI21xp33_ASAP7_75t_L g2557 ( 
.A1(n_2528),
.A2(n_2473),
.B(n_2498),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2536),
.B(n_2500),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2524),
.A2(n_2444),
.B1(n_2338),
.B2(n_2455),
.Y(n_2559)
);

OAI22xp33_ASAP7_75t_L g2560 ( 
.A1(n_2536),
.A2(n_2459),
.B1(n_2444),
.B2(n_2411),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2509),
.A2(n_2405),
.B1(n_2360),
.B2(n_2401),
.Y(n_2561)
);

AOI32xp33_ASAP7_75t_L g2562 ( 
.A1(n_2536),
.A2(n_2479),
.A3(n_2367),
.B1(n_2381),
.B2(n_2258),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2516),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2510),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2510),
.Y(n_2565)
);

NOR4xp25_ASAP7_75t_L g2566 ( 
.A(n_2507),
.B(n_2295),
.C(n_2408),
.D(n_2402),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2537),
.B(n_2479),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2535),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2513),
.A2(n_2479),
.B1(n_2405),
.B2(n_2425),
.Y(n_2569)
);

OAI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2514),
.A2(n_2475),
.B1(n_2456),
.B2(n_2454),
.Y(n_2570)
);

OAI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_2519),
.A2(n_2459),
.B1(n_2411),
.B2(n_2346),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2516),
.Y(n_2572)
);

OAI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2535),
.A2(n_2475),
.B1(n_2454),
.B2(n_2392),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2522),
.A2(n_2469),
.B1(n_2466),
.B2(n_2377),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2534),
.B(n_2537),
.Y(n_2575)
);

OAI33xp33_ASAP7_75t_L g2576 ( 
.A1(n_2529),
.A2(n_2370),
.A3(n_2457),
.B1(n_2431),
.B2(n_2429),
.B3(n_2423),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2568),
.B(n_2564),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2573),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2565),
.Y(n_2579)
);

NAND4xp25_ASAP7_75t_SL g2580 ( 
.A(n_2562),
.B(n_2317),
.C(n_2336),
.D(n_2316),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2575),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2550),
.Y(n_2582)
);

A2O1A1Ixp33_ASAP7_75t_L g2583 ( 
.A1(n_2554),
.A2(n_2546),
.B(n_2559),
.C(n_2557),
.Y(n_2583)
);

OAI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2559),
.A2(n_2525),
.B1(n_2534),
.B2(n_2522),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2543),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2545),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2548),
.Y(n_2587)
);

AOI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2566),
.A2(n_2542),
.B1(n_2539),
.B2(n_2530),
.C(n_2410),
.Y(n_2588)
);

AOI221xp5_ASAP7_75t_L g2589 ( 
.A1(n_2576),
.A2(n_2542),
.B1(n_2539),
.B2(n_2530),
.C(n_2422),
.Y(n_2589)
);

AOI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2555),
.A2(n_2530),
.B1(n_2409),
.B2(n_2420),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2547),
.Y(n_2591)
);

OAI31xp33_ASAP7_75t_L g2592 ( 
.A1(n_2570),
.A2(n_2530),
.A3(n_2420),
.B(n_2406),
.Y(n_2592)
);

OAI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2561),
.A2(n_2558),
.B(n_2549),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2551),
.B(n_2508),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2553),
.Y(n_2595)
);

OAI21xp33_ASAP7_75t_L g2596 ( 
.A1(n_2569),
.A2(n_2574),
.B(n_2561),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2578),
.B(n_2567),
.Y(n_2597)
);

INVxp67_ASAP7_75t_L g2598 ( 
.A(n_2580),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2577),
.B(n_2544),
.Y(n_2599)
);

OAI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2583),
.A2(n_2556),
.B1(n_2574),
.B2(n_2571),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2593),
.B(n_2552),
.Y(n_2601)
);

AOI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2588),
.A2(n_2560),
.B1(n_2414),
.B2(n_2413),
.C(n_2416),
.Y(n_2602)
);

INVx2_ASAP7_75t_SL g2603 ( 
.A(n_2585),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2577),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2581),
.Y(n_2605)
);

OAI21xp33_ASAP7_75t_SL g2606 ( 
.A1(n_2592),
.A2(n_2572),
.B(n_2563),
.Y(n_2606)
);

AOI321xp33_ASAP7_75t_L g2607 ( 
.A1(n_2596),
.A2(n_2409),
.A3(n_2462),
.B1(n_2425),
.B2(n_2420),
.C(n_2406),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2582),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2584),
.A2(n_2587),
.B(n_2589),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2579),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2595),
.B(n_2586),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2594),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2590),
.B(n_2508),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2591),
.B(n_2502),
.Y(n_2614)
);

AOI22xp33_ASAP7_75t_L g2615 ( 
.A1(n_2578),
.A2(n_2304),
.B1(n_2337),
.B2(n_2322),
.Y(n_2615)
);

AOI221xp5_ASAP7_75t_L g2616 ( 
.A1(n_2578),
.A2(n_2418),
.B1(n_2201),
.B2(n_2532),
.C(n_2527),
.Y(n_2616)
);

OAI221xp5_ASAP7_75t_SL g2617 ( 
.A1(n_2578),
.A2(n_2221),
.B1(n_2383),
.B2(n_2398),
.C(n_2393),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2579),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2596),
.A2(n_2406),
.B1(n_2425),
.B2(n_2490),
.Y(n_2619)
);

OAI221xp5_ASAP7_75t_L g2620 ( 
.A1(n_2583),
.A2(n_2357),
.B1(n_2326),
.B2(n_2324),
.C(n_2312),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2603),
.Y(n_2621)
);

AND3x1_ASAP7_75t_L g2622 ( 
.A(n_2616),
.B(n_2306),
.C(n_2281),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_SL g2623 ( 
.A1(n_2598),
.A2(n_2301),
.B(n_2218),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_SL g2624 ( 
.A(n_2620),
.B(n_2267),
.Y(n_2624)
);

BUFx2_ASAP7_75t_L g2625 ( 
.A(n_2598),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2611),
.Y(n_2626)
);

NOR3x1_ASAP7_75t_L g2627 ( 
.A(n_2600),
.B(n_2327),
.C(n_2384),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2609),
.B(n_2502),
.Y(n_2628)
);

NOR3x1_ASAP7_75t_L g2629 ( 
.A(n_2604),
.B(n_2386),
.C(n_2291),
.Y(n_2629)
);

O2A1O1Ixp5_ASAP7_75t_L g2630 ( 
.A1(n_2617),
.A2(n_2505),
.B(n_2504),
.C(n_2506),
.Y(n_2630)
);

AOI211xp5_ASAP7_75t_L g2631 ( 
.A1(n_2617),
.A2(n_2287),
.B(n_2279),
.C(n_2257),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2601),
.A2(n_2325),
.B1(n_2490),
.B2(n_2462),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2597),
.B(n_2504),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2614),
.Y(n_2634)
);

AOI221xp5_ASAP7_75t_L g2635 ( 
.A1(n_2606),
.A2(n_2541),
.B1(n_2540),
.B2(n_2511),
.C(n_2518),
.Y(n_2635)
);

OR2x2_ASAP7_75t_L g2636 ( 
.A(n_2605),
.B(n_2511),
.Y(n_2636)
);

INVx2_ASAP7_75t_SL g2637 ( 
.A(n_2608),
.Y(n_2637)
);

OAI21xp33_ASAP7_75t_SL g2638 ( 
.A1(n_2602),
.A2(n_2506),
.B(n_2518),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2631),
.A2(n_2619),
.B1(n_2615),
.B2(n_2613),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2633),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2626),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2622),
.A2(n_2615),
.B1(n_2599),
.B2(n_2612),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2631),
.A2(n_2613),
.B1(n_2618),
.B2(n_2610),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2637),
.Y(n_2644)
);

OAI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2625),
.A2(n_2613),
.B(n_2610),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2634),
.B(n_2618),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2621),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2623),
.A2(n_2288),
.B(n_2347),
.Y(n_2648)
);

AOI211x1_ASAP7_75t_L g2649 ( 
.A1(n_2628),
.A2(n_2607),
.B(n_2268),
.C(n_2240),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2636),
.Y(n_2650)
);

NOR2xp67_ASAP7_75t_L g2651 ( 
.A(n_2638),
.B(n_2333),
.Y(n_2651)
);

OAI21xp33_ASAP7_75t_SL g2652 ( 
.A1(n_2635),
.A2(n_2137),
.B(n_2541),
.Y(n_2652)
);

AOI211xp5_ASAP7_75t_L g2653 ( 
.A1(n_2624),
.A2(n_2292),
.B(n_2257),
.C(n_2351),
.Y(n_2653)
);

AOI221xp5_ASAP7_75t_L g2654 ( 
.A1(n_2644),
.A2(n_2622),
.B1(n_2630),
.B2(n_2627),
.C(n_2632),
.Y(n_2654)
);

A2O1A1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2651),
.A2(n_2355),
.B(n_2629),
.C(n_2368),
.Y(n_2655)
);

OAI211xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2647),
.A2(n_2267),
.B(n_2227),
.C(n_2255),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2641),
.B(n_2523),
.Y(n_2657)
);

NAND4xp25_ASAP7_75t_L g2658 ( 
.A(n_2653),
.B(n_2293),
.C(n_2269),
.D(n_2356),
.Y(n_2658)
);

OAI211xp5_ASAP7_75t_L g2659 ( 
.A1(n_2649),
.A2(n_2311),
.B(n_2389),
.C(n_2362),
.Y(n_2659)
);

OAI21xp33_ASAP7_75t_L g2660 ( 
.A1(n_2639),
.A2(n_2490),
.B(n_2505),
.Y(n_2660)
);

NAND4xp75_ASAP7_75t_L g2661 ( 
.A(n_2645),
.B(n_2224),
.C(n_2157),
.D(n_2169),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2646),
.Y(n_2662)
);

AOI221xp5_ASAP7_75t_L g2663 ( 
.A1(n_2642),
.A2(n_2424),
.B1(n_2436),
.B2(n_2540),
.C(n_2523),
.Y(n_2663)
);

AOI221xp5_ASAP7_75t_L g2664 ( 
.A1(n_2640),
.A2(n_2532),
.B1(n_2527),
.B2(n_2224),
.C(n_2481),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_SL g2665 ( 
.A1(n_2648),
.A2(n_2301),
.B(n_2254),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2650),
.A2(n_2505),
.B1(n_2441),
.B2(n_2461),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2662),
.B(n_2643),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2657),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2660),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2661),
.Y(n_2670)
);

A2O1A1Ixp33_ASAP7_75t_SL g2671 ( 
.A1(n_2665),
.A2(n_2652),
.B(n_2227),
.C(n_2255),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2654),
.A2(n_2169),
.B1(n_2231),
.B2(n_2220),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2655),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_2658),
.Y(n_2674)
);

OR2x2_ASAP7_75t_L g2675 ( 
.A(n_2666),
.B(n_2467),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2663),
.B(n_2533),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_2670),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2669),
.B(n_2664),
.Y(n_2678)
);

NOR3xp33_ASAP7_75t_L g2679 ( 
.A(n_2673),
.B(n_2656),
.C(n_2659),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2674),
.A2(n_2169),
.B1(n_2231),
.B2(n_2220),
.Y(n_2680)
);

NOR3xp33_ASAP7_75t_SL g2681 ( 
.A(n_2668),
.B(n_2231),
.C(n_2220),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2667),
.B(n_2533),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2676),
.Y(n_2683)
);

OAI221xp5_ASAP7_75t_L g2684 ( 
.A1(n_2672),
.A2(n_2262),
.B1(n_2254),
.B2(n_2180),
.C(n_2192),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2675),
.B(n_2671),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_L g2686 ( 
.A(n_2679),
.B(n_2193),
.C(n_2203),
.D(n_2212),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2677),
.Y(n_2687)
);

INVxp67_ASAP7_75t_L g2688 ( 
.A(n_2678),
.Y(n_2688)
);

INVxp33_ASAP7_75t_SL g2689 ( 
.A(n_2680),
.Y(n_2689)
);

INVx1_ASAP7_75t_SL g2690 ( 
.A(n_2687),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2688),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2689),
.Y(n_2692)
);

NOR2xp67_ASAP7_75t_L g2693 ( 
.A(n_2686),
.B(n_2682),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2687),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_2694),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2690),
.A2(n_2683),
.B1(n_2685),
.B2(n_2681),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2692),
.Y(n_2697)
);

OAI31xp33_ASAP7_75t_L g2698 ( 
.A1(n_2697),
.A2(n_2691),
.A3(n_2684),
.B(n_2693),
.Y(n_2698)
);

OAI22x1_ASAP7_75t_L g2699 ( 
.A1(n_2696),
.A2(n_2695),
.B1(n_2163),
.B2(n_2203),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2695),
.Y(n_2700)
);

NOR2x1p5_ASAP7_75t_L g2701 ( 
.A(n_2700),
.B(n_2219),
.Y(n_2701)
);

AOI21xp5_ASAP7_75t_L g2702 ( 
.A1(n_2701),
.A2(n_2698),
.B(n_2699),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_SL g2703 ( 
.A1(n_2702),
.A2(n_2362),
.B1(n_2318),
.B2(n_2225),
.Y(n_2703)
);

OR2x6_ASAP7_75t_L g2704 ( 
.A(n_2703),
.B(n_2262),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2704),
.A2(n_2362),
.B1(n_2318),
.B2(n_2262),
.Y(n_2705)
);


endmodule