module fake_jpeg_2398_n_462 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_462);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_462;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_53),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_26),
.Y(n_128)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_71),
.Y(n_123)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_1),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_83),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_36),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_76),
.Y(n_155)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_26),
.B1(n_19),
.B2(n_39),
.Y(n_127)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_50),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_101),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

CKINVDCx6p67_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_28),
.C(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_34),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_57),
.B(n_28),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_33),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_33),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_50),
.B1(n_49),
.B2(n_32),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_56),
.B1(n_95),
.B2(n_77),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_35),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_136),
.B1(n_153),
.B2(n_39),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_134),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_50),
.B1(n_49),
.B2(n_32),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_49),
.B1(n_42),
.B2(n_40),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_20),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_30),
.Y(n_198)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_166),
.B(n_169),
.Y(n_220)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_168),
.A2(n_180),
.B1(n_121),
.B2(n_136),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_170),
.Y(n_219)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_172),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g224 ( 
.A(n_175),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_176),
.A2(n_198),
.B(n_204),
.Y(n_239)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_109),
.A2(n_85),
.B1(n_78),
.B2(n_67),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_124),
.A2(n_35),
.B1(n_44),
.B2(n_19),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_195),
.B1(n_199),
.B2(n_205),
.Y(n_231)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_34),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_192),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_105),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_197),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_130),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_201),
.Y(n_217)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_203),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_115),
.B(n_30),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_207),
.B1(n_108),
.B2(n_162),
.Y(n_246)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_124),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_134),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_174),
.B(n_163),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_192),
.B(n_187),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_153),
.B1(n_119),
.B2(n_118),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_87),
.B1(n_170),
.B2(n_177),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_159),
.C(n_111),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_227),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_123),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_123),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_213),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_193),
.B1(n_167),
.B2(n_165),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_179),
.A2(n_156),
.B1(n_161),
.B2(n_120),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_29),
.B(n_27),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_114),
.C(n_106),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_173),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_246),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_142),
.B1(n_125),
.B2(n_143),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_247),
.A2(n_248),
.B1(n_266),
.B2(n_219),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_250),
.B(n_251),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_253),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_265),
.B(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_196),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_261),
.B1(n_268),
.B2(n_244),
.Y(n_277)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_262),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_213),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_210),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_187),
.B(n_195),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_222),
.B(n_219),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_264),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_197),
.B(n_202),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_104),
.B1(n_110),
.B2(n_113),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_29),
.B1(n_24),
.B2(n_194),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_191),
.B(n_206),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_223),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_276),
.B1(n_243),
.B2(n_240),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_199),
.B(n_164),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_212),
.B(n_235),
.Y(n_297)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_264),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_262),
.A2(n_255),
.B(n_247),
.C(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_288),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_284),
.A2(n_295),
.B1(n_296),
.B2(n_302),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_257),
.A2(n_217),
.B1(n_220),
.B2(n_240),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_221),
.C(n_217),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_239),
.C(n_211),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_245),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_212),
.C(n_235),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_253),
.C(n_270),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_222),
.B1(n_225),
.B2(n_243),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_256),
.A2(n_250),
.B1(n_251),
.B2(n_275),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_297),
.A2(n_299),
.B(n_258),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_267),
.B1(n_259),
.B2(n_271),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_248),
.A2(n_203),
.B1(n_185),
.B2(n_157),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_310),
.B1(n_311),
.B2(n_315),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_309),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_329),
.C(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_265),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_318),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_263),
.B(n_249),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_313),
.A2(n_323),
.B(n_324),
.Y(n_334)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_319),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_252),
.B1(n_276),
.B2(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_215),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_325),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_215),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_292),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_283),
.A2(n_297),
.B(n_300),
.Y(n_323)
);

NOR2x1_ASAP7_75t_SL g324 ( 
.A(n_291),
.B(n_283),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_281),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_326),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_278),
.B(n_282),
.Y(n_345)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

AOI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_218),
.B(n_279),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_274),
.C(n_218),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_303),
.B1(n_288),
.B2(n_278),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_330),
.A2(n_341),
.B1(n_68),
.B2(n_58),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_344),
.C(n_353),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_304),
.B(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_335),
.B(n_230),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_280),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_339),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_280),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_354),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_278),
.B1(n_301),
.B2(n_302),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_323),
.A2(n_313),
.B(n_324),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_343),
.A2(n_207),
.B(n_100),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_282),
.C(n_278),
.Y(n_344)
);

XOR2x1_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_348),
.Y(n_359)
);

AOI21xp33_ASAP7_75t_L g356 ( 
.A1(n_346),
.A2(n_326),
.B(n_319),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_308),
.C(n_320),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_347),
.B(n_344),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_279),
.B(n_234),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_316),
.A2(n_276),
.B1(n_252),
.B2(n_241),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_97),
.B1(n_96),
.B2(n_92),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_216),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_234),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_216),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_61),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_339),
.B(n_314),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_360),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_350),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_361),
.B(n_362),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_352),
.Y(n_363)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_367),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_368),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g369 ( 
.A(n_331),
.B(n_230),
.CI(n_93),
.CON(n_369),
.SN(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_141),
.B1(n_140),
.B2(n_152),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_152),
.B1(n_141),
.B2(n_140),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_338),
.B(n_2),
.CI(n_3),
.CON(n_372),
.SN(n_372)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_372),
.A2(n_373),
.B1(n_333),
.B2(n_341),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_348),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_375),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_80),
.C(n_70),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_377),
.C(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_378),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_366),
.Y(n_400)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_375),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_371),
.A2(n_330),
.B1(n_334),
.B2(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_392),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_335),
.C(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_394),
.A2(n_381),
.B1(n_380),
.B2(n_359),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_334),
.C(n_354),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_396),
.B(n_376),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_360),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_400),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_366),
.C(n_358),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_405),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_408),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_402),
.A2(n_395),
.B(n_390),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_365),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_409),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_389),
.B(n_365),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_386),
.A2(n_342),
.B1(n_372),
.B2(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_407),
.B(n_410),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_355),
.B(n_377),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_53),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_42),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_42),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_384),
.C(n_387),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_412),
.B(n_423),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_418),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_38),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_391),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_381),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_422),
.Y(n_432)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_411),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_399),
.B(n_382),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_408),
.A2(n_393),
.B(n_383),
.Y(n_424)
);

OAI21x1_ASAP7_75t_SL g428 ( 
.A1(n_424),
.A2(n_420),
.B(n_421),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_410),
.A2(n_383),
.B1(n_388),
.B2(n_40),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_38),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_400),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_429),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_434),
.B1(n_437),
.B2(n_415),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_409),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_420),
.A2(n_403),
.B(n_398),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_431),
.B(n_6),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_40),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_435),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_38),
.Y(n_435)
);

INVx11_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_440),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_417),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_442),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_417),
.C(n_32),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_4),
.C(n_5),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_446),
.B(n_7),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_8),
.Y(n_452)
);

A2O1A1O1Ixp25_ASAP7_75t_L g447 ( 
.A1(n_438),
.A2(n_437),
.B(n_439),
.C(n_443),
.D(n_445),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_447),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_439),
.A2(n_433),
.B(n_8),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_448),
.B(n_449),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_452),
.B(n_9),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_9),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_455),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_456),
.A2(n_451),
.B(n_10),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_458),
.A2(n_454),
.B(n_453),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_459),
.A2(n_457),
.B(n_10),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_9),
.C(n_11),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_12),
.Y(n_462)
);


endmodule