module fake_ariane_2146_n_58 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_58);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_58;

wire n_56;
wire n_24;
wire n_22;
wire n_43;
wire n_49;
wire n_27;
wire n_20;
wire n_48;
wire n_29;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_47;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_51;
wire n_45;
wire n_34;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_39;
wire n_40;
wire n_31;
wire n_42;
wire n_57;
wire n_53;
wire n_21;
wire n_23;
wire n_35;
wire n_54;
wire n_25;

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

OAI22x1_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_10),
.B1(n_7),
.B2(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_15),
.B1(n_11),
.B2(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_36),
.B(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_34),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_26),
.B(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_47),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_49),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OR2x6_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_48),
.Y(n_58)
);


endmodule