module real_jpeg_25791_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_39),
.B1(n_47),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_43),
.B1(n_60),
.B2(n_100),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_60),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_47),
.B(n_53),
.C(n_117),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_2),
.A2(n_39),
.B1(n_42),
.B2(n_47),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_26),
.C(n_87),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_70),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_79),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_39),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_39),
.B1(n_47),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_9),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_81),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_81),
.Y(n_153)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_14),
.A2(n_24),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_123),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_103),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_18),
.B(n_103),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_74),
.B2(n_75),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_48),
.B1(n_72),
.B2(n_73),
.Y(n_20)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_35),
.B2(n_36),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_25),
.A2(n_26),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_25),
.B(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_31),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B(n_41),
.C(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_38),
.B1(n_44),
.B2(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_46),
.C(n_47),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_41),
.A2(n_42),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_42),
.A2(n_51),
.B(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_42),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_42),
.B(n_85),
.Y(n_164)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_64),
.C(n_67),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_55),
.B(n_58),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_52),
.B1(n_86),
.B2(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_59),
.B(n_79),
.Y(n_137)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_62),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_71),
.B(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_70),
.A2(n_153),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_93),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_89),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_85),
.A2(n_89),
.B(n_133),
.Y(n_173)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_111),
.B1(n_113),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B(n_101),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_114),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_105),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_114),
.B1(n_115),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_112),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_112),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_118),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_151),
.B(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_138),
.B(n_183),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.C(n_134),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_177),
.B(n_182),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_167),
.B(n_176),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_154),
.B(n_166),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_149),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_162),
.B(n_165),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_173),
.C(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);


endmodule