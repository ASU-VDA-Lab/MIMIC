module fake_netlist_5_951_n_2794 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_785, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_802, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_753, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_788, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_755, n_6, n_509, n_568, n_39, n_147, n_373, n_757, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_375, n_301, n_779, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_741, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_752, n_331, n_10, n_24, n_406, n_519, n_470, n_782, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_760, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_442, n_157, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_798, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_144, n_114, n_96, n_772, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_236, n_388, n_761, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_770, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_745, n_627, n_767, n_172, n_206, n_217, n_440, n_726, n_478, n_793, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_794, n_768, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_797, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_766, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_799, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_764, n_200, n_162, n_64, n_759, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_747, n_52, n_278, n_784, n_110, n_2794);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_755;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_757;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_375;
input n_301;
input n_779;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_741;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_782;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_144;
input n_114;
input n_96;
input n_772;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_761;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_794;
input n_768;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_797;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_766;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_799;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_162;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_2794;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2561;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_897;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_1600;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_2331;
wire n_2293;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2342;
wire n_1832;
wire n_1851;
wire n_999;
wire n_2046;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2339;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_1159;
wire n_957;
wire n_2124;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2650;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_984;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_1232;
wire n_1603;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_1812;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_2421;
wire n_2286;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2430;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_2687;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2717;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2505;
wire n_2438;
wire n_2427;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_2704;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g803 ( 
.A(n_266),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_463),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_786),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_245),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_762),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_778),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_99),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_466),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_437),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_6),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_286),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_660),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_69),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_729),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_758),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_766),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_586),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_699),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_462),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_300),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_785),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_727),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_395),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_143),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_695),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_383),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_497),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_456),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_159),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_750),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_731),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_693),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_118),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_709),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_208),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_601),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_756),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_748),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_793),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_443),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_356),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_469),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_708),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_234),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_25),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_339),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_85),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_203),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_537),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_234),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_364),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_698),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_91),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_780),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_765),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_638),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_781),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_735),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_393),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_44),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_794),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_640),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_102),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_553),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_226),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_259),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_162),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_333),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_779),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_481),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_774),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_546),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_188),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_214),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_221),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_767),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_261),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_365),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_771),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_757),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_391),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_503),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_388),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_64),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_506),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_61),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_581),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_369),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_120),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_707),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_455),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_717),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_555),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_469),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_763),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_457),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_658),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_473),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_246),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_721),
.Y(n_904)
);

INVx4_ASAP7_75t_R g905 ( 
.A(n_400),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_445),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_715),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_238),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_162),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_351),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_417),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_661),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_612),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_711),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_53),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_776),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_281),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_610),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_716),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_189),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_391),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_499),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_24),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_431),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_420),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_456),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_718),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_634),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_253),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_713),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_247),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_454),
.Y(n_932)
);

BUFx10_ASAP7_75t_L g933 ( 
.A(n_67),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_51),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_796),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_300),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_755),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_492),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_678),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_777),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_381),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_580),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_801),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_136),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_739),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_115),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_468),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_607),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_171),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_106),
.Y(n_950)
);

BUFx10_ASAP7_75t_L g951 ( 
.A(n_618),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_710),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_753),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_215),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_80),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_298),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_599),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_104),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_788),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_760),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_768),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_730),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_462),
.Y(n_963)
);

BUFx10_ASAP7_75t_L g964 ( 
.A(n_434),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_791),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_712),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_792),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_425),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_543),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_338),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_327),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_784),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_384),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_770),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_720),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_782),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_726),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_594),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_432),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_759),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_140),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_800),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_752),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_532),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_633),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_520),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_648),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_301),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_606),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_505),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_516),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_579),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_743),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_403),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_754),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_761),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_121),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_725),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_59),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_723),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_260),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_322),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_772),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_440),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_131),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_798),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_151),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_733),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_161),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_507),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_736),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_379),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_326),
.Y(n_1013)
);

BUFx10_ASAP7_75t_L g1014 ( 
.A(n_539),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_353),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_388),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_458),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_392),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_311),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_253),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_764),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_3),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_642),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_751),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_327),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_728),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_737),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_799),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_49),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_246),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_464),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_416),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_620),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_57),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_697),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_399),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_632),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_96),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_20),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_459),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_269),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_461),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_403),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_355),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_472),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_509),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_742),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_0),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_775),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_94),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_572),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_639),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_347),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_367),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_176),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_465),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_769),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_305),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_288),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_285),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_732),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_113),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_336),
.Y(n_1063)
);

BUFx5_ASAP7_75t_L g1064 ( 
.A(n_371),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_32),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_376),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_475),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_740),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_783),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_714),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_460),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_326),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_552),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_746),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_457),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_239),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_500),
.Y(n_1077)
);

BUFx2_ASAP7_75t_R g1078 ( 
.A(n_156),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_773),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_719),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_460),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_166),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_333),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_789),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_548),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_363),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_795),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_356),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_65),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_444),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_749),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_722),
.Y(n_1092)
);

BUFx5_ASAP7_75t_L g1093 ( 
.A(n_797),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_209),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_432),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_316),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_443),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_106),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_545),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_802),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_140),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_668),
.Y(n_1102)
);

BUFx5_ASAP7_75t_L g1103 ( 
.A(n_576),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_790),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_135),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_747),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_71),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_316),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_467),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_309),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_214),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_421),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_687),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_745),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_267),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_7),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_314),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_386),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_787),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_283),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_738),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_626),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_485),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_285),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_242),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_374),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_744),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_724),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_741),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1064),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1064),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1064),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_855),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_805),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_859),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1064),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_935),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_808),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_817),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_819),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_821),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_834),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_837),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1064),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_840),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_841),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_870),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_846),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_942),
.B(n_1000),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_861),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_865),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_858),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_870),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_873),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_870),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_874),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_876),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_878),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_878),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_883),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_898),
.B(n_0),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_914),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_878),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_981),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_884),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_896),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_981),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_901),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1004),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1004),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_828),
.B(n_2),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_902),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_830),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1040),
.Y(n_1176)
);

INVxp33_ASAP7_75t_SL g1177 ( 
.A(n_925),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_951),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_924),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1040),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_912),
.B(n_2),
.Y(n_1181)
);

AND2x2_ASAP7_75t_SL g1182 ( 
.A(n_1173),
.B(n_1007),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1168),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1168),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1175),
.B(n_984),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1152),
.B(n_1051),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1178),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1147),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1153),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1155),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1158),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1159),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1149),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1130),
.A2(n_839),
.B(n_820),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1134),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1163),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1162),
.B(n_1102),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_SL g1198 ( 
.A(n_1161),
.B(n_1040),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1138),
.B(n_842),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1164),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1139),
.B(n_868),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1140),
.B(n_860),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1165),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1141),
.B(n_1101),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1170),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1171),
.Y(n_1206)
);

AND2x6_ASAP7_75t_L g1207 ( 
.A(n_1131),
.B(n_839),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1172),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1142),
.B(n_886),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1176),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1182),
.A2(n_1177),
.B1(n_1181),
.B2(n_1179),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1199),
.B(n_1143),
.Y(n_1212)
);

AND2x6_ASAP7_75t_L g1213 ( 
.A(n_1204),
.B(n_818),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1188),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1189),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1188),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1205),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1205),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1186),
.A2(n_1179),
.B1(n_1136),
.B2(n_1144),
.Y(n_1219)
);

AND2x2_ASAP7_75t_SL g1220 ( 
.A(n_1193),
.B(n_1108),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1191),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1193),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1202),
.B(n_1145),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1187),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1195),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1208),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1208),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1183),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1192),
.Y(n_1229)
);

AND3x2_ASAP7_75t_L g1230 ( 
.A(n_1185),
.B(n_1053),
.C(n_909),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1190),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1196),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1203),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1183),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1201),
.B(n_1146),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1206),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1197),
.B(n_926),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1200),
.Y(n_1238)
);

INVx8_ASAP7_75t_L g1239 ( 
.A(n_1207),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1207),
.A2(n_1198),
.B1(n_1132),
.B2(n_1054),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_1209),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1210),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1184),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1207),
.B(n_1148),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1184),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_L g1246 ( 
.A(n_1194),
.B(n_853),
.C(n_822),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1188),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1195),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1182),
.A2(n_1151),
.B1(n_1154),
.B2(n_1150),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1199),
.B(n_1156),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1195),
.B(n_963),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1188),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1199),
.B(n_1157),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1189),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1189),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1199),
.B(n_1166),
.C(n_1160),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1235),
.B(n_1212),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1246),
.A2(n_894),
.B1(n_897),
.B2(n_852),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1211),
.A2(n_1106),
.B1(n_1113),
.B2(n_978),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1223),
.B(n_1167),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1243),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1231),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1233),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1250),
.A2(n_1024),
.B1(n_1067),
.B2(n_1011),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1219),
.A2(n_815),
.B1(n_824),
.B2(n_809),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1215),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1253),
.B(n_1169),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1221),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1232),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1256),
.B(n_1174),
.Y(n_1270)
);

O2A1O1Ixp5_ASAP7_75t_L g1271 ( 
.A1(n_1238),
.A2(n_1119),
.B(n_835),
.C(n_857),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1249),
.B(n_1070),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1236),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1254),
.B(n_825),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1255),
.B(n_864),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1228),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1245),
.B(n_875),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1234),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1213),
.B(n_889),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1229),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1213),
.B(n_891),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1224),
.B(n_1220),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1224),
.B(n_1133),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1241),
.A2(n_1073),
.B1(n_1137),
.B2(n_1135),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1244),
.A2(n_916),
.B1(n_918),
.B2(n_904),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1213),
.A2(n_928),
.B1(n_930),
.B2(n_922),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1247),
.B(n_1121),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1216),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1242),
.Y(n_1289)
);

NAND2x1_ASAP7_75t_L g1290 ( 
.A(n_1247),
.B(n_818),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1217),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1222),
.B(n_851),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1240),
.B(n_907),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1239),
.B(n_913),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1239),
.B(n_919),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1225),
.B(n_806),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1237),
.B(n_851),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1218),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1237),
.A2(n_943),
.B1(n_945),
.B2(n_940),
.Y(n_1299)
);

NAND2x1p5_ASAP7_75t_L g1300 ( 
.A(n_1248),
.B(n_1226),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1252),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1227),
.A2(n_937),
.B(n_927),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1214),
.B(n_948),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1214),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1230),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1214),
.B(n_938),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1251),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1251),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1244),
.A2(n_952),
.B(n_939),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1212),
.A2(n_1012),
.B1(n_1098),
.B2(n_862),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1235),
.B(n_953),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1235),
.B(n_957),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1243),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1247),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1211),
.B(n_807),
.C(n_804),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1235),
.B(n_962),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1235),
.B(n_967),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1243),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1235),
.B(n_969),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1243),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_1180),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1247),
.Y(n_1322)
);

BUFx5_ASAP7_75t_L g1323 ( 
.A(n_1243),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1235),
.A2(n_960),
.B1(n_961),
.B2(n_959),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1225),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1243),
.Y(n_1326)
);

AO22x2_ASAP7_75t_L g1327 ( 
.A1(n_1211),
.A2(n_1110),
.B1(n_1078),
.B2(n_810),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1235),
.B(n_974),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1224),
.B(n_915),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1235),
.A2(n_972),
.B1(n_975),
.B2(n_966),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1235),
.B(n_976),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1224),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1243),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1235),
.A2(n_980),
.B1(n_982),
.B2(n_977),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1212),
.B(n_1127),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1212),
.B(n_1128),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1228),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1256),
.B(n_983),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1243),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1235),
.B(n_989),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1243),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1243),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1247),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1224),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1212),
.B(n_985),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1243),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1243),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1235),
.B(n_992),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1235),
.B(n_993),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1235),
.B(n_1003),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1256),
.B(n_986),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_SL g1352 ( 
.A(n_1222),
.B(n_1124),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1228),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1243),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1222),
.B(n_863),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1212),
.B(n_811),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1235),
.B(n_1033),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1237),
.B(n_832),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1224),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1257),
.A2(n_1049),
.B(n_1035),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1329),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1311),
.A2(n_1069),
.B(n_1057),
.Y(n_1362)
);

OAI21xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1312),
.A2(n_1087),
.B(n_1080),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1356),
.B(n_1091),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1316),
.A2(n_1319),
.B(n_1317),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1328),
.A2(n_1114),
.B1(n_1092),
.B2(n_1107),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1331),
.B(n_987),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1274),
.A2(n_827),
.B(n_803),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1340),
.A2(n_899),
.B(n_818),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1348),
.B(n_990),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1357),
.B(n_991),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1260),
.B(n_995),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1359),
.B(n_915),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1309),
.A2(n_998),
.B(n_996),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1267),
.B(n_1006),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1264),
.B(n_941),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1270),
.B(n_1008),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1292),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1335),
.A2(n_965),
.B(n_899),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1320),
.B(n_1010),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1275),
.A2(n_838),
.B(n_831),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1336),
.A2(n_965),
.B(n_899),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_1021),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1332),
.B(n_949),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1293),
.A2(n_1026),
.B(n_1023),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1282),
.B(n_1027),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1342),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1346),
.A2(n_845),
.B(n_844),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1314),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1345),
.A2(n_1318),
.B(n_1313),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1326),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1339),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1347),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1266),
.B(n_1028),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1268),
.B(n_1045),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1344),
.B(n_1047),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1341),
.A2(n_1037),
.B(n_965),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1259),
.A2(n_970),
.B1(n_1022),
.B2(n_956),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_L g1401 ( 
.A(n_1323),
.B(n_1093),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1269),
.B(n_1068),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1278),
.B(n_1074),
.Y(n_1403)
);

BUFx4_ASAP7_75t_SL g1404 ( 
.A(n_1305),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1315),
.A2(n_867),
.B(n_880),
.C(n_833),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1323),
.B(n_1077),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1354),
.A2(n_1084),
.B(n_1037),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1294),
.A2(n_1084),
.B(n_1037),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1325),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1314),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1295),
.A2(n_1084),
.B(n_1079),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1262),
.A2(n_854),
.B(n_847),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1337),
.B(n_1085),
.Y(n_1413)
);

O2A1O1Ixp5_ASAP7_75t_L g1414 ( 
.A1(n_1271),
.A2(n_1082),
.B(n_1056),
.C(n_879),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1263),
.A2(n_1100),
.B(n_1099),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1273),
.A2(n_881),
.B(n_866),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1338),
.A2(n_887),
.B(n_885),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1277),
.A2(n_1052),
.B(n_1046),
.C(n_893),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1321),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1353),
.A2(n_1122),
.B(n_1104),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1285),
.A2(n_1123),
.B(n_1129),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1276),
.A2(n_903),
.B(n_888),
.Y(n_1422)
);

INVx3_ASAP7_75t_SL g1423 ( 
.A(n_1358),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1265),
.A2(n_911),
.B(n_946),
.C(n_944),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1323),
.B(n_1093),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1308),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1351),
.A2(n_973),
.B(n_971),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1280),
.A2(n_997),
.B(n_988),
.Y(n_1428)
);

BUFx8_ASAP7_75t_L g1429 ( 
.A(n_1307),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1323),
.B(n_1093),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1352),
.B(n_951),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1272),
.A2(n_1103),
.B1(n_1093),
.B2(n_1044),
.Y(n_1432)
);

OAI21xp33_ASAP7_75t_L g1433 ( 
.A1(n_1355),
.A2(n_1327),
.B(n_1310),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1324),
.B(n_1093),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1289),
.A2(n_1017),
.B(n_1001),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1283),
.B(n_1014),
.Y(n_1437)
);

AND2x6_ASAP7_75t_L g1438 ( 
.A(n_1297),
.B(n_1291),
.Y(n_1438)
);

NOR3xp33_ASAP7_75t_L g1439 ( 
.A(n_1284),
.B(n_813),
.C(n_812),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1288),
.B(n_1103),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1301),
.A2(n_1019),
.B(n_1018),
.Y(n_1441)
);

A2O1A1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1258),
.A2(n_1030),
.B(n_1032),
.C(n_1029),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1322),
.A2(n_1055),
.B(n_1041),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1298),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1299),
.B(n_1014),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1279),
.A2(n_1081),
.B(n_1066),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1304),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1286),
.A2(n_1281),
.B(n_1306),
.C(n_1287),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1300),
.B(n_1061),
.Y(n_1449)
);

BUFx8_ASAP7_75t_L g1450 ( 
.A(n_1327),
.Y(n_1450)
);

AND2x4_ASAP7_75t_SL g1451 ( 
.A(n_1343),
.B(n_1061),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1303),
.A2(n_1302),
.B(n_1290),
.Y(n_1452)
);

O2A1O1Ixp5_ASAP7_75t_L g1453 ( 
.A1(n_1296),
.A2(n_1088),
.B(n_1105),
.C(n_1097),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1257),
.B(n_1103),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1257),
.A2(n_1115),
.B(n_1112),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1359),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1257),
.A2(n_1118),
.B(n_1117),
.Y(n_1457)
);

NOR3xp33_ASAP7_75t_L g1458 ( 
.A(n_1264),
.B(n_816),
.C(n_814),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1257),
.B(n_1103),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1257),
.A2(n_1125),
.B(n_1120),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1274),
.A2(n_1103),
.B(n_905),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1257),
.B(n_1059),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1257),
.B(n_823),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1257),
.A2(n_1016),
.B(n_908),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1257),
.B(n_826),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1257),
.B(n_1095),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1261),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1257),
.B(n_829),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1359),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1261),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1261),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1359),
.B(n_933),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1257),
.A2(n_1111),
.B(n_1094),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1257),
.B(n_836),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1257),
.A2(n_848),
.B1(n_849),
.B2(n_843),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1257),
.B(n_850),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1257),
.B(n_856),
.Y(n_1477)
);

O2A1O1Ixp5_ASAP7_75t_L g1478 ( 
.A1(n_1309),
.A2(n_964),
.B(n_1015),
.C(n_933),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1257),
.A2(n_1083),
.B(n_1076),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1257),
.A2(n_871),
.B(n_869),
.Y(n_1480)
);

BUFx2_ASAP7_75t_SL g1481 ( 
.A(n_1359),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1359),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1257),
.A2(n_877),
.B1(n_882),
.B2(n_872),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1329),
.Y(n_1484)
);

OAI321xp33_ASAP7_75t_L g1485 ( 
.A1(n_1310),
.A2(n_1015),
.A3(n_1090),
.B1(n_964),
.B2(n_900),
.C(n_892),
.Y(n_1485)
);

OR2x6_ASAP7_75t_SL g1486 ( 
.A(n_1264),
.B(n_921),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1257),
.B(n_890),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1257),
.A2(n_906),
.B(n_895),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1359),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1257),
.A2(n_917),
.B(n_910),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1320),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1261),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1257),
.B(n_920),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1257),
.A2(n_929),
.B(n_931),
.C(n_923),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1257),
.B(n_932),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1257),
.A2(n_936),
.B(n_947),
.C(n_934),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1257),
.B(n_950),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1257),
.A2(n_955),
.B(n_954),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1359),
.B(n_1090),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1257),
.B(n_958),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1257),
.A2(n_979),
.B(n_968),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1359),
.Y(n_1502)
);

BUFx4f_ASAP7_75t_L g1503 ( 
.A(n_1314),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1314),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1314),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1261),
.Y(n_1506)
);

O2A1O1Ixp5_ASAP7_75t_L g1507 ( 
.A1(n_1309),
.A2(n_999),
.B(n_1002),
.C(n_994),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1257),
.A2(n_1009),
.B(n_1013),
.C(n_1005),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1359),
.B(n_1020),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1257),
.A2(n_1031),
.B1(n_1034),
.B2(n_1025),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1257),
.A2(n_1038),
.B(n_1036),
.Y(n_1511)
);

AO22x1_ASAP7_75t_L g1512 ( 
.A1(n_1378),
.A2(n_1042),
.B1(n_1043),
.B2(n_1039),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1482),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1502),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1391),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1371),
.B(n_1048),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1468),
.B(n_1050),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1456),
.B(n_1058),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1365),
.A2(n_471),
.B(n_470),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1455),
.A2(n_1062),
.B(n_1063),
.C(n_1060),
.Y(n_1520)
);

OAI22x1_ASAP7_75t_L g1521 ( 
.A1(n_1462),
.A2(n_1071),
.B1(n_1072),
.B2(n_1065),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1503),
.B(n_474),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1389),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1476),
.B(n_1075),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1401),
.A2(n_477),
.B(n_476),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1395),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1373),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1460),
.A2(n_1366),
.B(n_1466),
.C(n_1360),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1086),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1406),
.A2(n_479),
.B(n_478),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1479),
.A2(n_1096),
.B(n_1109),
.C(n_1089),
.Y(n_1531)
);

CKINVDCx14_ASAP7_75t_R g1532 ( 
.A(n_1409),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1436),
.A2(n_482),
.B(n_480),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1361),
.B(n_1116),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1393),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1469),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1491),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1394),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1392),
.A2(n_484),
.B(n_483),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1364),
.A2(n_1126),
.B(n_4),
.C(n_1),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1489),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1463),
.B(n_1),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1467),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1484),
.B(n_486),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1433),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1470),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1465),
.A2(n_488),
.B1(n_489),
.B2(n_487),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1481),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1492),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1425),
.A2(n_491),
.B(n_490),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1474),
.B(n_493),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1506),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_5),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1373),
.Y(n_1554)
);

NOR3xp33_ASAP7_75t_SL g1555 ( 
.A(n_1485),
.B(n_6),
.C(n_7),
.Y(n_1555)
);

NOR3xp33_ASAP7_75t_L g1556 ( 
.A(n_1400),
.B(n_8),
.C(n_9),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1430),
.A2(n_495),
.B(n_494),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1471),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1410),
.B(n_496),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1374),
.A2(n_501),
.B(n_498),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1391),
.Y(n_1561)
);

OAI22x1_ASAP7_75t_L g1562 ( 
.A1(n_1431),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1391),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1505),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1477),
.B(n_1487),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1427),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1423),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1471),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1495),
.B(n_502),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_11),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1500),
.B(n_12),
.Y(n_1571)
);

OR2x6_ASAP7_75t_SL g1572 ( 
.A(n_1510),
.B(n_13),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1377),
.A2(n_1459),
.B(n_1454),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1386),
.B(n_13),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1447),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1505),
.B(n_14),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1444),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1367),
.A2(n_508),
.B1(n_510),
.B2(n_504),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1412),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1448),
.A2(n_512),
.B(n_511),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1375),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1507),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1416),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1472),
.B(n_15),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1458),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1585)
);

BUFx8_ASAP7_75t_L g1586 ( 
.A(n_1505),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1370),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1444),
.Y(n_1588)
);

XOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_1388),
.B(n_517),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1440),
.A2(n_519),
.B(n_518),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1504),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1372),
.B(n_17),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1390),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1432),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1499),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1452),
.A2(n_522),
.B(n_521),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1419),
.Y(n_1597)
);

O2A1O1Ixp5_ASAP7_75t_L g1598 ( 
.A1(n_1379),
.A2(n_1376),
.B(n_1434),
.C(n_1421),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1457),
.B(n_19),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1494),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1380),
.B(n_1439),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1480),
.B(n_21),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1368),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1445),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1383),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1488),
.B(n_25),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1490),
.B(n_1498),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1496),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1382),
.A2(n_524),
.B1(n_525),
.B2(n_523),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1426),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1398),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1501),
.B(n_26),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1405),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1385),
.A2(n_527),
.B(n_526),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1417),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1396),
.B(n_528),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1438),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1461),
.A2(n_530),
.B(n_529),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1429),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1511),
.B(n_1397),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1478),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_R g1622 ( 
.A(n_1429),
.B(n_531),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1402),
.A2(n_534),
.B(n_533),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1414),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1486),
.B(n_30),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1387),
.A2(n_1483),
.B1(n_1475),
.B2(n_1403),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1413),
.A2(n_536),
.B(n_535),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1381),
.A2(n_540),
.B(n_538),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1508),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1464),
.B(n_33),
.Y(n_1630)
);

AOI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1573),
.A2(n_1411),
.B(n_1384),
.Y(n_1631)
);

AO31x2_ASAP7_75t_L g1632 ( 
.A1(n_1580),
.A2(n_1446),
.A3(n_1418),
.B(n_1362),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1620),
.A2(n_1598),
.B(n_1565),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1596),
.A2(n_1408),
.B(n_1369),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1513),
.Y(n_1635)
);

O2A1O1Ixp5_ASAP7_75t_L g1636 ( 
.A1(n_1517),
.A2(n_1529),
.B(n_1626),
.C(n_1571),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_SL g1637 ( 
.A1(n_1528),
.A2(n_1437),
.B(n_1442),
.C(n_1449),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_SL g1638 ( 
.A1(n_1545),
.A2(n_1424),
.B(n_1473),
.C(n_1435),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1516),
.B(n_1438),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1523),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1570),
.A2(n_1363),
.B(n_1420),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1574),
.A2(n_1453),
.B(n_1443),
.C(n_1422),
.Y(n_1642)
);

AOI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1593),
.A2(n_1415),
.B(n_1407),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1586),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1514),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1524),
.B(n_1438),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1526),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1607),
.A2(n_1399),
.B(n_1441),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1519),
.A2(n_1428),
.B(n_1451),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1605),
.A2(n_1438),
.B(n_1450),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1581),
.A2(n_1450),
.B1(n_1404),
.B2(n_36),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1551),
.A2(n_542),
.B(n_541),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1569),
.A2(n_547),
.B(n_544),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1579),
.A2(n_550),
.B(n_549),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1539),
.A2(n_554),
.B(n_551),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1624),
.A2(n_557),
.B(n_556),
.Y(n_1656)
);

AOI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1531),
.A2(n_34),
.B(n_35),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1590),
.A2(n_1618),
.B(n_1615),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1537),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1535),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1538),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1546),
.Y(n_1662)
);

O2A1O1Ixp5_ASAP7_75t_L g1663 ( 
.A1(n_1592),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_R g1664 ( 
.A1(n_1567),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1603),
.A2(n_559),
.A3(n_560),
.B(n_558),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1543),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1586),
.Y(n_1667)
);

AOI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1583),
.A2(n_562),
.B(n_561),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1556),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1542),
.B(n_40),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1536),
.B(n_563),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1588),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1672)
);

NAND3x1_ASAP7_75t_L g1673 ( 
.A(n_1625),
.B(n_41),
.C(n_42),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1601),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1553),
.B(n_43),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1541),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1616),
.A2(n_565),
.B(n_564),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1611),
.A2(n_1595),
.B1(n_1544),
.B2(n_1518),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_SL g1679 ( 
.A1(n_1594),
.A2(n_567),
.B(n_568),
.C(n_566),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1548),
.B(n_1610),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1563),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_SL g1682 ( 
.A1(n_1566),
.A2(n_570),
.B(n_571),
.C(n_569),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_R g1683 ( 
.A(n_1515),
.B(n_573),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1602),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1549),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1527),
.A2(n_1577),
.B1(n_1554),
.B2(n_1568),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1533),
.A2(n_575),
.B(n_574),
.Y(n_1687)
);

AOI31xp67_ASAP7_75t_L g1688 ( 
.A1(n_1630),
.A2(n_578),
.A3(n_582),
.B(n_577),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1564),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1575),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1520),
.A2(n_584),
.B(n_583),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1552),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1527),
.B(n_46),
.Y(n_1693)
);

AOI221x1_ASAP7_75t_L g1694 ( 
.A1(n_1582),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.C(n_50),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1525),
.A2(n_587),
.B(n_585),
.Y(n_1695)
);

AOI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1606),
.A2(n_589),
.B(n_588),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1530),
.A2(n_591),
.B(n_590),
.Y(n_1697)
);

AOI221x1_ASAP7_75t_L g1698 ( 
.A1(n_1600),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.C(n_52),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1512),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1560),
.A2(n_593),
.B(n_592),
.Y(n_1700)
);

AO21x1_ASAP7_75t_L g1701 ( 
.A1(n_1612),
.A2(n_56),
.B(n_55),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1532),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1584),
.B(n_54),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1558),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1550),
.A2(n_596),
.B(n_595),
.Y(n_1705)
);

AOI31xp67_ASAP7_75t_L g1706 ( 
.A1(n_1599),
.A2(n_598),
.A3(n_600),
.B(n_597),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1614),
.A2(n_1623),
.B(n_1557),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1597),
.Y(n_1708)
);

OAI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1572),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1534),
.B(n_60),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1627),
.A2(n_603),
.B(n_602),
.Y(n_1711)
);

O2A1O1Ixp33_ASAP7_75t_SL g1712 ( 
.A1(n_1608),
.A2(n_605),
.B(n_608),
.C(n_604),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1578),
.A2(n_611),
.B(n_609),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1515),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1629),
.A2(n_614),
.B(n_613),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1521),
.B(n_61),
.Y(n_1716)
);

AOI221x1_ASAP7_75t_L g1717 ( 
.A1(n_1585),
.A2(n_1562),
.B1(n_1547),
.B2(n_1587),
.C(n_1609),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1619),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1591),
.B(n_62),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1555),
.B(n_62),
.C(n_63),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1561),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_SL g1722 ( 
.A1(n_1604),
.A2(n_617),
.B(n_619),
.C(n_615),
.Y(n_1722)
);

AO31x2_ASAP7_75t_L g1723 ( 
.A1(n_1628),
.A2(n_622),
.A3(n_623),
.B(n_621),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1613),
.A2(n_625),
.B(n_624),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1591),
.B(n_629),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1621),
.A2(n_628),
.B(n_627),
.Y(n_1726)
);

AO31x2_ASAP7_75t_L g1727 ( 
.A1(n_1540),
.A2(n_1617),
.A3(n_1589),
.B(n_1522),
.Y(n_1727)
);

AOI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1576),
.A2(n_631),
.B(n_630),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_L g1729 ( 
.A(n_1576),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1617),
.B(n_63),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1617),
.A2(n_636),
.B(n_635),
.Y(n_1731)
);

BUFx2_ASAP7_75t_R g1732 ( 
.A(n_1559),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1622),
.B(n_64),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1596),
.A2(n_641),
.B(n_637),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1514),
.Y(n_1735)
);

OAI22x1_ASAP7_75t_L g1736 ( 
.A1(n_1574),
.A2(n_67),
.B1(n_68),
.B2(n_66),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1565),
.B(n_65),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1532),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1513),
.B(n_66),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1596),
.A2(n_644),
.B(n_643),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1573),
.A2(n_646),
.B(n_645),
.Y(n_1741)
);

AO21x1_ASAP7_75t_L g1742 ( 
.A1(n_1528),
.A2(n_70),
.B(n_69),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1565),
.B(n_68),
.Y(n_1743)
);

AO32x2_ASAP7_75t_L g1744 ( 
.A1(n_1626),
.A2(n_72),
.A3(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_1744)
);

AO32x2_ASAP7_75t_L g1745 ( 
.A1(n_1626),
.A2(n_74),
.A3(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_1745)
);

AO21x1_ASAP7_75t_L g1746 ( 
.A1(n_1528),
.A2(n_76),
.B(n_75),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1528),
.A2(n_649),
.B(n_647),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1596),
.A2(n_651),
.B(n_650),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1523),
.Y(n_1749)
);

AOI21x1_ASAP7_75t_SL g1750 ( 
.A1(n_1602),
.A2(n_74),
.B(n_76),
.Y(n_1750)
);

O2A1O1Ixp5_ASAP7_75t_L g1751 ( 
.A1(n_1517),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_1751)
);

OAI21x1_ASAP7_75t_L g1752 ( 
.A1(n_1596),
.A2(n_653),
.B(n_652),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1586),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1513),
.Y(n_1754)
);

AO32x2_ASAP7_75t_L g1755 ( 
.A1(n_1626),
.A2(n_79),
.A3(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1573),
.A2(n_655),
.B(n_654),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1536),
.B(n_656),
.Y(n_1757)
);

AOI221x1_ASAP7_75t_L g1758 ( 
.A1(n_1556),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.C(n_84),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1573),
.A2(n_659),
.B(n_657),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1573),
.A2(n_663),
.B(n_662),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1573),
.A2(n_665),
.B(n_664),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1523),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1553),
.B(n_81),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1528),
.A2(n_667),
.B(n_666),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1517),
.B(n_82),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1536),
.B(n_669),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1528),
.A2(n_671),
.B(n_670),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1523),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1765),
.A2(n_91),
.B1(n_99),
.B2(n_83),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1635),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1657),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1710),
.A2(n_95),
.B1(n_104),
.B2(n_86),
.Y(n_1772)
);

CKINVDCx11_ASAP7_75t_R g1773 ( 
.A(n_1738),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_87),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1754),
.Y(n_1775)
);

CKINVDCx6p67_ASAP7_75t_R g1776 ( 
.A(n_1667),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1702),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1644),
.B(n_672),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1645),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1763),
.B(n_87),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_88),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1640),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1736),
.A2(n_1664),
.B1(n_1719),
.B2(n_1716),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1659),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1681),
.Y(n_1785)
);

INVx5_ASAP7_75t_L g1786 ( 
.A(n_1635),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1691),
.A2(n_1764),
.B1(n_1747),
.B2(n_1720),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1729),
.A2(n_97),
.B1(n_108),
.B2(n_88),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1647),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1678),
.A2(n_92),
.B1(n_89),
.B2(n_90),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1735),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1680),
.Y(n_1793)
);

CKINVDCx6p67_ASAP7_75t_R g1794 ( 
.A(n_1753),
.Y(n_1794)
);

OAI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1674),
.A2(n_92),
.B1(n_89),
.B2(n_90),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1689),
.B(n_673),
.Y(n_1796)
);

CKINVDCx14_ASAP7_75t_R g1797 ( 
.A(n_1739),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1660),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1669),
.A2(n_1699),
.B1(n_1684),
.B2(n_1742),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1676),
.Y(n_1800)
);

AOI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1636),
.A2(n_93),
.B(n_94),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1766),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_SL g1803 ( 
.A1(n_1670),
.A2(n_103),
.B1(n_113),
.B2(n_93),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1714),
.B(n_674),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1666),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1718),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1762),
.B(n_1768),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1692),
.B(n_95),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1746),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1701),
.A2(n_101),
.B1(n_98),
.B2(n_100),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1708),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1703),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1721),
.B(n_675),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1690),
.Y(n_1814)
);

BUFx4f_ASAP7_75t_SL g1815 ( 
.A(n_1661),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1662),
.Y(n_1816)
);

BUFx12f_ASAP7_75t_L g1817 ( 
.A(n_1671),
.Y(n_1817)
);

INVx8_ASAP7_75t_L g1818 ( 
.A(n_1671),
.Y(n_1818)
);

BUFx12f_ASAP7_75t_L g1819 ( 
.A(n_1725),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1685),
.Y(n_1820)
);

BUFx8_ASAP7_75t_SL g1821 ( 
.A(n_1733),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1693),
.Y(n_1822)
);

CKINVDCx6p67_ASAP7_75t_R g1823 ( 
.A(n_1675),
.Y(n_1823)
);

CKINVDCx11_ASAP7_75t_R g1824 ( 
.A(n_1732),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1686),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1673),
.A2(n_107),
.B1(n_103),
.B2(n_105),
.Y(n_1826)
);

INVx6_ASAP7_75t_L g1827 ( 
.A(n_1683),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1709),
.A2(n_108),
.B1(n_105),
.B2(n_107),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1639),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1829)
);

INVx5_ASAP7_75t_L g1830 ( 
.A(n_1750),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1758),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1744),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1651),
.A2(n_115),
.B(n_114),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1727),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1646),
.A2(n_116),
.B1(n_112),
.B2(n_114),
.Y(n_1835)
);

INVx8_ASAP7_75t_L g1836 ( 
.A(n_1757),
.Y(n_1836)
);

INVx8_ASAP7_75t_L g1837 ( 
.A(n_1728),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1642),
.A2(n_117),
.B1(n_112),
.B2(n_116),
.Y(n_1838)
);

CKINVDCx11_ASAP7_75t_R g1839 ( 
.A(n_1704),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1744),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1658),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1713),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1745),
.Y(n_1843)
);

INVx6_ASAP7_75t_L g1844 ( 
.A(n_1730),
.Y(n_1844)
);

BUFx2_ASAP7_75t_SL g1845 ( 
.A(n_1731),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1650),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1641),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1696),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1672),
.A2(n_130),
.B1(n_138),
.B2(n_122),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1717),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1850)
);

INVx6_ASAP7_75t_L g1851 ( 
.A(n_1727),
.Y(n_1851)
);

CKINVDCx11_ASAP7_75t_R g1852 ( 
.A(n_1663),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1715),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1745),
.Y(n_1854)
);

AO22x1_ASAP7_75t_L g1855 ( 
.A1(n_1755),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1755),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1633),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1751),
.Y(n_1858)
);

INVx6_ASAP7_75t_L g1859 ( 
.A(n_1637),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1698),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1665),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1649),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1724),
.A2(n_138),
.B1(n_147),
.B2(n_129),
.Y(n_1863)
);

CKINVDCx20_ASAP7_75t_R g1864 ( 
.A(n_1677),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1665),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1694),
.B(n_131),
.Y(n_1866)
);

INVx6_ASAP7_75t_L g1867 ( 
.A(n_1767),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1726),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1638),
.Y(n_1869)
);

BUFx10_ASAP7_75t_L g1870 ( 
.A(n_1688),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1723),
.Y(n_1871)
);

NAND2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1705),
.B(n_676),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1707),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1652),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1697),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1643),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1723),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1653),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1741),
.A2(n_141),
.B1(n_137),
.B2(n_139),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1668),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1756),
.A2(n_1759),
.B1(n_1761),
.B2(n_1760),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1679),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1706),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1700),
.B(n_139),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1656),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1655),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1682),
.Y(n_1887)
);

BUFx2_ASAP7_75t_R g1888 ( 
.A(n_1712),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1632),
.B(n_144),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1695),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1734),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1711),
.Y(n_1892)
);

CKINVDCx12_ASAP7_75t_R g1893 ( 
.A(n_1722),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1687),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1654),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1740),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_1748),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1648),
.A2(n_1631),
.B(n_1752),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1632),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1634),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1782),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1791),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1783),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1789),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1792),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1784),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1786),
.B(n_677),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1811),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1798),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1814),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1805),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1816),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1807),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1786),
.Y(n_1914)
);

AO21x2_ASAP7_75t_L g1915 ( 
.A1(n_1880),
.A2(n_150),
.B(n_151),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1820),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1834),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1822),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1787),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1825),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1858),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1770),
.B(n_679),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1785),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1779),
.Y(n_1924)
);

INVxp33_ASAP7_75t_L g1925 ( 
.A(n_1800),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1883),
.A2(n_152),
.B(n_153),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1889),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1871),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1861),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1881),
.A2(n_681),
.B(n_680),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1773),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1775),
.B(n_154),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1851),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1876),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1859),
.Y(n_1935)
);

OR2x6_ASAP7_75t_L g1936 ( 
.A(n_1818),
.B(n_682),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1823),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1781),
.B(n_1774),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1891),
.A2(n_684),
.B(n_683),
.Y(n_1939)
);

OAI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1896),
.A2(n_686),
.B(n_685),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1808),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1851),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1790),
.B(n_155),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1832),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1840),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1806),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1813),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1884),
.A2(n_157),
.B(n_158),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1799),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1815),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1843),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1780),
.B(n_688),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1776),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1869),
.Y(n_1954)
);

INVx6_ASAP7_75t_L g1955 ( 
.A(n_1844),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1848),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1793),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1854),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1856),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1899),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1794),
.Y(n_1961)
);

AO21x2_ASAP7_75t_L g1962 ( 
.A1(n_1898),
.A2(n_160),
.B(n_161),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1833),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1797),
.B(n_689),
.Y(n_1964)
);

OR2x6_ASAP7_75t_L g1965 ( 
.A(n_1818),
.B(n_690),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1882),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1846),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1802),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1830),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1772),
.B(n_691),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1841),
.A2(n_694),
.B(n_692),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1887),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1836),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1802),
.B(n_696),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1836),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1777),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1827),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1830),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1877),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1866),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1850),
.B(n_163),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1865),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1895),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1902),
.B(n_1796),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1963),
.A2(n_1826),
.B1(n_1828),
.B2(n_1888),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1914),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1927),
.B(n_1852),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1967),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1948),
.A2(n_1874),
.B(n_1801),
.C(n_1847),
.Y(n_1989)
);

NAND2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1914),
.B(n_1853),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1930),
.A2(n_1868),
.B(n_1897),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1903),
.A2(n_1769),
.B1(n_1809),
.B2(n_1810),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1921),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1912),
.B(n_1875),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1904),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1905),
.B(n_1778),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1908),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1910),
.B(n_1778),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1913),
.B(n_1870),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1980),
.B(n_1863),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1918),
.B(n_1894),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1949),
.A2(n_1812),
.B1(n_1831),
.B2(n_1849),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1946),
.B(n_1864),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1916),
.B(n_1817),
.Y(n_2004)
);

INVx11_ASAP7_75t_L g2005 ( 
.A(n_1955),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1941),
.B(n_1855),
.Y(n_2006)
);

OR2x6_ASAP7_75t_L g2007 ( 
.A(n_1936),
.B(n_1837),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1925),
.B(n_1803),
.Y(n_2008)
);

NOR2x1_ASAP7_75t_SL g2009 ( 
.A(n_1962),
.B(n_1819),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1981),
.A2(n_1838),
.B(n_1892),
.C(n_1771),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1955),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1919),
.A2(n_1886),
.B(n_1885),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1983),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1938),
.B(n_1788),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1943),
.A2(n_1839),
.B1(n_1827),
.B2(n_1860),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1937),
.A2(n_1842),
.B(n_1857),
.C(n_1873),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1924),
.B(n_1835),
.Y(n_2017)
);

O2A1O1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1957),
.A2(n_1795),
.B(n_1879),
.C(n_1890),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1901),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1970),
.A2(n_1900),
.B1(n_1867),
.B2(n_1878),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1979),
.B(n_1862),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1906),
.B(n_1829),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1969),
.A2(n_1804),
.B(n_1872),
.Y(n_2023)
);

OAI21xp33_ASAP7_75t_L g2024 ( 
.A1(n_1932),
.A2(n_1893),
.B(n_1821),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1929),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1964),
.B(n_1845),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_SL g2027 ( 
.A(n_1953),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1920),
.B(n_1837),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1935),
.A2(n_1867),
.B1(n_1824),
.B2(n_166),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1952),
.B(n_164),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1911),
.B(n_165),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1909),
.B(n_167),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_1915),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.C(n_170),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_SL g2034 ( 
.A1(n_1936),
.A2(n_701),
.B(n_700),
.Y(n_2034)
);

NOR3xp33_ASAP7_75t_SL g2035 ( 
.A(n_1942),
.B(n_168),
.C(n_169),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_SL g2036 ( 
.A(n_1917),
.B(n_702),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1947),
.B(n_170),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1928),
.Y(n_2038)
);

A2O1A1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1978),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1966),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1933),
.B(n_703),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1931),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1944),
.B(n_172),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1933),
.B(n_704),
.Y(n_2044)
);

AO32x2_ASAP7_75t_L g2045 ( 
.A1(n_1945),
.A2(n_175),
.A3(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1968),
.B(n_705),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1951),
.B(n_174),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1965),
.A2(n_178),
.B1(n_175),
.B2(n_177),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1958),
.B(n_177),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1950),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1923),
.B(n_706),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1959),
.B(n_178),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1934),
.B(n_179),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1972),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_1940),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1956),
.B(n_180),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1960),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1976),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1988),
.B(n_1961),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1995),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_1994),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2015),
.A2(n_1965),
.B1(n_1977),
.B2(n_1973),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1993),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2001),
.B(n_1997),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2025),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2003),
.B(n_1987),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2038),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2004),
.B(n_1982),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1999),
.B(n_1954),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1996),
.B(n_1975),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2013),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2057),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2019),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2040),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_2024),
.B(n_1922),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2054),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2000),
.B(n_1926),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1998),
.B(n_2026),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1984),
.B(n_1922),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2028),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2008),
.B(n_1974),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2021),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2047),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1990),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2017),
.B(n_1974),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2053),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_2058),
.B(n_1907),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2056),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2007),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2032),
.Y(n_2090)
);

AOI22xp33_ASAP7_75t_L g2091 ( 
.A1(n_1985),
.A2(n_1926),
.B1(n_1939),
.B2(n_1971),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2006),
.B(n_181),
.Y(n_2092)
);

INVxp67_ASAP7_75t_L g2093 ( 
.A(n_1986),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2011),
.B(n_182),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2043),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_SL g2096 ( 
.A1(n_1992),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2049),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2014),
.B(n_183),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2050),
.B(n_184),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1986),
.Y(n_2100)
);

NOR2x1p5_ASAP7_75t_L g2101 ( 
.A(n_2042),
.B(n_185),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2052),
.B(n_185),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_2007),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2023),
.B(n_186),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2045),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_2022),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2037),
.B(n_186),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2045),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2031),
.B(n_187),
.Y(n_2109)
);

INVxp67_ASAP7_75t_SL g2110 ( 
.A(n_2009),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_2027),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2036),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_2005),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2036),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_2041),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_2051),
.B(n_187),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2030),
.B(n_188),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1991),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2010),
.B(n_189),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2044),
.B(n_2020),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_2046),
.B(n_190),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2029),
.B(n_190),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2055),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2018),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_2035),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2048),
.B(n_191),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2034),
.B(n_191),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1989),
.B(n_192),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2033),
.B(n_192),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2039),
.B(n_193),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2012),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_2002),
.B(n_193),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2016),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1988),
.B(n_194),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1993),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1988),
.B(n_194),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_1985),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1988),
.B(n_195),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1993),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2139),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_L g2141 ( 
.A(n_2132),
.B(n_198),
.C(n_196),
.D(n_197),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2106),
.B(n_198),
.Y(n_2142)
);

OAI31xp33_ASAP7_75t_L g2143 ( 
.A1(n_2133),
.A2(n_201),
.A3(n_199),
.B(n_200),
.Y(n_2143)
);

AO21x2_ASAP7_75t_L g2144 ( 
.A1(n_2110),
.A2(n_199),
.B(n_200),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2082),
.B(n_201),
.Y(n_2145)
);

AO21x2_ASAP7_75t_L g2146 ( 
.A1(n_2118),
.A2(n_202),
.B(n_203),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2078),
.B(n_202),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_2061),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2139),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2063),
.Y(n_2150)
);

NAND4xp25_ASAP7_75t_L g2151 ( 
.A(n_2128),
.B(n_206),
.C(n_204),
.D(n_205),
.Y(n_2151)
);

AOI211xp5_ASAP7_75t_L g2152 ( 
.A1(n_2119),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2111),
.B(n_207),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2061),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_2096),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_2111),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_SL g2157 ( 
.A1(n_2137),
.A2(n_210),
.B(n_211),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2060),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2065),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2089),
.B(n_210),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2070),
.B(n_211),
.Y(n_2161)
);

OAI21xp33_ASAP7_75t_L g2162 ( 
.A1(n_2123),
.A2(n_212),
.B(n_213),
.Y(n_2162)
);

OAI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_2131),
.A2(n_212),
.B(n_213),
.Y(n_2163)
);

AOI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2124),
.A2(n_2129),
.B1(n_2123),
.B2(n_2130),
.C(n_2125),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2067),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2103),
.Y(n_2166)
);

NAND3xp33_ASAP7_75t_L g2167 ( 
.A(n_2077),
.B(n_215),
.C(n_216),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2071),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_2104),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2169)
);

INVxp67_ASAP7_75t_L g2170 ( 
.A(n_2086),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_2103),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2135),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2080),
.B(n_2059),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2074),
.B(n_217),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2064),
.B(n_218),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2104),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_2084),
.B(n_219),
.Y(n_2177)
);

INVx4_ASAP7_75t_L g2178 ( 
.A(n_2121),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2072),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2076),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2073),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2066),
.B(n_220),
.Y(n_2182)
);

AO21x2_ASAP7_75t_L g2183 ( 
.A1(n_2105),
.A2(n_222),
.B(n_223),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2092),
.B(n_222),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2083),
.B(n_223),
.Y(n_2185)
);

OA21x2_ASAP7_75t_L g2186 ( 
.A1(n_2105),
.A2(n_224),
.B(n_225),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2095),
.B(n_224),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2068),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2069),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2097),
.B(n_225),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2108),
.Y(n_2191)
);

AOI221xp5_ASAP7_75t_L g2192 ( 
.A1(n_2108),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2088),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2090),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2112),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2085),
.B(n_227),
.Y(n_2196)
);

INVx2_ASAP7_75t_SL g2197 ( 
.A(n_2100),
.Y(n_2197)
);

CKINVDCx20_ASAP7_75t_R g2198 ( 
.A(n_2113),
.Y(n_2198)
);

OAI31xp33_ASAP7_75t_L g2199 ( 
.A1(n_2127),
.A2(n_230),
.A3(n_228),
.B(n_229),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_2121),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2062),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2201)
);

OAI21xp33_ASAP7_75t_L g2202 ( 
.A1(n_2126),
.A2(n_231),
.B(n_232),
.Y(n_2202)
);

OAI33xp33_ASAP7_75t_L g2203 ( 
.A1(n_2098),
.A2(n_2109),
.A3(n_2107),
.B1(n_2093),
.B2(n_2114),
.B3(n_236),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2134),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2115),
.B(n_233),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2079),
.B(n_233),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2081),
.B(n_235),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2136),
.Y(n_2208)
);

NAND4xp25_ASAP7_75t_L g2209 ( 
.A(n_2122),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_2209)
);

BUFx2_ASAP7_75t_L g2210 ( 
.A(n_2115),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2120),
.B(n_237),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_2091),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2138),
.Y(n_2213)
);

NAND4xp25_ASAP7_75t_SL g2214 ( 
.A(n_2099),
.B(n_242),
.C(n_240),
.D(n_241),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2075),
.A2(n_244),
.B1(n_241),
.B2(n_243),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2094),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2102),
.Y(n_2217)
);

BUFx2_ASAP7_75t_L g2218 ( 
.A(n_2101),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2087),
.B(n_243),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2117),
.B(n_244),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_2116),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2133),
.A2(n_248),
.B1(n_245),
.B2(n_247),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2082),
.Y(n_2223)
);

INVx5_ASAP7_75t_SL g2224 ( 
.A(n_2121),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2060),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2060),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2133),
.B(n_248),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2106),
.B(n_249),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2060),
.Y(n_2229)
);

INVxp67_ASAP7_75t_SL g2230 ( 
.A(n_2106),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2139),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2106),
.B(n_249),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2139),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2133),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2139),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2106),
.B(n_250),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2106),
.B(n_251),
.Y(n_2237)
);

NOR3xp33_ASAP7_75t_L g2238 ( 
.A(n_2128),
.B(n_252),
.C(n_254),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2148),
.B(n_254),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2189),
.B(n_255),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2166),
.B(n_255),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2171),
.B(n_256),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2195),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2223),
.B(n_256),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2140),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2210),
.B(n_2230),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2154),
.B(n_257),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_2186),
.Y(n_2248)
);

AND2x4_ASAP7_75t_SL g2249 ( 
.A(n_2198),
.B(n_257),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2173),
.B(n_258),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2188),
.B(n_258),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2156),
.B(n_259),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2149),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2231),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2170),
.B(n_260),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2194),
.B(n_261),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2233),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2235),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2193),
.B(n_262),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2150),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_2178),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_2191),
.B(n_262),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2204),
.B(n_2208),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2213),
.B(n_263),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2159),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2165),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2216),
.B(n_263),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2172),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2168),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_2218),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2180),
.B(n_264),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2158),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2217),
.B(n_264),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_2227),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_2225),
.B(n_265),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2179),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2197),
.B(n_2200),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_2218),
.Y(n_2278)
);

BUFx3_ASAP7_75t_L g2279 ( 
.A(n_2205),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2181),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2226),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_2177),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2229),
.B(n_265),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2174),
.B(n_266),
.Y(n_2284)
);

AND2x4_ASAP7_75t_SL g2285 ( 
.A(n_2160),
.B(n_267),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2186),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2175),
.B(n_268),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2187),
.Y(n_2288)
);

AOI21xp33_ASAP7_75t_L g2289 ( 
.A1(n_2152),
.A2(n_268),
.B(n_269),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2145),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2236),
.B(n_270),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2185),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_2238),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2142),
.B(n_271),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2228),
.B(n_2232),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2237),
.B(n_272),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2224),
.B(n_2147),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2146),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2183),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2190),
.Y(n_2300)
);

NAND2xp67_ASAP7_75t_L g2301 ( 
.A(n_2211),
.B(n_273),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2224),
.B(n_273),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_2206),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2161),
.B(n_274),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_2144),
.Y(n_2305)
);

OAI31xp33_ASAP7_75t_L g2306 ( 
.A1(n_2167),
.A2(n_276),
.A3(n_274),
.B(n_275),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2196),
.B(n_275),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2207),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2203),
.B(n_2184),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2182),
.B(n_276),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2164),
.B(n_277),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2153),
.B(n_277),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2220),
.Y(n_2313)
);

AND2x4_ASAP7_75t_SL g2314 ( 
.A(n_2219),
.B(n_278),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2209),
.B(n_278),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2212),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2199),
.B(n_279),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2221),
.Y(n_2318)
);

INVxp67_ASAP7_75t_L g2319 ( 
.A(n_2214),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2151),
.B(n_279),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2202),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2169),
.B(n_280),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2201),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2162),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2176),
.B(n_280),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2141),
.B(n_281),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2215),
.B(n_282),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2163),
.B(n_282),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2143),
.B(n_2234),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2192),
.B(n_283),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2222),
.B(n_284),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2155),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2157),
.B(n_284),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2203),
.B(n_286),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2230),
.B(n_287),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2140),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2230),
.B(n_287),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2189),
.B(n_288),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2148),
.B(n_289),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_2186),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2140),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2148),
.B(n_289),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2218),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2148),
.B(n_290),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2148),
.B(n_290),
.Y(n_2345)
);

AND2x4_ASAP7_75t_SL g2346 ( 
.A(n_2198),
.B(n_291),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2186),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2189),
.B(n_291),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2189),
.B(n_292),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2148),
.B(n_292),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2253),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_2278),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2249),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2282),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2270),
.B(n_293),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2343),
.B(n_293),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2254),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2309),
.B(n_294),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2298),
.Y(n_2359)
);

OA21x2_ASAP7_75t_L g2360 ( 
.A1(n_2248),
.A2(n_294),
.B(n_295),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2257),
.Y(n_2361)
);

INVxp67_ASAP7_75t_L g2362 ( 
.A(n_2305),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2289),
.A2(n_295),
.B(n_296),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_2274),
.B(n_296),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2246),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2336),
.Y(n_2366)
);

INVx2_ASAP7_75t_SL g2367 ( 
.A(n_2282),
.Y(n_2367)
);

O2A1O1Ixp33_ASAP7_75t_L g2368 ( 
.A1(n_2311),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2341),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2305),
.B(n_297),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2346),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2243),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2261),
.B(n_299),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_L g2374 ( 
.A(n_2329),
.B(n_301),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2269),
.Y(n_2375)
);

OR2x2_ASAP7_75t_L g2376 ( 
.A(n_2313),
.B(n_2290),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2280),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2277),
.B(n_302),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2288),
.B(n_302),
.Y(n_2379)
);

INVx2_ASAP7_75t_SL g2380 ( 
.A(n_2279),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2240),
.B(n_303),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2272),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2260),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_2271),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2245),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2265),
.Y(n_2386)
);

AND2x4_ASAP7_75t_SL g2387 ( 
.A(n_2318),
.B(n_303),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2303),
.B(n_304),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2266),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2292),
.B(n_304),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2268),
.Y(n_2391)
);

INVxp67_ASAP7_75t_SL g2392 ( 
.A(n_2248),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2276),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2258),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2281),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2338),
.B(n_305),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2348),
.B(n_306),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2340),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2263),
.B(n_306),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2349),
.B(n_307),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2340),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2347),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2347),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2295),
.B(n_307),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2271),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2308),
.B(n_308),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2286),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2299),
.B(n_308),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2300),
.B(n_309),
.Y(n_2409)
);

OR2x6_ASAP7_75t_L g2410 ( 
.A(n_2241),
.B(n_310),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2275),
.Y(n_2411)
);

AND2x4_ASAP7_75t_SL g2412 ( 
.A(n_2297),
.B(n_310),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2262),
.Y(n_2413)
);

INVxp67_ASAP7_75t_L g2414 ( 
.A(n_2334),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2264),
.B(n_311),
.Y(n_2415)
);

NOR2x1_ASAP7_75t_L g2416 ( 
.A(n_2335),
.B(n_2337),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2250),
.B(n_2239),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_SL g2418 ( 
.A1(n_2321),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_2418)
);

NOR2x1p5_ASAP7_75t_SL g2419 ( 
.A(n_2323),
.B(n_312),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2339),
.B(n_313),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2283),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2342),
.B(n_315),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2344),
.B(n_315),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2259),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2256),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2255),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2345),
.B(n_317),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2251),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2256),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2244),
.Y(n_2430)
);

OR2x2_ASAP7_75t_L g2431 ( 
.A(n_2316),
.B(n_317),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2267),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2273),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2247),
.Y(n_2434)
);

INVxp67_ASAP7_75t_L g2435 ( 
.A(n_2324),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2242),
.B(n_318),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2350),
.B(n_318),
.Y(n_2437)
);

OR2x6_ASAP7_75t_L g2438 ( 
.A(n_2302),
.B(n_319),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_2332),
.B(n_319),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2252),
.B(n_320),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2291),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_2284),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2287),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2294),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2301),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2319),
.B(n_320),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2312),
.B(n_321),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2315),
.B(n_321),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2326),
.Y(n_2449)
);

NOR2x1_ASAP7_75t_L g2450 ( 
.A(n_2296),
.B(n_322),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2304),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2307),
.B(n_323),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2310),
.B(n_323),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2328),
.B(n_324),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2317),
.Y(n_2455)
);

OR2x6_ASAP7_75t_L g2456 ( 
.A(n_2333),
.B(n_324),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2327),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2320),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2285),
.B(n_325),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2330),
.Y(n_2460)
);

INVx3_ASAP7_75t_L g2461 ( 
.A(n_2314),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2322),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2325),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2331),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2306),
.B(n_325),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2293),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2270),
.B(n_328),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2253),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2253),
.Y(n_2469)
);

AOI22x1_ASAP7_75t_L g2470 ( 
.A1(n_2305),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2253),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2270),
.B(n_329),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2253),
.Y(n_2473)
);

NAND2xp33_ASAP7_75t_L g2474 ( 
.A(n_2329),
.B(n_330),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2270),
.B(n_331),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2253),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2305),
.B(n_331),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2305),
.B(n_332),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2305),
.B(n_332),
.Y(n_2479)
);

NAND2x1_ASAP7_75t_L g2480 ( 
.A(n_2248),
.B(n_334),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2309),
.B(n_334),
.Y(n_2481)
);

OR2x2_ASAP7_75t_L g2482 ( 
.A(n_2270),
.B(n_335),
.Y(n_2482)
);

HB1xp67_ASAP7_75t_L g2483 ( 
.A(n_2298),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2270),
.B(n_335),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2270),
.B(n_336),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2329),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_2249),
.Y(n_2487)
);

OR2x2_ASAP7_75t_L g2488 ( 
.A(n_2270),
.B(n_337),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2305),
.B(n_340),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2270),
.B(n_340),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2253),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2305),
.B(n_341),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2270),
.B(n_341),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2309),
.B(n_342),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2282),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2270),
.B(n_342),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2253),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2309),
.A2(n_343),
.B(n_344),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2278),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2253),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2253),
.Y(n_2501)
);

AND2x4_ASAP7_75t_SL g2502 ( 
.A(n_2318),
.B(n_343),
.Y(n_2502)
);

INVx1_ASAP7_75t_SL g2503 ( 
.A(n_2249),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2270),
.B(n_344),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2289),
.A2(n_345),
.B(n_346),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2253),
.Y(n_2506)
);

INVxp67_ASAP7_75t_L g2507 ( 
.A(n_2305),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2298),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2253),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2253),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2305),
.B(n_345),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2270),
.B(n_346),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2309),
.B(n_347),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2305),
.B(n_348),
.Y(n_2514)
);

CKINVDCx16_ASAP7_75t_R g2515 ( 
.A(n_2279),
.Y(n_2515)
);

NAND2xp33_ASAP7_75t_SL g2516 ( 
.A(n_2305),
.B(n_348),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2278),
.B(n_349),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2455),
.B(n_349),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2449),
.B(n_350),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2515),
.B(n_350),
.Y(n_2520)
);

NAND4xp25_ASAP7_75t_L g2521 ( 
.A(n_2358),
.B(n_353),
.C(n_351),
.D(n_352),
.Y(n_2521)
);

OR2x2_ASAP7_75t_L g2522 ( 
.A(n_2376),
.B(n_352),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2407),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_2441),
.B(n_354),
.Y(n_2524)
);

AOI211xp5_ASAP7_75t_L g2525 ( 
.A1(n_2374),
.A2(n_357),
.B(n_354),
.C(n_355),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2384),
.B(n_357),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2365),
.B(n_358),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2444),
.B(n_358),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2460),
.B(n_359),
.Y(n_2529)
);

OR2x2_ASAP7_75t_L g2530 ( 
.A(n_2435),
.B(n_359),
.Y(n_2530)
);

INVx1_ASAP7_75t_SL g2531 ( 
.A(n_2353),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2398),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2352),
.B(n_360),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2380),
.B(n_360),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2405),
.B(n_361),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2499),
.B(n_361),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_2457),
.B(n_362),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2443),
.B(n_2411),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2414),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2425),
.B(n_365),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2351),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2357),
.Y(n_2542)
);

OR2x2_ASAP7_75t_L g2543 ( 
.A(n_2413),
.B(n_366),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2464),
.B(n_366),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2429),
.B(n_367),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2361),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2366),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2516),
.Y(n_2548)
);

NOR2x1_ASAP7_75t_L g2549 ( 
.A(n_2360),
.B(n_368),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2430),
.B(n_368),
.Y(n_2550)
);

BUFx2_ASAP7_75t_L g2551 ( 
.A(n_2442),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2426),
.B(n_369),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2392),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2354),
.B(n_370),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2367),
.B(n_370),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2495),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2424),
.B(n_2458),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2462),
.B(n_371),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2369),
.Y(n_2559)
);

NOR2xp67_ASAP7_75t_L g2560 ( 
.A(n_2362),
.B(n_372),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2434),
.B(n_372),
.Y(n_2561)
);

OR2x6_ASAP7_75t_L g2562 ( 
.A(n_2480),
.B(n_373),
.Y(n_2562)
);

OR2x2_ASAP7_75t_L g2563 ( 
.A(n_2372),
.B(n_373),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2421),
.B(n_374),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2468),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_SL g2566 ( 
.A(n_2371),
.B(n_375),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2463),
.B(n_2416),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2428),
.B(n_2370),
.Y(n_2568)
);

NOR2xp67_ASAP7_75t_L g2569 ( 
.A(n_2507),
.B(n_375),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2451),
.B(n_376),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2477),
.B(n_377),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2375),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2478),
.B(n_377),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2417),
.B(n_378),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2382),
.B(n_378),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2498),
.A2(n_379),
.B(n_380),
.Y(n_2576)
);

AND3x1_ASAP7_75t_L g2577 ( 
.A(n_2481),
.B(n_2513),
.C(n_2494),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2432),
.B(n_380),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2433),
.B(n_381),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2378),
.B(n_382),
.Y(n_2580)
);

NAND2xp33_ASAP7_75t_SL g2581 ( 
.A(n_2465),
.B(n_382),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2469),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2474),
.A2(n_383),
.B(n_384),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2399),
.B(n_385),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2404),
.B(n_385),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2401),
.B(n_386),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2402),
.Y(n_2587)
);

NAND3xp33_ASAP7_75t_L g2588 ( 
.A(n_2368),
.B(n_387),
.C(n_389),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2385),
.Y(n_2589)
);

INVxp67_ASAP7_75t_L g2590 ( 
.A(n_2360),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2355),
.B(n_387),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2471),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2403),
.B(n_389),
.Y(n_2593)
);

NOR2x1_ASAP7_75t_L g2594 ( 
.A(n_2479),
.B(n_390),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2473),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2476),
.Y(n_2596)
);

INVx2_ASAP7_75t_SL g2597 ( 
.A(n_2517),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2356),
.B(n_2467),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2395),
.B(n_2394),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2489),
.A2(n_390),
.B(n_392),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2491),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_SL g2602 ( 
.A(n_2492),
.B(n_393),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2359),
.Y(n_2603)
);

OR2x2_ASAP7_75t_L g2604 ( 
.A(n_2408),
.B(n_394),
.Y(n_2604)
);

OR2x2_ASAP7_75t_L g2605 ( 
.A(n_2431),
.B(n_394),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2497),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2472),
.B(n_395),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2475),
.B(n_396),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2511),
.B(n_396),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2484),
.B(n_397),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2500),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2514),
.B(n_397),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2461),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2501),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2490),
.B(n_398),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2466),
.B(n_398),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2506),
.Y(n_2617)
);

OR2x2_ASAP7_75t_L g2618 ( 
.A(n_2377),
.B(n_399),
.Y(n_2618)
);

OAI31xp33_ASAP7_75t_SL g2619 ( 
.A1(n_2450),
.A2(n_402),
.A3(n_400),
.B(n_401),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2517),
.Y(n_2620)
);

CKINVDCx16_ASAP7_75t_R g2621 ( 
.A(n_2438),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2445),
.B(n_401),
.Y(n_2622)
);

INVx1_ASAP7_75t_SL g2623 ( 
.A(n_2487),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2509),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2510),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2383),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2483),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2493),
.B(n_402),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2386),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2389),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2496),
.B(n_404),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2391),
.Y(n_2632)
);

OR2x2_ASAP7_75t_L g2633 ( 
.A(n_2393),
.B(n_404),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2448),
.B(n_405),
.Y(n_2634)
);

OR2x2_ASAP7_75t_L g2635 ( 
.A(n_2379),
.B(n_405),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2508),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2390),
.Y(n_2637)
);

INVx1_ASAP7_75t_SL g2638 ( 
.A(n_2503),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2504),
.B(n_406),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2409),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2512),
.B(n_406),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2551),
.B(n_2482),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2531),
.B(n_2439),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2553),
.Y(n_2644)
);

AOI221xp5_ASAP7_75t_L g2645 ( 
.A1(n_2577),
.A2(n_2446),
.B1(n_2486),
.B2(n_2363),
.C(n_2505),
.Y(n_2645)
);

OAI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2621),
.A2(n_2456),
.B1(n_2470),
.B2(n_2410),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2587),
.Y(n_2647)
);

OAI21xp33_ASAP7_75t_L g2648 ( 
.A1(n_2619),
.A2(n_2418),
.B(n_2419),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2523),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2538),
.Y(n_2650)
);

NAND2x1_ASAP7_75t_L g2651 ( 
.A(n_2549),
.B(n_2410),
.Y(n_2651)
);

NOR2x1_ASAP7_75t_L g2652 ( 
.A(n_2560),
.B(n_2438),
.Y(n_2652)
);

OAI221xp5_ASAP7_75t_L g2653 ( 
.A1(n_2576),
.A2(n_2456),
.B1(n_2364),
.B2(n_2454),
.C(n_2447),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2613),
.Y(n_2654)
);

AOI21xp33_ASAP7_75t_L g2655 ( 
.A1(n_2590),
.A2(n_2396),
.B(n_2381),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2581),
.A2(n_2397),
.B1(n_2400),
.B2(n_2412),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2629),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2623),
.B(n_2638),
.Y(n_2658)
);

O2A1O1Ixp33_ASAP7_75t_L g2659 ( 
.A1(n_2548),
.A2(n_2488),
.B(n_2485),
.C(n_2437),
.Y(n_2659)
);

OR2x2_ASAP7_75t_L g2660 ( 
.A(n_2637),
.B(n_2436),
.Y(n_2660)
);

AO221x1_ASAP7_75t_L g2661 ( 
.A1(n_2532),
.A2(n_2388),
.B1(n_2502),
.B2(n_2387),
.C(n_2373),
.Y(n_2661)
);

OAI221xp5_ASAP7_75t_L g2662 ( 
.A1(n_2588),
.A2(n_2525),
.B1(n_2583),
.B2(n_2602),
.C(n_2521),
.Y(n_2662)
);

INVx1_ASAP7_75t_SL g2663 ( 
.A(n_2520),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2556),
.B(n_2406),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2586),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2597),
.B(n_2420),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2598),
.B(n_2422),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_L g2668 ( 
.A1(n_2567),
.A2(n_2440),
.B1(n_2427),
.B2(n_2423),
.C(n_2459),
.Y(n_2668)
);

NAND3xp33_ASAP7_75t_SL g2669 ( 
.A(n_2600),
.B(n_2453),
.C(n_2452),
.Y(n_2669)
);

INVx2_ASAP7_75t_SL g2670 ( 
.A(n_2620),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2640),
.B(n_2415),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2539),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_2672)
);

OAI221xp5_ASAP7_75t_L g2673 ( 
.A1(n_2557),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.C(n_410),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2630),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2541),
.Y(n_2675)
);

OAI221xp5_ASAP7_75t_L g2676 ( 
.A1(n_2568),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.C(n_413),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2558),
.B(n_411),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2542),
.Y(n_2678)
);

NAND3xp33_ASAP7_75t_SL g2679 ( 
.A(n_2566),
.B(n_412),
.C(n_413),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2546),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2547),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2574),
.B(n_414),
.Y(n_2682)
);

AOI221xp5_ASAP7_75t_L g2683 ( 
.A1(n_2603),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_L g2684 ( 
.A(n_2519),
.B(n_415),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2569),
.B(n_418),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2518),
.B(n_2550),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2570),
.B(n_418),
.Y(n_2687)
);

NAND4xp75_ASAP7_75t_SL g2688 ( 
.A(n_2634),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_2688)
);

OAI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2562),
.A2(n_423),
.B1(n_419),
.B2(n_422),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2522),
.B(n_422),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2586),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2562),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2559),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2529),
.B(n_423),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2578),
.B(n_424),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2594),
.B(n_424),
.Y(n_2696)
);

OAI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2622),
.A2(n_425),
.B(n_426),
.Y(n_2697)
);

OAI22xp33_ASAP7_75t_L g2698 ( 
.A1(n_2627),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_2698)
);

OA222x2_ASAP7_75t_L g2699 ( 
.A1(n_2636),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.C1(n_430),
.C2(n_431),
.Y(n_2699)
);

OAI32xp33_ASAP7_75t_L g2700 ( 
.A1(n_2534),
.A2(n_433),
.A3(n_429),
.B1(n_430),
.B2(n_434),
.Y(n_2700)
);

AOI321xp33_ASAP7_75t_L g2701 ( 
.A1(n_2616),
.A2(n_433),
.A3(n_435),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_2701)
);

INVx2_ASAP7_75t_SL g2702 ( 
.A(n_2593),
.Y(n_2702)
);

AND2x2_ASAP7_75t_SL g2703 ( 
.A(n_2658),
.B(n_2526),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2644),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2647),
.Y(n_2705)
);

NAND4xp25_ASAP7_75t_SL g2706 ( 
.A(n_2645),
.B(n_2662),
.C(n_2652),
.D(n_2683),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2665),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2671),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2663),
.B(n_2593),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2692),
.B(n_2533),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2665),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2667),
.B(n_2702),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2691),
.B(n_2579),
.Y(n_2713)
);

NAND3xp33_ASAP7_75t_SL g2714 ( 
.A(n_2651),
.B(n_2604),
.C(n_2573),
.Y(n_2714)
);

AOI221xp5_ASAP7_75t_L g2715 ( 
.A1(n_2646),
.A2(n_2582),
.B1(n_2595),
.B2(n_2592),
.C(n_2565),
.Y(n_2715)
);

XNOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2688),
.B(n_2641),
.Y(n_2716)
);

A2O1A1Ixp33_ASAP7_75t_L g2717 ( 
.A1(n_2648),
.A2(n_2530),
.B(n_2605),
.C(n_2571),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2657),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2642),
.Y(n_2719)
);

O2A1O1Ixp33_ASAP7_75t_L g2720 ( 
.A1(n_2679),
.A2(n_2612),
.B(n_2609),
.C(n_2544),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2643),
.A2(n_2589),
.B1(n_2564),
.B2(n_2561),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2670),
.B(n_2536),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2664),
.B(n_2572),
.Y(n_2723)
);

OAI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2673),
.A2(n_2633),
.B1(n_2618),
.B2(n_2528),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2674),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2649),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_SL g2727 ( 
.A1(n_2661),
.A2(n_2607),
.B1(n_2608),
.B2(n_2591),
.Y(n_2727)
);

AOI322xp5_ASAP7_75t_L g2728 ( 
.A1(n_2669),
.A2(n_2639),
.A3(n_2631),
.B1(n_2628),
.B2(n_2610),
.C1(n_2615),
.C2(n_2584),
.Y(n_2728)
);

OAI322xp33_ASAP7_75t_L g2729 ( 
.A1(n_2676),
.A2(n_2611),
.A3(n_2632),
.B1(n_2626),
.B2(n_2625),
.C1(n_2624),
.C2(n_2617),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2668),
.B(n_2535),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2654),
.B(n_2563),
.Y(n_2731)
);

OAI211xp5_ASAP7_75t_L g2732 ( 
.A1(n_2701),
.A2(n_2596),
.B(n_2606),
.C(n_2601),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2659),
.A2(n_2552),
.B(n_2524),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2686),
.B(n_2575),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2650),
.Y(n_2735)
);

OAI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2697),
.A2(n_2599),
.B(n_2543),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2706),
.A2(n_2655),
.B(n_2696),
.Y(n_2737)
);

OAI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2727),
.A2(n_2672),
.B(n_2689),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2735),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2711),
.B(n_2666),
.Y(n_2740)
);

INVx2_ASAP7_75t_SL g2741 ( 
.A(n_2707),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2703),
.Y(n_2742)
);

OAI21xp33_ASAP7_75t_L g2743 ( 
.A1(n_2730),
.A2(n_2660),
.B(n_2675),
.Y(n_2743)
);

INVxp67_ASAP7_75t_L g2744 ( 
.A(n_2710),
.Y(n_2744)
);

OAI21x1_ASAP7_75t_L g2745 ( 
.A1(n_2735),
.A2(n_2680),
.B(n_2678),
.Y(n_2745)
);

AOI221x1_ASAP7_75t_L g2746 ( 
.A1(n_2733),
.A2(n_2685),
.B1(n_2684),
.B2(n_2694),
.C(n_2693),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2728),
.B(n_2656),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2723),
.Y(n_2748)
);

OR2x2_ASAP7_75t_L g2749 ( 
.A(n_2709),
.B(n_2690),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2708),
.Y(n_2750)
);

OR2x2_ASAP7_75t_L g2751 ( 
.A(n_2713),
.B(n_2681),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2714),
.A2(n_2724),
.B1(n_2732),
.B2(n_2715),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2704),
.Y(n_2753)
);

XNOR2x1_ASAP7_75t_L g2754 ( 
.A(n_2716),
.B(n_2635),
.Y(n_2754)
);

OAI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2719),
.A2(n_2653),
.B1(n_2698),
.B2(n_2537),
.Y(n_2755)
);

NAND2x1_ASAP7_75t_L g2756 ( 
.A(n_2739),
.B(n_2722),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2749),
.Y(n_2757)
);

NAND4xp25_ASAP7_75t_L g2758 ( 
.A(n_2752),
.B(n_2712),
.C(n_2717),
.D(n_2705),
.Y(n_2758)
);

NOR3x1_ASAP7_75t_L g2759 ( 
.A(n_2738),
.B(n_2734),
.C(n_2731),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2751),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2754),
.B(n_2744),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2742),
.B(n_2736),
.Y(n_2762)
);

NAND4xp25_ASAP7_75t_L g2763 ( 
.A(n_2737),
.B(n_2720),
.C(n_2725),
.D(n_2718),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2740),
.B(n_2721),
.Y(n_2764)
);

AOI321xp33_ASAP7_75t_L g2765 ( 
.A1(n_2761),
.A2(n_2747),
.A3(n_2743),
.B1(n_2755),
.B2(n_2748),
.C(n_2750),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2758),
.B(n_2741),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2763),
.A2(n_2753),
.B1(n_2726),
.B2(n_2614),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_R g2768 ( 
.A(n_2757),
.B(n_2760),
.Y(n_2768)
);

NAND3xp33_ASAP7_75t_L g2769 ( 
.A(n_2756),
.B(n_2746),
.C(n_2687),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2762),
.A2(n_2729),
.B1(n_2745),
.B2(n_2682),
.Y(n_2770)
);

AOI221xp5_ASAP7_75t_L g2771 ( 
.A1(n_2764),
.A2(n_2700),
.B1(n_2695),
.B2(n_2677),
.C(n_2699),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_SL g2772 ( 
.A(n_2759),
.B(n_2580),
.Y(n_2772)
);

AOI311xp33_ASAP7_75t_L g2773 ( 
.A1(n_2766),
.A2(n_2545),
.A3(n_2540),
.B(n_2555),
.C(n_2554),
.Y(n_2773)
);

INVx1_ASAP7_75t_SL g2774 ( 
.A(n_2772),
.Y(n_2774)
);

AOI221xp5_ASAP7_75t_L g2775 ( 
.A1(n_2770),
.A2(n_2585),
.B1(n_2527),
.B2(n_438),
.C(n_435),
.Y(n_2775)
);

AOI221xp5_ASAP7_75t_L g2776 ( 
.A1(n_2769),
.A2(n_440),
.B1(n_436),
.B2(n_439),
.C(n_441),
.Y(n_2776)
);

AOI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_2771),
.A2(n_2768),
.B1(n_2767),
.B2(n_2765),
.C(n_442),
.Y(n_2777)
);

AND3x2_ASAP7_75t_L g2778 ( 
.A(n_2776),
.B(n_439),
.C(n_441),
.Y(n_2778)
);

NOR3xp33_ASAP7_75t_L g2779 ( 
.A(n_2777),
.B(n_442),
.C(n_444),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2779),
.A2(n_2774),
.B1(n_2775),
.B2(n_2773),
.Y(n_2780)
);

AOI211xp5_ASAP7_75t_L g2781 ( 
.A1(n_2780),
.A2(n_2778),
.B(n_447),
.C(n_445),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2781),
.Y(n_2782)
);

NOR2x1_ASAP7_75t_L g2783 ( 
.A(n_2782),
.B(n_446),
.Y(n_2783)
);

XOR2x1_ASAP7_75t_L g2784 ( 
.A(n_2782),
.B(n_446),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2784),
.Y(n_2785)
);

CKINVDCx20_ASAP7_75t_R g2786 ( 
.A(n_2783),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2785),
.B(n_447),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2787),
.B(n_2786),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2788),
.B(n_448),
.Y(n_2789)
);

OAI21x1_ASAP7_75t_L g2790 ( 
.A1(n_2788),
.A2(n_448),
.B(n_449),
.Y(n_2790)
);

XNOR2xp5_ASAP7_75t_L g2791 ( 
.A(n_2789),
.B(n_449),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2790),
.Y(n_2792)
);

AOI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_2792),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.C(n_453),
.Y(n_2793)
);

AOI211xp5_ASAP7_75t_L g2794 ( 
.A1(n_2793),
.A2(n_2791),
.B(n_452),
.C(n_450),
.Y(n_2794)
);


endmodule