module real_aes_7124_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_575;
wire n_210;
wire n_325;
wire n_212;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g574 ( .A1(n_0), .A2(n_174), .B(n_575), .C(n_578), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_1), .B(n_520), .Y(n_579) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g127 ( .A(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g208 ( .A(n_3), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_4), .B(n_166), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_489), .B(n_514), .Y(n_513) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_6), .A2(n_151), .B(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_7), .A2(n_36), .B1(n_160), .B2(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_8), .B(n_151), .Y(n_177) );
AND2x6_ASAP7_75t_L g175 ( .A(n_9), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_10), .A2(n_175), .B(n_479), .C(n_481), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_11), .A2(n_460), .B1(n_752), .B2(n_753), .C1(n_762), .C2(n_766), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_12), .B(n_37), .Y(n_128) );
INVx1_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
INVx1_ASAP7_75t_L g201 ( .A(n_14), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_15), .B(n_164), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_16), .B(n_166), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_17), .B(n_152), .Y(n_213) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_18), .A2(n_151), .A3(n_181), .B1(n_192), .B2(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_19), .B(n_160), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_20), .B(n_152), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_21), .A2(n_56), .B1(n_160), .B2(n_238), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g260 ( .A1(n_22), .A2(n_84), .B1(n_160), .B2(n_164), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_23), .B(n_160), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_24), .A2(n_192), .B(n_479), .C(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_25), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_25), .Y(n_754) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_26), .A2(n_192), .B(n_479), .C(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_27), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_28), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_29), .A2(n_489), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_30), .B(n_194), .Y(n_232) );
INVx2_ASAP7_75t_L g162 ( .A(n_31), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_32), .A2(n_491), .B(n_499), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_33), .B(n_160), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_34), .B(n_194), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_35), .B(n_246), .Y(n_509) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_38), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_39), .B(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_40), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_41), .A2(n_80), .B1(n_758), .B2(n_759), .Y(n_757) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_41), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_42), .B(n_166), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_43), .B(n_489), .Y(n_506) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_44), .A2(n_81), .B1(n_141), .B2(n_142), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_44), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_45), .A2(n_491), .B(n_493), .C(n_499), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_46), .A2(n_757), .B1(n_760), .B2(n_761), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_46), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_47), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g576 ( .A(n_48), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_49), .A2(n_93), .B1(n_238), .B2(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g494 ( .A(n_50), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_51), .B(n_160), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_52), .B(n_160), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_53), .A2(n_131), .B1(n_132), .B2(n_135), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_53), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_54), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_55), .B(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_SL g217 ( .A1(n_57), .A2(n_61), .B1(n_160), .B2(n_164), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_58), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_59), .B(n_160), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_60), .B(n_160), .Y(n_243) );
INVx1_ASAP7_75t_L g176 ( .A(n_62), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_63), .B(n_489), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_64), .B(n_520), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_65), .A2(n_172), .B(n_204), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_66), .B(n_160), .Y(n_209) );
INVx1_ASAP7_75t_L g155 ( .A(n_67), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_68), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_69), .B(n_166), .Y(n_530) );
AO32x2_ASAP7_75t_L g256 ( .A1(n_70), .A2(n_151), .A3(n_192), .B1(n_257), .B2(n_261), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_71), .B(n_167), .Y(n_482) );
INVx1_ASAP7_75t_L g187 ( .A(n_72), .Y(n_187) );
INVx1_ASAP7_75t_L g227 ( .A(n_73), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g573 ( .A(n_74), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_75), .B(n_496), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_76), .A2(n_479), .B(n_499), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_77), .B(n_164), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_78), .Y(n_515) );
INVx1_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_80), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_81), .Y(n_142) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_81), .A2(n_142), .B1(n_143), .B2(n_453), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_82), .A2(n_89), .B1(n_133), .B2(n_134), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_82), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_83), .B(n_495), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_85), .B(n_238), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_86), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_87), .B(n_164), .Y(n_231) );
INVx2_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_89), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_90), .B(n_191), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_91), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
OR2x2_ASAP7_75t_L g124 ( .A(n_92), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_126), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_94), .A2(n_104), .B1(n_164), .B2(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_95), .B(n_489), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_96), .Y(n_529) );
INVxp67_ASAP7_75t_L g518 ( .A(n_97), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_98), .A2(n_106), .B1(n_117), .B2(n_771), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_99), .B(n_164), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g475 ( .A(n_101), .Y(n_475) );
INVx1_ASAP7_75t_L g553 ( .A(n_102), .Y(n_553) );
AND2x2_ASAP7_75t_L g501 ( .A(n_103), .B(n_194), .Y(n_501) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx12_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g772 ( .A(n_109), .Y(n_772) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
OR2x2_ASAP7_75t_L g751 ( .A(n_113), .B(n_126), .Y(n_751) );
NOR2x2_ASAP7_75t_L g768 ( .A(n_113), .B(n_125), .Y(n_768) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_458), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g770 ( .A(n_120), .Y(n_770) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B(n_454), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g457 ( .A(n_124), .Y(n_457) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
XOR2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_136), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_134), .B(n_218), .Y(n_557) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B1(n_143), .B2(n_453), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g453 ( .A(n_143), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_377), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_335), .Y(n_144) );
NOR4xp25_ASAP7_75t_L g145 ( .A(n_146), .B(n_275), .C(n_311), .D(n_325), .Y(n_145) );
OAI221xp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_219), .B1(n_251), .B2(n_262), .C(n_266), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_147), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_195), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_178), .Y(n_149) );
AND2x2_ASAP7_75t_L g272 ( .A(n_150), .B(n_179), .Y(n_272) );
INVx3_ASAP7_75t_L g280 ( .A(n_150), .Y(n_280) );
AND2x2_ASAP7_75t_L g334 ( .A(n_150), .B(n_198), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_150), .B(n_197), .Y(n_370) );
AND2x2_ASAP7_75t_L g428 ( .A(n_150), .B(n_290), .Y(n_428) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_157), .B(n_177), .Y(n_150) );
INVx4_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_151), .A2(n_506), .B(n_507), .Y(n_505) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_151), .Y(n_512) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_153), .B(n_154), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_169), .B(n_175), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_166), .Y(n_158) );
INVx3_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_160), .Y(n_555) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g238 ( .A(n_161), .Y(n_238) );
BUFx3_ASAP7_75t_L g259 ( .A(n_161), .Y(n_259) );
AND2x6_ASAP7_75t_L g479 ( .A(n_161), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
INVx1_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
INVx2_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_166), .A2(n_184), .B(n_185), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_SL g225 ( .A1(n_166), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_166), .B(n_518), .Y(n_517) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g257 ( .A1(n_167), .A2(n_191), .B1(n_258), .B2(n_260), .Y(n_257) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_168), .Y(n_191) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_168), .Y(n_206) );
INVx1_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
AND2x2_ASAP7_75t_L g477 ( .A(n_168), .B(n_173), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_168), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_174), .Y(n_169) );
INVx2_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_174), .A2(n_188), .B(n_208), .C(n_209), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_174), .A2(n_191), .B1(n_216), .B2(n_217), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_174), .A2(n_191), .B1(n_237), .B2(n_239), .Y(n_236) );
BUFx3_ASAP7_75t_L g192 ( .A(n_175), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_175), .A2(n_200), .B(n_207), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_175), .A2(n_225), .B(n_229), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_175), .A2(n_242), .B(n_247), .Y(n_241) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_175), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g489 ( .A(n_175), .B(n_477), .Y(n_489) );
INVx4_ASAP7_75t_SL g500 ( .A(n_175), .Y(n_500) );
AND2x2_ASAP7_75t_L g263 ( .A(n_178), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_178), .B(n_198), .Y(n_277) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_179), .B(n_198), .Y(n_292) );
AND2x2_ASAP7_75t_L g304 ( .A(n_179), .B(n_280), .Y(n_304) );
OR2x2_ASAP7_75t_L g306 ( .A(n_179), .B(n_264), .Y(n_306) );
AND2x2_ASAP7_75t_L g341 ( .A(n_179), .B(n_264), .Y(n_341) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_179), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_179), .Y(n_394) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_182), .B(n_193), .Y(n_179) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_180), .A2(n_199), .B(n_210), .Y(n_198) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_181), .B(n_485), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_192), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .C(n_190), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_188), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_190), .A2(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx4_ASAP7_75t_L g577 ( .A(n_191), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g214 ( .A(n_192), .B(n_215), .C(n_218), .Y(n_214) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_194), .A2(n_224), .B(n_232), .Y(n_223) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_194), .A2(n_241), .B(n_250), .Y(n_240) );
INVx2_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_194), .A2(n_488), .B(n_490), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_194), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g546 ( .A(n_194), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_195), .A2(n_312), .B1(n_316), .B2(n_320), .C(n_321), .Y(n_311) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g271 ( .A(n_196), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
INVx2_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
AND2x2_ASAP7_75t_L g323 ( .A(n_197), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g342 ( .A(n_197), .B(n_280), .Y(n_342) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g405 ( .A(n_198), .B(n_280), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .C(n_204), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_202), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_202), .A2(n_509), .B(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_204), .A2(n_553), .B(n_554), .C(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_230), .B(n_231), .Y(n_229) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g496 ( .A(n_206), .Y(n_496) );
AND2x2_ASAP7_75t_L g327 ( .A(n_211), .B(n_272), .Y(n_327) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_211), .A2(n_351), .A3(n_396), .B1(n_398), .B2(n_401), .C1(n_403), .C2(n_407), .Y(n_395) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_212), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g291 ( .A(n_212), .Y(n_291) );
AND2x2_ASAP7_75t_L g400 ( .A(n_212), .B(n_280), .Y(n_400) );
AND2x2_ASAP7_75t_L g432 ( .A(n_212), .B(n_304), .Y(n_432) );
OR2x2_ASAP7_75t_L g435 ( .A(n_212), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
AO21x1_ASAP7_75t_L g264 ( .A1(n_215), .A2(n_218), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_218), .A2(n_474), .B(n_484), .Y(n_473) );
INVx3_ASAP7_75t_L g520 ( .A(n_218), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_218), .B(n_532), .Y(n_531) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_218), .A2(n_550), .B(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_233), .Y(n_220) );
INVx1_ASAP7_75t_L g448 ( .A(n_221), .Y(n_448) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g253 ( .A(n_222), .B(n_240), .Y(n_253) );
INVx2_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g310 ( .A(n_223), .Y(n_310) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
OR2x2_ASAP7_75t_L g442 ( .A(n_223), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g267 ( .A(n_233), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g307 ( .A(n_233), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g359 ( .A(n_233), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
AND2x2_ASAP7_75t_L g254 ( .A(n_234), .B(n_255), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g314 ( .A(n_234), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_256), .Y(n_368) );
OR2x2_ASAP7_75t_L g376 ( .A(n_234), .B(n_310), .Y(n_376) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
BUFx2_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_235), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g319 ( .A(n_235), .B(n_240), .Y(n_319) );
AND2x2_ASAP7_75t_L g383 ( .A(n_235), .B(n_256), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_240), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_240), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g296 ( .A(n_240), .Y(n_296) );
INVx1_ASAP7_75t_L g301 ( .A(n_240), .Y(n_301) );
AND2x2_ASAP7_75t_L g313 ( .A(n_240), .B(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_240), .Y(n_391) );
INVx1_ASAP7_75t_L g443 ( .A(n_240), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_245), .Y(n_242) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_329), .Y(n_420) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g347 ( .A(n_254), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g446 ( .A(n_254), .B(n_381), .Y(n_446) );
INVx1_ASAP7_75t_L g268 ( .A(n_255), .Y(n_268) );
AND2x2_ASAP7_75t_L g294 ( .A(n_255), .B(n_288), .Y(n_294) );
BUFx2_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
INVx1_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_259), .Y(n_498) );
INVx2_ASAP7_75t_L g578 ( .A(n_259), .Y(n_578) );
INVx1_ASAP7_75t_L g543 ( .A(n_261), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g422 ( .A(n_262), .B(n_269), .Y(n_422) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI32xp33_ASAP7_75t_L g266 ( .A1(n_263), .A2(n_267), .A3(n_269), .B1(n_271), .B2(n_273), .Y(n_266) );
AND2x2_ASAP7_75t_L g406 ( .A(n_263), .B(n_279), .Y(n_406) );
AND2x2_ASAP7_75t_L g444 ( .A(n_263), .B(n_342), .Y(n_444) );
INVx1_ASAP7_75t_L g324 ( .A(n_264), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_268), .B(n_330), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_269), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_269), .B(n_272), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_269), .B(n_341), .Y(n_423) );
OR2x2_ASAP7_75t_L g437 ( .A(n_269), .B(n_306), .Y(n_437) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g364 ( .A(n_270), .B(n_272), .Y(n_364) );
OR2x2_ASAP7_75t_L g373 ( .A(n_270), .B(n_360), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_272), .B(n_323), .Y(n_345) );
INVx2_ASAP7_75t_L g360 ( .A(n_274), .Y(n_360) );
OR2x2_ASAP7_75t_L g375 ( .A(n_274), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g390 ( .A(n_274), .B(n_391), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_274), .A2(n_367), .B(n_448), .C(n_449), .Y(n_447) );
OAI321xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_281), .A3(n_286), .B1(n_289), .B2(n_293), .C(n_297), .Y(n_275) );
INVx1_ASAP7_75t_L g388 ( .A(n_276), .Y(n_388) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g399 ( .A(n_277), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g351 ( .A(n_279), .Y(n_351) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_280), .B(n_394), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_281), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_424), .Y(n_418) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g356 ( .A(n_283), .B(n_330), .Y(n_356) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_284), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g371 ( .A1(n_286), .A2(n_327), .B(n_372), .C(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g338 ( .A(n_288), .B(n_295), .Y(n_338) );
BUFx2_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g363 ( .A(n_288), .Y(n_363) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
OR2x2_ASAP7_75t_L g369 ( .A(n_291), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g452 ( .A(n_291), .Y(n_452) );
INVx1_ASAP7_75t_L g445 ( .A(n_292), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g298 ( .A(n_294), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g402 ( .A(n_294), .B(n_319), .Y(n_402) );
INVx1_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B1(n_305), .B2(n_307), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_299), .B(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g367 ( .A(n_300), .B(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_301), .B(n_310), .Y(n_330) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g322 ( .A(n_304), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g332 ( .A(n_306), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_309), .A2(n_427), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g315 ( .A(n_310), .Y(n_315) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_310), .Y(n_381) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_313), .B(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_314), .A2(n_319), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_317), .B(n_327), .Y(n_424) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g393 ( .A(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g352 ( .A(n_319), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g441 ( .A(n_319), .Y(n_441) );
INVx1_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
INVx1_ASAP7_75t_L g412 ( .A(n_323), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_331), .B2(n_332), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_329), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g397 ( .A(n_330), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_330), .B(n_368), .Y(n_434) );
OR2x2_ASAP7_75t_L g407 ( .A(n_331), .B(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_334), .B(n_385), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_354), .C(n_365), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_343), .C(n_349), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_338), .A2(n_409), .B1(n_413), .B2(n_416), .C(n_418), .Y(n_408) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g350 ( .A(n_341), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g404 ( .A(n_341), .B(n_405), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_342), .A2(n_390), .B(n_392), .C(n_394), .Y(n_389) );
INVx2_ASAP7_75t_L g436 ( .A(n_342), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_346), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g415 ( .A(n_348), .B(n_368), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
OAI21xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_357), .B(n_358), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_364), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_359), .B(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_364), .B(n_451), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B(n_371), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g392 ( .A(n_368), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND4x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_408), .C(n_425), .D(n_447), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_395), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_384), .B(n_387), .C(n_389), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_383), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_394), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
INVx2_ASAP7_75t_SL g417 ( .A(n_405), .Y(n_417) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g425 ( .A(n_426), .B(n_433), .Y(n_425) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
OAI221xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_454), .B(n_459), .C(n_769), .Y(n_458) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_462), .B1(n_465), .B2(n_749), .Y(n_460) );
INVx1_ASAP7_75t_L g763 ( .A(n_461), .Y(n_763) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g764 ( .A(n_463), .Y(n_764) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_466), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
OR3x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_647), .C(n_712), .Y(n_466) );
NAND4xp25_ASAP7_75t_SL g467 ( .A(n_468), .B(n_588), .C(n_614), .D(n_637), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_521), .B1(n_558), .B2(n_565), .C(n_580), .Y(n_468) );
CKINVDCx14_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_470), .A2(n_581), .B1(n_605), .B2(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_502), .Y(n_470) );
INVx1_ASAP7_75t_SL g641 ( .A(n_471), .Y(n_641) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_486), .Y(n_471) );
OR2x2_ASAP7_75t_L g563 ( .A(n_472), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g583 ( .A(n_472), .B(n_503), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_472), .B(n_511), .Y(n_596) );
AND2x2_ASAP7_75t_L g613 ( .A(n_472), .B(n_486), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_472), .B(n_561), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_472), .B(n_612), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_472), .B(n_502), .Y(n_734) );
AOI211xp5_ASAP7_75t_SL g745 ( .A1(n_472), .A2(n_651), .B(n_746), .C(n_747), .Y(n_745) );
INVx5_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_473), .B(n_503), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_473), .B(n_504), .Y(n_620) );
OR2x2_ASAP7_75t_L g665 ( .A(n_473), .B(n_503), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_473), .B(n_511), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .Y(n_474) );
INVx5_ASAP7_75t_L g492 ( .A(n_479), .Y(n_492) );
INVx5_ASAP7_75t_SL g564 ( .A(n_486), .Y(n_564) );
AND2x2_ASAP7_75t_L g582 ( .A(n_486), .B(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_486), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_486), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g700 ( .A(n_486), .B(n_511), .Y(n_700) );
OR2x2_ASAP7_75t_L g706 ( .A(n_486), .B(n_596), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_486), .B(n_656), .Y(n_715) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_501), .Y(n_486) );
BUFx2_ASAP7_75t_L g538 ( .A(n_489), .Y(n_538) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_492), .A2(n_500), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g572 ( .A1(n_492), .A2(n_500), .B(n_573), .C(n_574), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_497), .C(n_498), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_495), .A2(n_498), .B(n_529), .C(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
AND2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_564), .Y(n_597) );
INVx1_ASAP7_75t_SL g610 ( .A(n_503), .Y(n_610) );
OR2x2_ASAP7_75t_L g645 ( .A(n_503), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g651 ( .A(n_503), .B(n_511), .Y(n_651) );
AND2x2_ASAP7_75t_L g709 ( .A(n_503), .B(n_561), .Y(n_709) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_504), .B(n_564), .Y(n_636) );
INVx3_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
OR2x2_ASAP7_75t_L g602 ( .A(n_511), .B(n_564), .Y(n_602) );
AND2x2_ASAP7_75t_L g612 ( .A(n_511), .B(n_610), .Y(n_612) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_511), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_511), .B(n_583), .Y(n_669) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_520), .A2(n_571), .B(n_579), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_521), .A2(n_686), .B1(n_688), .B2(n_690), .C(n_693), .Y(n_685) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
AND2x2_ASAP7_75t_L g659 ( .A(n_523), .B(n_640), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_523), .B(n_718), .Y(n_722) );
OR2x2_ASAP7_75t_L g743 ( .A(n_523), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_523), .B(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx5_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g667 ( .A(n_524), .B(n_535), .Y(n_667) );
AND2x2_ASAP7_75t_L g728 ( .A(n_524), .B(n_607), .Y(n_728) );
AND2x2_ASAP7_75t_L g741 ( .A(n_524), .B(n_561), .Y(n_741) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_547), .Y(n_533) );
AND2x4_ASAP7_75t_L g568 ( .A(n_534), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_534), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g593 ( .A(n_534), .Y(n_593) );
AND2x2_ASAP7_75t_L g662 ( .A(n_534), .B(n_640), .Y(n_662) );
AND2x2_ASAP7_75t_L g672 ( .A(n_534), .B(n_590), .Y(n_672) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_534), .Y(n_680) );
AND2x2_ASAP7_75t_L g692 ( .A(n_534), .B(n_570), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_534), .B(n_624), .Y(n_696) );
AND2x2_ASAP7_75t_L g733 ( .A(n_534), .B(n_728), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_534), .B(n_607), .Y(n_744) );
OR2x2_ASAP7_75t_L g746 ( .A(n_534), .B(n_682), .Y(n_746) );
INVx5_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g632 ( .A(n_535), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g642 ( .A(n_535), .B(n_587), .Y(n_642) );
AND2x2_ASAP7_75t_L g654 ( .A(n_535), .B(n_570), .Y(n_654) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_535), .Y(n_684) );
AND2x4_ASAP7_75t_L g718 ( .A(n_535), .B(n_569), .Y(n_718) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_544), .Y(n_535) );
AOI21xp5_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_539), .B(n_543), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
BUFx2_ASAP7_75t_L g567 ( .A(n_547), .Y(n_567) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g607 ( .A(n_548), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_548), .B(n_570), .Y(n_640) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g587 ( .A(n_549), .B(n_570), .Y(n_587) );
BUFx2_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_556), .Y(n_550) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_560), .B(n_641), .Y(n_720) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_561), .B(n_583), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_561), .B(n_564), .Y(n_622) );
AND2x2_ASAP7_75t_L g677 ( .A(n_561), .B(n_613), .Y(n_677) );
AOI221xp5_ASAP7_75t_SL g614 ( .A1(n_562), .A2(n_615), .B1(n_623), .B2(n_625), .C(n_629), .Y(n_614) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g609 ( .A(n_563), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g650 ( .A(n_563), .B(n_651), .Y(n_650) );
OAI321xp33_ASAP7_75t_L g657 ( .A1(n_563), .A2(n_616), .A3(n_658), .B1(n_660), .B2(n_661), .C(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_564), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_567), .B(n_718), .Y(n_736) );
AND2x2_ASAP7_75t_L g623 ( .A(n_568), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_568), .B(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_569), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_569), .B(n_681), .Y(n_711) );
INVx1_ASAP7_75t_L g748 ( .A(n_569), .Y(n_748) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B(n_585), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g740 ( .A1(n_582), .A2(n_692), .B(n_741), .C(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_583), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_583), .B(n_621), .Y(n_687) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g630 ( .A(n_587), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_587), .B(n_590), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_587), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_587), .B(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_603), .B2(n_608), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g604 ( .A(n_590), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g627 ( .A(n_590), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g639 ( .A(n_590), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_590), .B(n_633), .Y(n_675) );
OR2x2_ASAP7_75t_L g682 ( .A(n_590), .B(n_607), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_590), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g732 ( .A(n_590), .B(n_718), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B1(n_598), .B2(n_600), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g638 ( .A(n_593), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_596), .A2(n_611), .B1(n_679), .B2(n_683), .Y(n_678) );
INVx1_ASAP7_75t_L g726 ( .A(n_597), .Y(n_726) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_601), .A2(n_638), .B1(n_641), .B2(n_642), .C(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g616 ( .A(n_602), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_606), .B(n_672), .Y(n_704) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_607), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_607), .Y(n_628) );
NAND2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g646 ( .A(n_613), .Y(n_646) );
AND2x2_ASAP7_75t_L g655 ( .A(n_613), .B(n_656), .Y(n_655) );
NAND2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g699 ( .A(n_620), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_623), .A2(n_649), .B1(n_652), .B2(n_655), .C(n_657), .Y(n_648) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_627), .B(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_631), .B(n_634), .Y(n_629) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_634), .Y(n_731) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x2_ASAP7_75t_L g673 ( .A(n_636), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g694 ( .A(n_639), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_639), .B(n_699), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_642), .B(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_666), .C(n_685), .D(n_698), .Y(n_647) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g656 ( .A(n_651), .Y(n_656) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g689 ( .A(n_660), .B(n_665), .Y(n_689) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B(n_670), .C(n_678), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g737 ( .A1(n_668), .A2(n_710), .B(n_738), .C(n_745), .Y(n_737) );
INVx1_ASAP7_75t_SL g697 ( .A(n_669), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B1(n_675), .B2(n_676), .Y(n_670) );
INVx1_ASAP7_75t_L g701 ( .A(n_675), .Y(n_701) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_681), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_681), .B(n_692), .Y(n_725) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g702 ( .A(n_692), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_697), .Y(n_693) );
INVxp33_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .A3(n_702), .B1(n_703), .B2(n_705), .C1(n_707), .C2(n_710), .Y(n_698) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_730), .C(n_737), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B1(n_719), .B2(n_721), .C(n_723), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g729 ( .A(n_718), .Y(n_729) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_730) );
NAND2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g765 ( .A(n_750), .Y(n_765) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx16_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_757), .Y(n_760) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
endmodule