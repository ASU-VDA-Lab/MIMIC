module fake_jpeg_10888_n_648 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_648);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_73),
.Y(n_137)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_14),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_109),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_22),
.B(n_14),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_85),
.Y(n_146)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_14),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_107),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_13),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_46),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_97),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_96),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_21),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_22),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_58),
.Y(n_166)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_117),
.Y(n_127)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_0),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_120),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_25),
.B(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_49),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_130),
.B(n_164),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_31),
.B1(n_52),
.B2(n_35),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_132),
.A2(n_44),
.B(n_43),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_54),
.B1(n_46),
.B2(n_27),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_134),
.A2(n_142),
.B1(n_158),
.B2(n_173),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_84),
.A2(n_54),
.B1(n_30),
.B2(n_52),
.Y(n_142)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_153),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_72),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_157),
.B(n_170),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_75),
.A2(n_54),
.B1(n_30),
.B2(n_52),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_66),
.B(n_59),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_162),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_58),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_166),
.B(n_177),
.Y(n_252)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_95),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_175),
.B(n_181),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_100),
.B(n_58),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_179),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_72),
.A2(n_27),
.B(n_35),
.C(n_31),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_80),
.B(n_54),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_89),
.B(n_25),
.Y(n_181)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_25),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_79),
.A2(n_48),
.B1(n_41),
.B2(n_34),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_196),
.B1(n_39),
.B2(n_53),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_111),
.B(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_201),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_87),
.A2(n_48),
.B1(n_41),
.B2(n_34),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_98),
.A2(n_41),
.B1(n_34),
.B2(n_28),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_198),
.B1(n_43),
.B2(n_38),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_101),
.A2(n_28),
.B1(n_44),
.B2(n_29),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_113),
.B(n_29),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_60),
.B(n_44),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_179),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_146),
.A2(n_86),
.B1(n_76),
.B2(n_90),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_204),
.A2(n_216),
.B1(n_219),
.B2(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_149),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_207),
.B(n_225),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_83),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_213),
.C(n_215),
.Y(n_278)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_209),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_210),
.B(n_212),
.Y(n_324)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_94),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_127),
.B(n_91),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_214),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_123),
.B(n_104),
.C(n_116),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_134),
.A2(n_71),
.B1(n_67),
.B2(n_61),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_140),
.A2(n_196),
.B1(n_189),
.B2(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_220),
.B(n_229),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_269),
.B(n_210),
.Y(n_279)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_223),
.Y(n_326)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_224),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_176),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_226),
.Y(n_317)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_227),
.Y(n_333)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_125),
.B(n_63),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_133),
.C(n_136),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_38),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_232),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_233),
.B(n_241),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_234),
.B(n_235),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_137),
.B(n_102),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_158),
.A2(n_103),
.B1(n_115),
.B2(n_108),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_246),
.Y(n_288)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_130),
.B(n_155),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_249),
.Y(n_315)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_240),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_143),
.B(n_102),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_147),
.A2(n_118),
.B1(n_24),
.B2(n_37),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_129),
.B(n_24),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_145),
.B(n_24),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_265),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_105),
.B1(n_131),
.B2(n_182),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_253),
.A2(n_257),
.B(n_183),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_142),
.A2(n_106),
.B1(n_99),
.B2(n_68),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_254),
.A2(n_259),
.B1(n_260),
.B2(n_264),
.Y(n_292)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_191),
.A2(n_131),
.B1(n_151),
.B2(n_182),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_193),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_258),
.B(n_262),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_124),
.A2(n_39),
.B1(n_53),
.B2(n_50),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_124),
.A2(n_39),
.B1(n_53),
.B2(n_50),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_195),
.A2(n_96),
.B1(n_50),
.B2(n_43),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_151),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_23),
.B1(n_168),
.B2(n_169),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_147),
.A2(n_38),
.B1(n_37),
.B2(n_23),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_171),
.B1(n_205),
.B2(n_264),
.Y(n_301)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_156),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_273),
.Y(n_339)
);

CKINVDCx6p67_ASAP7_75t_R g270 ( 
.A(n_153),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_270),
.Y(n_287)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_161),
.Y(n_271)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_165),
.B(n_37),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_0),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_165),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_276),
.B(n_9),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_167),
.A2(n_23),
.B1(n_20),
.B2(n_96),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_236),
.B1(n_269),
.B2(n_216),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_279),
.A2(n_310),
.B1(n_336),
.B2(n_337),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_282),
.A2(n_298),
.B1(n_299),
.B2(n_304),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_148),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_300),
.C(n_307),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_229),
.A2(n_133),
.B(n_200),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_296),
.B(n_303),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_252),
.A2(n_169),
.B1(n_168),
.B2(n_126),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_206),
.A2(n_192),
.B1(n_172),
.B2(n_183),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_220),
.B(n_242),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_301),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_206),
.A2(n_266),
.B1(n_251),
.B2(n_219),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_311),
.B1(n_331),
.B2(n_335),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_208),
.B(n_161),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_185),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_312),
.C(n_313),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_218),
.A2(n_192),
.B1(n_159),
.B2(n_171),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_215),
.A2(n_186),
.B1(n_161),
.B2(n_178),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_242),
.A2(n_178),
.B(n_138),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_212),
.A2(n_40),
.B(n_20),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_212),
.A2(n_40),
.B(n_20),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_319),
.C(n_327),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_249),
.A2(n_40),
.B(n_20),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_239),
.B(n_186),
.C(n_40),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_335),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_250),
.A2(n_186),
.B1(n_21),
.B2(n_2),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_230),
.B(n_272),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_203),
.C(n_237),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_275),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_204),
.A2(n_228),
.B1(n_214),
.B2(n_232),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_228),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_340),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_324),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_343),
.B(n_367),
.Y(n_397)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_344),
.Y(n_396)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_347),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_281),
.B(n_207),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_351),
.B(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_221),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_294),
.B(n_255),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_357),
.B(n_360),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_291),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_286),
.B(n_231),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g363 ( 
.A(n_300),
.B(n_227),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_262),
.B1(n_226),
.B2(n_265),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_374),
.B1(n_377),
.B2(n_292),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_288),
.B(n_256),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_339),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_368),
.Y(n_437)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_370),
.B(n_372),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_278),
.B(n_211),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_378),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_286),
.B(n_247),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_243),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_373),
.B(n_375),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_226),
.B1(n_248),
.B2(n_217),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_231),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_376),
.B(n_381),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_290),
.A2(n_324),
.B1(n_298),
.B2(n_282),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_278),
.B(n_268),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_283),
.B(n_274),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_380),
.B(n_382),
.Y(n_428)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_284),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_284),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_383),
.B(n_384),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_261),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_291),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_390),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_303),
.A2(n_223),
.B1(n_263),
.B2(n_238),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_287),
.B1(n_326),
.B2(n_331),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_328),
.B(n_203),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_307),
.Y(n_402)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_280),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_293),
.Y(n_426)
);

AOI32xp33_ASAP7_75t_L g393 ( 
.A1(n_313),
.A2(n_244),
.A3(n_270),
.B1(n_273),
.B2(n_209),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_393),
.A2(n_289),
.B(n_279),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_394),
.A2(n_398),
.B(n_401),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_285),
.B(n_324),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g399 ( 
.A1(n_385),
.A2(n_358),
.A3(n_386),
.B1(n_343),
.B2(n_371),
.C1(n_378),
.C2(n_389),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_399),
.B(n_422),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_285),
.B(n_314),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_350),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_319),
.B(n_311),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_409),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_408),
.A2(n_414),
.B1(n_416),
.B2(n_423),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_388),
.A2(n_323),
.B(n_312),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_349),
.A2(n_336),
.B1(n_292),
.B2(n_310),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_377),
.A2(n_337),
.B1(n_296),
.B2(n_299),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_418),
.A2(n_431),
.B1(n_381),
.B2(n_375),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_350),
.B(n_308),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_380),
.C(n_391),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_386),
.A2(n_327),
.B(n_315),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_349),
.A2(n_315),
.B1(n_287),
.B2(n_326),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_366),
.A2(n_306),
.B(n_325),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_424),
.B(n_409),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_352),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_346),
.A2(n_326),
.B1(n_332),
.B2(n_306),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_427),
.A2(n_438),
.B1(n_355),
.B2(n_344),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_244),
.B(n_332),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_363),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_358),
.A2(n_330),
.B1(n_309),
.B2(n_302),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_348),
.A2(n_309),
.B1(n_322),
.B2(n_341),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_435),
.A2(n_418),
.B1(n_431),
.B2(n_382),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_346),
.A2(n_374),
.B1(n_365),
.B2(n_384),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_441),
.A2(n_473),
.B(n_400),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_423),
.B1(n_427),
.B2(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_452),
.C(n_454),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_360),
.C(n_354),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_447),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_426),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_432),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_448),
.B(n_449),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_433),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_413),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_451),
.B(n_457),
.Y(n_501)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_363),
.C(n_383),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_463),
.B1(n_467),
.B2(n_470),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_406),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_462),
.B1(n_471),
.B2(n_474),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_461),
.Y(n_496)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_408),
.A2(n_414),
.B1(n_416),
.B2(n_438),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_361),
.C(n_345),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_465),
.C(n_466),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_356),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_402),
.B(n_370),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_437),
.B(n_362),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_468),
.B(n_395),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_426),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_469),
.Y(n_512)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_364),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_410),
.B(n_392),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_476),
.C(n_419),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_413),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_417),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_412),
.A2(n_342),
.B1(n_369),
.B2(n_359),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_477),
.B1(n_469),
.B2(n_447),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_387),
.C(n_342),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_445),
.B(n_422),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_480),
.B(n_500),
.Y(n_532)
);

A2O1A1Ixp33_ASAP7_75t_SL g484 ( 
.A1(n_478),
.A2(n_398),
.B(n_401),
.C(n_394),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_SL g531 ( 
.A(n_484),
.B(n_489),
.C(n_470),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_462),
.A2(n_399),
.B1(n_406),
.B2(n_397),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_485),
.A2(n_491),
.B1(n_497),
.B2(n_320),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_486),
.A2(n_495),
.B1(n_503),
.B2(n_459),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_488),
.B(n_495),
.Y(n_519)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_454),
.B(n_409),
.CI(n_403),
.CON(n_489),
.SN(n_489)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_458),
.A2(n_397),
.B1(n_405),
.B2(n_430),
.Y(n_491)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_434),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_424),
.C(n_428),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_506),
.C(n_508),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_455),
.A2(n_405),
.B1(n_428),
.B2(n_412),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_458),
.A2(n_430),
.B1(n_419),
.B2(n_415),
.Y(n_497)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_498),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_435),
.B(n_415),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_499),
.A2(n_467),
.B(n_461),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_436),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_436),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_502),
.B(n_504),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_473),
.A2(n_400),
.B1(n_420),
.B2(n_425),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_425),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_443),
.B(n_395),
.C(n_435),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_450),
.B(n_411),
.Y(n_508)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_460),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_443),
.B(n_429),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_514),
.C(n_440),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_443),
.B(n_322),
.C(n_341),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_471),
.Y(n_515)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_516),
.A2(n_482),
.B1(n_518),
.B2(n_515),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_472),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_519),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_476),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_520),
.B(n_525),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_521),
.A2(n_507),
.B1(n_505),
.B2(n_494),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_463),
.Y(n_522)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_481),
.A2(n_477),
.B1(n_474),
.B2(n_444),
.Y(n_523)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_523),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_506),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_533),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_439),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_489),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_529),
.A2(n_530),
.B(n_491),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_513),
.B(n_453),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_531),
.B(n_537),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_499),
.A2(n_429),
.B(n_434),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_347),
.C(n_434),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_535),
.C(n_514),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_434),
.C(n_379),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_536),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_497),
.A2(n_271),
.B1(n_273),
.B2(n_240),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_538),
.A2(n_542),
.B1(n_487),
.B2(n_486),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_293),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_543),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_501),
.B(n_329),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_540),
.B(n_511),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_280),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_544),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_546),
.B(n_562),
.C(n_563),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_547),
.A2(n_564),
.B1(n_295),
.B2(n_270),
.Y(n_589)
);

FAx1_ASAP7_75t_SL g548 ( 
.A(n_519),
.B(n_489),
.CI(n_531),
.CON(n_548),
.SN(n_548)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_522),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_551),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_550),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_480),
.C(n_493),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_SL g553 ( 
.A(n_527),
.B(n_484),
.C(n_508),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_553),
.B(n_557),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_492),
.C(n_488),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_520),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_569),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_504),
.C(n_502),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_532),
.C(n_524),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_526),
.B(n_485),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_565),
.B(n_273),
.Y(n_587)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_566),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_532),
.B(n_528),
.C(n_541),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_541),
.C(n_484),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_525),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_571),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_576),
.B(n_585),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_530),
.C(n_533),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_578),
.C(n_579),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_530),
.C(n_529),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_557),
.B(n_542),
.C(n_484),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_581),
.A2(n_587),
.B(n_590),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_555),
.A2(n_543),
.B1(n_539),
.B2(n_224),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_582),
.A2(n_567),
.B1(n_553),
.B2(n_548),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_295),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_583),
.B(n_554),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_558),
.B(n_329),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_591),
.Y(n_599)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_320),
.C(n_270),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_558),
.C(n_556),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_589),
.B(n_550),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_569),
.A2(n_561),
.B(n_559),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_562),
.B(n_570),
.Y(n_591)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_592),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_572),
.B(n_568),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_594),
.B(n_600),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_596),
.B(n_601),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_576),
.B(n_556),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_597),
.B(n_598),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_559),
.C(n_552),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_580),
.A2(n_574),
.B1(n_582),
.B2(n_579),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_602),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_575),
.B(n_571),
.C(n_578),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_603),
.A2(n_605),
.B(n_606),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_577),
.A2(n_548),
.B1(n_1),
.B2(n_3),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_588),
.A2(n_0),
.B(n_3),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_3),
.C(n_4),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_607),
.A2(n_608),
.B(n_7),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_573),
.B(n_4),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_573),
.C(n_584),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_SL g625 ( 
.A(n_610),
.B(n_612),
.Y(n_625)
);

AOI21x1_ASAP7_75t_SL g611 ( 
.A1(n_604),
.A2(n_586),
.B(n_5),
.Y(n_611)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_611),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_600),
.B(n_4),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_595),
.B(n_4),
.C(n_6),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_615),
.B(n_616),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_6),
.C(n_7),
.Y(n_616)
);

BUFx24_ASAP7_75t_SL g618 ( 
.A(n_609),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_599),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_593),
.B(n_6),
.Y(n_622)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_622),
.Y(n_628)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_623),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_602),
.A2(n_7),
.B(n_8),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_605),
.B1(n_598),
.B2(n_596),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_607),
.Y(n_626)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_626),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_630),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_633),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_617),
.B(n_597),
.C(n_599),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_632),
.B(n_610),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_619),
.A2(n_7),
.B1(n_8),
.B2(n_613),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_635),
.B(n_639),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_620),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_617),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_632),
.B(n_615),
.Y(n_643)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_636),
.A2(n_625),
.B(n_621),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_641),
.A2(n_643),
.B1(n_637),
.B2(n_638),
.Y(n_644)
);

AOI221xp5_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_645),
.B1(n_627),
.B2(n_628),
.C(n_611),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_642),
.B(n_638),
.C(n_633),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_645),
.B1(n_616),
.B2(n_629),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_8),
.Y(n_648)
);


endmodule