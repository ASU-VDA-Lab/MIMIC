module real_jpeg_27948_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_0),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_65),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_48),
.B1(n_61),
.B2(n_62),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_40),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_54),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_11),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_79),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_79),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_56),
.B(n_60),
.C(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_12),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_58),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_12),
.B(n_38),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_38),
.B(n_42),
.C(n_182),
.D(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_12),
.B(n_70),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_12),
.A2(n_25),
.B(n_195),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g225 ( 
.A1(n_12),
.A2(n_62),
.B(n_73),
.C(n_111),
.D(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_12),
.B(n_62),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_13),
.A2(n_38),
.B(n_43),
.C(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_26),
.Y(n_183)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_21),
.B(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_22),
.B(n_80),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_52),
.C(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_36),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_25),
.A2(n_34),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_25),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_84),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_33),
.B1(n_104),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_25),
.B(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_30),
.A2(n_83),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_32),
.A2(n_39),
.A3(n_45),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_32),
.B(n_215),
.Y(n_214)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_37),
.A2(n_49),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_38),
.A2(n_61),
.A3(n_226),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_39),
.B(n_235),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_41),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_42),
.A2(n_46),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_42),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_42),
.A2(n_46),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_49),
.B(n_148),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_49),
.A2(n_146),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_49),
.B(n_99),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_57),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_58),
.B(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_62),
.B(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_62),
.B1(n_71),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_64),
.Y(n_128)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_72),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_69),
.B1(n_107),
.B2(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_78),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_69),
.A2(n_72),
.B(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_70),
.A2(n_73),
.B1(n_109),
.B2(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_71),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_86),
.Y(n_123)
);

INVx5_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_83),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_83),
.A2(n_211),
.B(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_88),
.A2(n_89),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.C(n_105),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_91),
.B1(n_105),
.B2(n_106),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_97),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_99),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_102),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_133),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_121),
.A2(n_202),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_132),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_174),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_158),
.B(n_173),
.Y(n_137)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.C(n_152),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_159),
.B(n_161),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_162),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_165),
.B(n_167),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_168),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_170),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_255),
.C(n_256),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_250),
.B(n_254),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_238),
.B(n_249),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_221),
.B(n_237),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_198),
.B(n_220),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_184),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_185),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_194),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_206),
.B(n_219),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_218),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_223),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.C(n_230),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.Y(n_245)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_245),
.C(n_246),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);


endmodule