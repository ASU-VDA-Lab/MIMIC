module real_aes_5356_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_174;
wire n_904;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_954;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g204 ( .A(n_0), .B(n_184), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_1), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_2), .A2(n_127), .B(n_257), .C(n_258), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_3), .A2(n_80), .B1(n_125), .B2(n_156), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_4), .A2(n_30), .B1(n_557), .B2(n_558), .Y(n_556) );
INVxp67_ASAP7_75t_L g514 ( .A(n_5), .Y(n_514) );
INVx1_ASAP7_75t_L g929 ( .A(n_5), .Y(n_929) );
INVx1_ASAP7_75t_L g934 ( .A(n_5), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_6), .A2(n_87), .B1(n_609), .B2(n_610), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_7), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g153 ( .A1(n_8), .A2(n_66), .B1(n_154), .B2(n_156), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_9), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_10), .A2(n_31), .B1(n_579), .B2(n_580), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_11), .Y(n_949) );
INVx2_ASAP7_75t_L g703 ( .A(n_12), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_13), .A2(n_58), .B1(n_125), .B2(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_14), .A2(n_65), .B(n_142), .Y(n_141) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_14), .A2(n_65), .B(n_142), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_15), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g701 ( .A(n_16), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_17), .B(n_160), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_18), .Y(n_230) );
BUFx3_ASAP7_75t_L g537 ( .A(n_19), .Y(n_537) );
BUFx8_ASAP7_75t_SL g958 ( .A(n_19), .Y(n_958) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_20), .A2(n_210), .B(n_263), .C(n_264), .Y(n_262) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_21), .A2(n_46), .B1(n_125), .B2(n_174), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_22), .A2(n_29), .B1(n_174), .B2(n_179), .Y(n_194) );
O2A1O1Ixp5_ASAP7_75t_L g652 ( .A1(n_23), .A2(n_560), .B(n_653), .C(n_656), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_24), .B(n_564), .Y(n_642) );
XOR2xp5_ASAP7_75t_L g935 ( .A(n_25), .B(n_936), .Y(n_935) );
O2A1O1Ixp5_ASAP7_75t_L g120 ( .A1(n_26), .A2(n_121), .B(n_124), .C(n_127), .Y(n_120) );
INVx1_ASAP7_75t_L g519 ( .A(n_27), .Y(n_519) );
INVx1_ASAP7_75t_SL g661 ( .A(n_28), .Y(n_661) );
AND2x2_ASAP7_75t_L g533 ( .A(n_32), .B(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_33), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_34), .B(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_35), .A2(n_39), .B1(n_563), .B2(n_565), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_36), .A2(n_64), .B1(n_565), .B2(n_597), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_37), .B(n_559), .Y(n_641) );
INVx2_ASAP7_75t_L g522 ( .A(n_38), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_40), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_41), .B(n_247), .Y(n_615) );
OAI22xp33_ASAP7_75t_SL g109 ( .A1(n_42), .A2(n_92), .B1(n_110), .B2(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_42), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_43), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_44), .A2(n_210), .B(n_699), .C(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g682 ( .A(n_45), .Y(n_682) );
INVx2_ASAP7_75t_L g662 ( .A(n_47), .Y(n_662) );
INVx1_ASAP7_75t_L g142 ( .A(n_48), .Y(n_142) );
AND2x4_ASAP7_75t_L g137 ( .A(n_49), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g159 ( .A(n_49), .B(n_138), .Y(n_159) );
INVx2_ASAP7_75t_L g598 ( .A(n_50), .Y(n_598) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_51), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_52), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_53), .Y(n_134) );
INVx2_ASAP7_75t_L g180 ( .A(n_54), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_55), .A2(n_127), .B(n_233), .C(n_234), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_56), .Y(n_217) );
INVx1_ASAP7_75t_SL g657 ( .A(n_57), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_59), .A2(n_75), .B1(n_196), .B2(n_197), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_60), .B(n_160), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_61), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_62), .Y(n_221) );
NAND2xp33_ASAP7_75t_R g161 ( .A(n_63), .B(n_146), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_63), .A2(n_102), .B1(n_200), .B2(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_67), .B(n_527), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_68), .A2(n_210), .B(n_557), .C(n_600), .Y(n_599) );
OR2x6_ASAP7_75t_L g516 ( .A(n_69), .B(n_517), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_70), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g668 ( .A(n_71), .Y(n_668) );
INVx1_ASAP7_75t_L g678 ( .A(n_72), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_73), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_74), .B(n_579), .Y(n_646) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_76), .B(n_121), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_77), .A2(n_127), .B(n_594), .C(n_596), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_77), .A2(n_127), .B(n_594), .C(n_596), .Y(n_627) );
INVx1_ASAP7_75t_L g518 ( .A(n_78), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_79), .A2(n_91), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_79), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_81), .A2(n_94), .B1(n_583), .B2(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g534 ( .A(n_82), .Y(n_534) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
BUFx5_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
INVx1_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
INVx2_ASAP7_75t_L g268 ( .A(n_84), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_85), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g237 ( .A(n_86), .Y(n_237) );
AOI22xp5_ASAP7_75t_SL g936 ( .A1(n_88), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_88), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_89), .Y(n_265) );
INVx2_ASAP7_75t_SL g138 ( .A(n_90), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_91), .Y(n_941) );
INVx1_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_95), .B(n_146), .Y(n_679) );
INVx1_ASAP7_75t_SL g572 ( .A(n_96), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_97), .B(n_602), .Y(n_664) );
INVx2_ASAP7_75t_L g144 ( .A(n_98), .Y(n_144) );
AND2x2_ASAP7_75t_L g587 ( .A(n_99), .B(n_171), .Y(n_587) );
OAI21xp33_ASAP7_75t_SL g228 ( .A1(n_100), .A2(n_125), .B(n_229), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_101), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_101), .Y(n_523) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_102), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_102), .B(n_200), .Y(n_291) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_529), .B(n_538), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_526), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B1(n_508), .B2(n_525), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OA22x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_109), .B1(n_112), .B2(n_507), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g507 ( .A(n_112), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g112 ( .A(n_113), .B(n_365), .C(n_436), .D(n_474), .Y(n_112) );
AND4x2_ASAP7_75t_L g930 ( .A(n_113), .B(n_365), .C(n_436), .D(n_474), .Y(n_930) );
NOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_303), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_115), .B(n_283), .Y(n_114) );
O2A1O1Ixp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_162), .B(n_186), .C(n_238), .Y(n_115) );
AND2x2_ASAP7_75t_L g297 ( .A(n_116), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_116), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g351 ( .A(n_116), .Y(n_351) );
AND2x2_ASAP7_75t_L g435 ( .A(n_116), .B(n_415), .Y(n_435) );
AND2x2_ASAP7_75t_L g442 ( .A(n_116), .B(n_240), .Y(n_442) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_147), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_117), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g499 ( .A(n_117), .B(n_399), .Y(n_499) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g270 ( .A(n_118), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g277 ( .A(n_118), .Y(n_277) );
BUFx2_ASAP7_75t_R g337 ( .A(n_118), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_118), .B(n_254), .Y(n_407) );
AND2x2_ASAP7_75t_L g411 ( .A(n_118), .B(n_253), .Y(n_411) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_139), .B(n_143), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_129), .C(n_136), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g130 ( .A(n_122), .Y(n_130) );
INVx1_ASAP7_75t_L g233 ( .A(n_122), .Y(n_233) );
INVx2_ASAP7_75t_L g559 ( .A(n_122), .Y(n_559) );
INVx2_ASAP7_75t_L g610 ( .A(n_122), .Y(n_610) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
INVx2_ASAP7_75t_L g156 ( .A(n_123), .Y(n_156) );
INVx6_ASAP7_75t_L g174 ( .A(n_123), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_125), .B(n_134), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_125), .A2(n_174), .B1(n_175), .B2(n_176), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g216 ( .A1(n_125), .A2(n_174), .B1(n_217), .B2(n_218), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_125), .A2(n_152), .B1(n_220), .B2(n_221), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_125), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g564 ( .A(n_125), .Y(n_564) );
INVx2_ASAP7_75t_L g579 ( .A(n_125), .Y(n_579) );
INVx2_ASAP7_75t_L g585 ( .A(n_125), .Y(n_585) );
INVx1_ASAP7_75t_L g595 ( .A(n_125), .Y(n_595) );
INVx2_ASAP7_75t_L g609 ( .A(n_125), .Y(n_609) );
NAND2xp33_ASAP7_75t_L g694 ( .A(n_125), .B(n_695), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_127), .A2(n_135), .B1(n_151), .B2(n_153), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g172 ( .A1(n_127), .A2(n_135), .B1(n_173), .B2(n_177), .Y(n_172) );
OAI221xp5_ASAP7_75t_L g215 ( .A1(n_127), .A2(n_159), .B1(n_210), .B2(n_216), .C(n_219), .Y(n_215) );
INVx1_ASAP7_75t_L g296 ( .A(n_127), .Y(n_296) );
INVx2_ASAP7_75t_SL g614 ( .A(n_127), .Y(n_614) );
INVx1_ASAP7_75t_L g647 ( .A(n_127), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_127), .B(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_127), .B(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_128), .B(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_128), .Y(n_193) );
INVx1_ASAP7_75t_L g198 ( .A(n_128), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_128), .B(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g210 ( .A(n_128), .Y(n_210) );
INVxp67_ASAP7_75t_L g612 ( .A(n_128), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B1(n_133), .B2(n_135), .Y(n_129) );
INVx2_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_SL g667 ( .A1(n_135), .A2(n_668), .B(n_669), .C(n_672), .Y(n_667) );
NOR2xp33_ASAP7_75t_SL g266 ( .A(n_136), .B(n_184), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_136), .A2(n_231), .B1(n_294), .B2(n_295), .C(n_296), .Y(n_293) );
NOR4xp25_ASAP7_75t_L g592 ( .A(n_136), .B(n_593), .C(n_599), .D(n_602), .Y(n_592) );
NOR2x1_ASAP7_75t_SL g691 ( .A(n_136), .B(n_214), .Y(n_691) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_137), .B(n_170), .Y(n_191) );
AND2x2_ASAP7_75t_L g225 ( .A(n_137), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_139), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g638 ( .A(n_139), .Y(n_638) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_140), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_140), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
BUFx3_ASAP7_75t_L g247 ( .A(n_141), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx1_ASAP7_75t_L g226 ( .A(n_146), .Y(n_226) );
INVx2_ASAP7_75t_L g384 ( .A(n_146), .Y(n_384) );
INVx1_ASAP7_75t_L g591 ( .A(n_146), .Y(n_591) );
INVx1_ASAP7_75t_SL g164 ( .A(n_147), .Y(n_164) );
INVx1_ASAP7_75t_L g278 ( .A(n_147), .Y(n_278) );
AND2x2_ASAP7_75t_L g360 ( .A(n_147), .B(n_253), .Y(n_360) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g271 ( .A(n_148), .Y(n_271) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_148), .Y(n_287) );
AND2x2_ASAP7_75t_L g408 ( .A(n_148), .B(n_167), .Y(n_408) );
AND2x2_ASAP7_75t_L g446 ( .A(n_148), .B(n_277), .Y(n_446) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_161), .Y(n_148) );
AND2x2_ASAP7_75t_L g381 ( .A(n_149), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_157), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g263 ( .A(n_152), .Y(n_263) );
INVx2_ASAP7_75t_L g580 ( .A(n_152), .Y(n_580) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_152), .Y(n_699) );
INVx2_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx2_ASAP7_75t_L g597 ( .A(n_156), .Y(n_597) );
INVx1_ASAP7_75t_L g673 ( .A(n_156), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_158), .B(n_247), .Y(n_663) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_159), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_185), .Y(n_211) );
INVx3_ASAP7_75t_L g570 ( .A(n_159), .Y(n_570) );
AND2x2_ASAP7_75t_L g586 ( .A(n_159), .B(n_246), .Y(n_586) );
INVxp67_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_165), .B(n_269), .Y(n_496) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g362 ( .A(n_167), .B(n_254), .Y(n_362) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_181), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_169), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_169), .B(n_246), .Y(n_624) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
INVx2_ASAP7_75t_SL g197 ( .A(n_174), .Y(n_197) );
INVx2_ASAP7_75t_L g259 ( .A(n_174), .Y(n_259) );
INVx1_ASAP7_75t_L g645 ( .A(n_174), .Y(n_645) );
INVx2_ASAP7_75t_L g655 ( .A(n_174), .Y(n_655) );
INVx1_ASAP7_75t_L g671 ( .A(n_174), .Y(n_671) );
INVx1_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_179), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_179), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g565 ( .A(n_179), .Y(n_565) );
INVx2_ASAP7_75t_L g584 ( .A(n_179), .Y(n_584) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx2_ASAP7_75t_L g214 ( .A(n_183), .Y(n_214) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
NOR2xp33_ASAP7_75t_SL g267 ( .A(n_185), .B(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_201), .Y(n_187) );
AND2x4_ASAP7_75t_L g280 ( .A(n_188), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g364 ( .A(n_189), .B(n_333), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_189), .B(n_358), .Y(n_448) );
OR2x2_ASAP7_75t_L g481 ( .A(n_189), .B(n_398), .Y(n_481) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g317 ( .A(n_190), .Y(n_317) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_199), .Y(n_190) );
INVx1_ASAP7_75t_L g245 ( .A(n_192), .Y(n_245) );
OA22x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_198), .Y(n_192) );
INVx4_ASAP7_75t_L g560 ( .A(n_193), .Y(n_560) );
INVx1_ASAP7_75t_L g257 ( .A(n_196), .Y(n_257) );
INVx3_ASAP7_75t_L g557 ( .A(n_196), .Y(n_557) );
INVx1_ASAP7_75t_L g248 ( .A(n_199), .Y(n_248) );
INVx2_ASAP7_75t_L g568 ( .A(n_200), .Y(n_568) );
BUFx2_ASAP7_75t_SL g345 ( .A(n_201), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
INVx1_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g282 ( .A(n_203), .Y(n_282) );
INVx3_ASAP7_75t_L g319 ( .A(n_203), .Y(n_319) );
AND2x2_ASAP7_75t_L g354 ( .A(n_203), .B(n_320), .Y(n_354) );
AND2x2_ASAP7_75t_L g454 ( .A(n_203), .B(n_223), .Y(n_454) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
INVx3_ASAP7_75t_L g566 ( .A(n_210), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
INVx2_ASAP7_75t_L g249 ( .A(n_213), .Y(n_249) );
INVx2_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_213) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_320) );
INVx1_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
AND2x2_ASAP7_75t_L g301 ( .A(n_223), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g327 ( .A(n_223), .B(n_282), .Y(n_327) );
INVx2_ASAP7_75t_L g333 ( .A(n_223), .Y(n_333) );
AND2x2_ASAP7_75t_L g358 ( .A(n_223), .B(n_319), .Y(n_358) );
BUFx2_ASAP7_75t_L g388 ( .A(n_223), .Y(n_388) );
INVx2_ASAP7_75t_L g399 ( .A(n_223), .Y(n_399) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_236), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_231), .B(n_232), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_231), .A2(n_641), .B(n_642), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_250), .B1(n_272), .B2(n_279), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g339 ( .A(n_243), .B(n_332), .Y(n_339) );
INVx2_ASAP7_75t_SL g394 ( .A(n_243), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_243), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
OR2x2_ASAP7_75t_L g325 ( .A(n_244), .B(n_320), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_248), .Y(n_244) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g281 ( .A(n_249), .B(n_282), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_250), .B(n_306), .C(n_310), .Y(n_305) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_269), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g298 ( .A(n_254), .B(n_290), .Y(n_298) );
INVx1_ASAP7_75t_L g309 ( .A(n_254), .Y(n_309) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
OR2x2_ASAP7_75t_L g342 ( .A(n_254), .B(n_290), .Y(n_342) );
INVx1_ASAP7_75t_L g416 ( .A(n_254), .Y(n_416) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_254), .Y(n_501) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_261), .A3(n_266), .B(n_267), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_259), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_263), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
OR2x2_ASAP7_75t_L g328 ( .A(n_269), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g340 ( .A(n_270), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g349 ( .A(n_270), .B(n_298), .Y(n_349) );
AND2x4_ASAP7_75t_L g455 ( .A(n_270), .B(n_362), .Y(n_455) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g391 ( .A(n_275), .B(n_313), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_276), .B(n_290), .Y(n_432) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g417 ( .A(n_277), .B(n_380), .Y(n_417) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_277), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_279), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g424 ( .A(n_280), .B(n_375), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_281), .B(n_388), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_281), .B(n_429), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_281), .B(n_364), .Y(n_485) );
AND2x2_ASAP7_75t_L g347 ( .A(n_282), .B(n_317), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_297), .B(n_299), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x2_ASAP7_75t_L g307 ( .A(n_286), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_286), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_286), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g458 ( .A(n_286), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g395 ( .A(n_288), .Y(n_395) );
INVx1_ASAP7_75t_L g505 ( .A(n_289), .Y(n_505) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_309), .Y(n_308) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_290), .Y(n_464) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g380 ( .A(n_292), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_298), .B(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_298), .Y(n_402) );
AOI22xp5_ASAP7_75t_SL g450 ( .A1(n_299), .A2(n_451), .B1(n_452), .B2(n_455), .Y(n_450) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_338), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_314), .B(n_321), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
OR2x2_ASAP7_75t_L g378 ( .A(n_309), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g490 ( .A(n_309), .B(n_408), .Y(n_490) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_310), .Y(n_451) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
OR2x2_ASAP7_75t_L g421 ( .A(n_315), .B(n_327), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_315), .A2(n_454), .B(n_457), .C(n_460), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_315), .B(n_318), .Y(n_493) );
AND2x2_ASAP7_75t_L g506 ( .A(n_315), .B(n_354), .Y(n_506) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g374 ( .A(n_316), .B(n_318), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_316), .B(n_354), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_316), .B(n_358), .Y(n_477) );
AND2x2_ASAP7_75t_L g482 ( .A(n_316), .B(n_454), .Y(n_482) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g441 ( .A(n_317), .Y(n_441) );
AND2x2_ASAP7_75t_L g488 ( .A(n_317), .B(n_320), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_318), .B(n_388), .Y(n_420) );
AND2x2_ASAP7_75t_L g465 ( .A(n_318), .B(n_364), .Y(n_465) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_319), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g440 ( .A(n_320), .B(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_328), .B1(n_330), .B2(n_334), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AND2x2_ASAP7_75t_L g331 ( .A(n_324), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_324), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g356 ( .A(n_325), .Y(n_356) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g385 ( .A(n_333), .B(n_354), .Y(n_385) );
INVx1_ASAP7_75t_L g430 ( .A(n_333), .Y(n_430) );
AND2x2_ASAP7_75t_L g468 ( .A(n_333), .B(n_347), .Y(n_468) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_335), .A2(n_435), .B1(n_480), .B2(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g370 ( .A(n_337), .Y(n_370) );
AOI211xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_340), .B(n_343), .C(n_350), .Y(n_338) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_340), .B(n_405), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_341), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_348), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI332xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .A3(n_353), .B1(n_355), .B2(n_357), .B3(n_359), .C1(n_361), .C2(n_363), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_354), .A2(n_405), .B1(n_409), .B2(n_410), .Y(n_404) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_355), .Y(n_409) );
INVx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g503 ( .A(n_357), .Y(n_503) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g431 ( .A(n_360), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g504 ( .A(n_360), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g459 ( .A(n_362), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_362), .B(n_446), .Y(n_460) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_403), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_371), .B(n_376), .C(n_392), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g486 ( .A(n_375), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_385), .B1(n_386), .B2(n_389), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_378), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g500 ( .A(n_379), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g423 ( .A(n_380), .Y(n_423) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_384), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g602 ( .A(n_384), .Y(n_602) );
INVx1_ASAP7_75t_L g469 ( .A(n_385), .Y(n_469) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI32xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_400), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI321xp33_ASAP7_75t_L g494 ( .A1(n_396), .A2(n_409), .A3(n_439), .B1(n_495), .B2(n_497), .C(n_502), .Y(n_494) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND3xp33_ASAP7_75t_SL g403 ( .A(n_404), .B(n_412), .C(n_425), .Y(n_403) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g410 ( .A(n_408), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_408), .A2(n_503), .B1(n_504), .B2(n_506), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_418), .B1(n_422), .B2(n_424), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2x1p5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_417), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .C(n_421), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_421), .A2(n_476), .B(n_478), .C(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND4x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_450), .C(n_456), .D(n_461), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_442), .B(n_443), .C(n_449), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_459), .A2(n_467), .B(n_469), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B(n_466), .C(n_470), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .C(n_494), .Y(n_474) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B(n_489), .C(n_491), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_520), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_509), .B(n_521), .Y(n_525) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx8_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx12f_ASAP7_75t_L g528 ( .A(n_512), .Y(n_528) );
INVx2_ASAP7_75t_SL g541 ( .A(n_512), .Y(n_541) );
BUFx6f_ASAP7_75t_L g961 ( .A(n_512), .Y(n_961) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OR2x6_ASAP7_75t_L g928 ( .A(n_515), .B(n_929), .Y(n_928) );
INVx8_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g933 ( .A(n_516), .B(n_934), .Y(n_933) );
OR2x6_ASAP7_75t_L g952 ( .A(n_516), .B(n_934), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_522), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_522), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_524), .B(n_954), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_SL g531 ( .A(n_532), .B(n_535), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_532), .B(n_544), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
OA21x2_ASAP7_75t_L g956 ( .A1(n_533), .A2(n_957), .B(n_959), .Y(n_956) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
CKINVDCx6p67_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_537), .Y(n_544) );
OAI21xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_545), .B(n_953), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_935), .B1(n_942), .B2(n_943), .C(n_948), .Y(n_545) );
OAI22x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_925), .B1(n_930), .B2(n_931), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g945 ( .A(n_548), .Y(n_945) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_815), .Y(n_548) );
NAND4xp25_ASAP7_75t_L g549 ( .A(n_550), .B(n_741), .C(n_775), .D(n_784), .Y(n_549) );
O2A1O1Ixp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_616), .B(n_632), .C(n_684), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_573), .Y(n_551) );
INVxp67_ASAP7_75t_L g749 ( .A(n_552), .Y(n_749) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_619), .Y(n_618) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_553), .B(n_631), .Y(n_764) );
NOR2x1_ASAP7_75t_L g773 ( .A(n_553), .B(n_623), .Y(n_773) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g712 ( .A(n_554), .Y(n_712) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_561), .B(n_571), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_557), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_560), .B(n_582), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_566), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_566), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AOI21x1_ASAP7_75t_L g619 ( .A1(n_568), .A2(n_620), .B(n_621), .Y(n_619) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_569), .A2(n_640), .B(n_643), .Y(n_639) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_570), .A2(n_638), .B(n_679), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g818 ( .A1(n_573), .A2(n_760), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g822 ( .A(n_573), .Y(n_822) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_588), .Y(n_573) );
INVx1_ASAP7_75t_L g732 ( .A(n_574), .Y(n_732) );
AND2x6_ASAP7_75t_SL g747 ( .A(n_574), .B(n_618), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_574), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_574), .B(n_773), .Y(n_772) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_575), .B(n_604), .Y(n_707) );
AND2x2_ASAP7_75t_L g852 ( .A(n_575), .B(n_589), .Y(n_852) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g631 ( .A(n_576), .Y(n_631) );
AO31x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .A3(n_586), .B(n_587), .Y(n_576) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g676 ( .A(n_585), .Y(n_676) );
INVx1_ASAP7_75t_L g867 ( .A(n_588), .Y(n_867) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_603), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_589), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g752 ( .A(n_589), .Y(n_752) );
AND2x4_ASAP7_75t_L g778 ( .A(n_589), .B(n_630), .Y(n_778) );
INVx1_ASAP7_75t_L g788 ( .A(n_589), .Y(n_788) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_590), .Y(n_629) );
INVx1_ASAP7_75t_L g605 ( .A(n_591), .Y(n_605) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_597), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g660 ( .A(n_597), .Y(n_660) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_599), .Y(n_628) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g731 ( .A(n_604), .B(n_718), .Y(n_731) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_604), .Y(n_740) );
INVx1_ASAP7_75t_L g907 ( .A(n_604), .Y(n_907) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_615), .Y(n_604) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_605), .A2(n_639), .B(n_648), .Y(n_729) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_607), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_611), .A2(n_659), .B(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g621 ( .A(n_615), .Y(n_621) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .Y(n_617) );
AND2x2_ASAP7_75t_L g838 ( .A(n_618), .B(n_757), .Y(n_838) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_618), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_618), .B(n_901), .Y(n_900) );
OR2x2_ASAP7_75t_L g717 ( .A(n_619), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g809 ( .A(n_619), .Y(n_809) );
AND2x2_ASAP7_75t_L g738 ( .A(n_622), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g761 ( .A(n_622), .B(n_749), .Y(n_761) );
AND2x4_ASAP7_75t_L g924 ( .A(n_622), .B(n_777), .Y(n_924) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_630), .Y(n_622) );
AND2x4_ASAP7_75t_L g758 ( .A(n_623), .B(n_718), .Y(n_758) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_623), .Y(n_904) );
OA21x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_629), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g716 ( .A(n_630), .Y(n_716) );
BUFx2_ASAP7_75t_SL g757 ( .A(n_630), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_630), .B(n_809), .Y(n_889) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_632), .A2(n_758), .B1(n_776), .B2(n_779), .C(n_782), .Y(n_775) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_634), .B(n_649), .Y(n_633) );
INVx2_ASAP7_75t_L g781 ( .A(n_634), .Y(n_781) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g794 ( .A(n_635), .B(n_727), .Y(n_794) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_635), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_635), .B(n_665), .Y(n_836) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g755 ( .A(n_636), .B(n_666), .Y(n_755) );
AND2x2_ASAP7_75t_L g798 ( .A(n_636), .B(n_650), .Y(n_798) );
AND2x2_ASAP7_75t_L g873 ( .A(n_636), .B(n_737), .Y(n_873) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI21x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_648), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_647), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_647), .A2(n_693), .B(n_696), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_649), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_665), .Y(n_649) );
INVx2_ASAP7_75t_SL g722 ( .A(n_650), .Y(n_722) );
BUFx2_ASAP7_75t_L g901 ( .A(n_650), .Y(n_901) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g688 ( .A(n_651), .Y(n_688) );
INVx3_ASAP7_75t_L g730 ( .A(n_651), .Y(n_730) );
OA21x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_658), .B(n_664), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g689 ( .A(n_665), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g859 ( .A(n_665), .B(n_690), .Y(n_859) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g745 ( .A(n_666), .B(n_729), .Y(n_745) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_674), .B(n_683), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_667), .A2(n_674), .B(n_683), .Y(n_724) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_670), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND3x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .C(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_704), .B(n_713), .C(n_725), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
AND2x2_ASAP7_75t_L g834 ( .A(n_687), .B(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_687), .B(n_854), .Y(n_853) );
OR2x2_ASAP7_75t_L g858 ( .A(n_687), .B(n_859), .Y(n_858) );
INVx2_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g803 ( .A(n_688), .Y(n_803) );
INVx2_ASAP7_75t_L g774 ( .A(n_689), .Y(n_774) );
AND2x2_ASAP7_75t_L g780 ( .A(n_689), .B(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_689), .B(n_803), .Y(n_802) );
OAI322xp33_ASAP7_75t_L g830 ( .A1(n_689), .A2(n_760), .A3(n_831), .B1(n_833), .B2(n_837), .C1(n_839), .C2(n_845), .Y(n_830) );
AND2x2_ASAP7_75t_L g918 ( .A(n_689), .B(n_873), .Y(n_918) );
OR2x2_ASAP7_75t_L g723 ( .A(n_690), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_690), .Y(n_727) );
INVx1_ASAP7_75t_L g735 ( .A(n_690), .Y(n_735) );
AND2x2_ASAP7_75t_L g909 ( .A(n_690), .B(n_724), .Y(n_909) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_690), .Y(n_921) );
AO31x2_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .A3(n_697), .B(n_702), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g808 ( .A(n_711), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g814 ( .A(n_711), .Y(n_814) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_711), .Y(n_913) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g718 ( .A(n_712), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_719), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g746 ( .A(n_714), .B(n_747), .C(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
AND2x2_ASAP7_75t_L g807 ( .A(n_716), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g877 ( .A(n_716), .Y(n_877) );
INVx2_ASAP7_75t_L g777 ( .A(n_717), .Y(n_777) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
AND2x2_ASAP7_75t_L g923 ( .A(n_721), .B(n_755), .Y(n_923) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g754 ( .A(n_722), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g779 ( .A(n_722), .B(n_780), .Y(n_779) );
OR2x2_ASAP7_75t_L g829 ( .A(n_722), .B(n_723), .Y(n_829) );
NOR3xp33_ASAP7_75t_L g903 ( .A(n_722), .B(n_877), .C(n_904), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_723), .A2(n_818), .B(n_820), .Y(n_817) );
OAI31xp33_ASAP7_75t_L g821 ( .A1(n_723), .A2(n_822), .A3(n_823), .B(n_824), .Y(n_821) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_731), .A3(n_732), .B1(n_733), .B2(n_738), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
AND2x2_ASAP7_75t_L g791 ( .A(n_727), .B(n_737), .Y(n_791) );
INVx1_ASAP7_75t_L g843 ( .A(n_727), .Y(n_843) );
INVx1_ASAP7_75t_L g855 ( .A(n_727), .Y(n_855) );
AND2x2_ASAP7_75t_L g868 ( .A(n_727), .B(n_755), .Y(n_868) );
INVx1_ASAP7_75t_L g872 ( .A(n_727), .Y(n_872) );
OR2x2_ASAP7_75t_L g875 ( .A(n_727), .B(n_841), .Y(n_875) );
INVx1_ASAP7_75t_L g765 ( .A(n_728), .Y(n_765) );
INVx1_ASAP7_75t_L g896 ( .A(n_728), .Y(n_896) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g736 ( .A(n_729), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_730), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_730), .B(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g800 ( .A(n_731), .Y(n_800) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g744 ( .A(n_735), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g895 ( .A(n_735), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g760 ( .A(n_736), .Y(n_760) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_736), .Y(n_823) );
AND2x2_ASAP7_75t_L g793 ( .A(n_737), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g804 ( .A(n_738), .Y(n_804) );
INVx1_ASAP7_75t_L g851 ( .A(n_739), .Y(n_851) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g770 ( .A(n_740), .Y(n_770) );
NOR2x1p5_ASAP7_75t_L g827 ( .A(n_740), .B(n_764), .Y(n_827) );
NAND2x1p5_ASAP7_75t_L g879 ( .A(n_740), .B(n_758), .Y(n_879) );
NOR2xp33_ASAP7_75t_SL g741 ( .A(n_742), .B(n_762), .Y(n_741) );
OAI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B(n_753), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_744), .B(n_756), .Y(n_783) );
AND2x2_ASAP7_75t_L g790 ( .A(n_745), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g854 ( .A(n_745), .B(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_745), .B(n_803), .Y(n_874) );
INVx1_ASAP7_75t_L g824 ( .A(n_747), .Y(n_824) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g905 ( .A(n_749), .B(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_751), .B(n_841), .Y(n_844) );
INVx1_ASAP7_75t_L g826 ( .A(n_752), .Y(n_826) );
AND2x2_ASAP7_75t_L g832 ( .A(n_752), .B(n_814), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B1(n_759), .B2(n_761), .Y(n_753) );
OAI21xp5_ASAP7_75t_SL g792 ( .A1(n_754), .A2(n_793), .B(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g841 ( .A(n_755), .Y(n_841) );
AND2x4_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B(n_766), .C(n_774), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g866 ( .A(n_764), .B(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g864 ( .A(n_765), .Y(n_864) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_768), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_768), .B(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g862 ( .A(n_772), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_773), .A2(n_864), .B1(n_865), .B2(n_868), .Y(n_863) );
AND2x2_ASAP7_75t_L g887 ( .A(n_773), .B(n_888), .Y(n_887) );
AND2x4_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_778), .Y(n_795) );
INVx2_ASAP7_75t_SL g801 ( .A(n_778), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_778), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g912 ( .A(n_778), .B(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g820 ( .A(n_780), .Y(n_820) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI211xp5_ASAP7_75t_SL g784 ( .A1(n_785), .A2(n_786), .B(n_796), .C(n_805), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_789), .B(n_792), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g812 ( .A(n_791), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g922 ( .A1(n_794), .A2(n_923), .B(n_924), .Y(n_922) );
OAI22xp33_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_799), .B1(n_802), .B2(n_804), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g819 ( .A(n_798), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_798), .B(n_915), .Y(n_914) );
NAND2x1_ASAP7_75t_SL g920 ( .A(n_798), .B(n_921), .Y(n_920) );
OR2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_810), .B1(n_812), .B2(n_813), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g882 ( .A(n_808), .Y(n_882) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_812), .B(n_861), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_847), .C(n_890), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_821), .B1(n_825), .B2(n_828), .C(n_830), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_820), .A2(n_881), .B1(n_883), .B2(n_884), .C(n_885), .Y(n_880) );
INVx1_ASAP7_75t_L g892 ( .A(n_825), .Y(n_892) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_827), .Y(n_917) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g884 ( .A(n_832), .Y(n_884) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g861 ( .A(n_835), .Y(n_861) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_838), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
INVx2_ASAP7_75t_SL g883 ( .A(n_840), .Y(n_883) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g886 ( .A(n_841), .Y(n_886) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NOR3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_869), .C(n_880), .Y(n_847) );
OAI211xp5_ASAP7_75t_SL g848 ( .A1(n_849), .A2(n_853), .B(n_856), .C(n_863), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g915 ( .A(n_855), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_860), .B(n_862), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AOI31xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_874), .A3(n_875), .B(n_876), .Y(n_869) );
NAND2xp5_ASAP7_75t_SL g894 ( .A(n_870), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_877), .Y(n_899) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g893 ( .A(n_887), .Y(n_893) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AOI211xp5_ASAP7_75t_SL g890 ( .A1(n_891), .A2(n_894), .B(n_897), .C(n_910), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
O2A1O1Ixp33_ASAP7_75t_SL g897 ( .A1(n_898), .A2(n_900), .B(n_902), .C(n_908), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI211xp5_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_914), .B(n_916), .C(n_922), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_SL g919 ( .A(n_920), .Y(n_919) );
BUFx3_ASAP7_75t_L g947 ( .A(n_925), .Y(n_947) );
BUFx12f_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
CKINVDCx11_ASAP7_75t_R g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AOI22x1_ASAP7_75t_L g944 ( .A1(n_930), .A2(n_932), .B1(n_945), .B2(n_946), .Y(n_944) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_932), .Y(n_931) );
BUFx8_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g942 ( .A(n_935), .Y(n_942) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
BUFx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
CKINVDCx8_ASAP7_75t_R g955 ( .A(n_956), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_958), .Y(n_957) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx5_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
endmodule