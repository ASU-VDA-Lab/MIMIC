module real_jpeg_5684_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_0),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_0),
.A2(n_104),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_0),
.A2(n_104),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_1),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_1),
.Y(n_463)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_2),
.Y(n_153)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_2),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_64),
.B1(n_147),
.B2(n_172),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_64),
.B1(n_162),
.B2(n_230),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_3),
.A2(n_64),
.B1(n_189),
.B2(n_192),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_4),
.A2(n_53),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_4),
.A2(n_53),
.B1(n_286),
.B2(n_359),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_4),
.A2(n_53),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_5),
.Y(n_519)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_7),
.A2(n_254),
.B1(n_256),
.B2(n_260),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_7),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_7),
.B(n_268),
.C(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_7),
.B(n_117),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_7),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_7),
.B(n_97),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_7),
.B(n_235),
.Y(n_349)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_8),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_9),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_9),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_9),
.A2(n_136),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_136),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_12),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_13),
.A2(n_232),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_13),
.A2(n_278),
.B1(n_293),
.B2(n_314),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_13),
.A2(n_293),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_13),
.A2(n_61),
.B1(n_293),
.B2(n_467),
.Y(n_466)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_16),
.A2(n_61),
.B1(n_63),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_16),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_16),
.A2(n_241),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_16),
.A2(n_241),
.B1(n_266),
.B2(n_340),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_16),
.A2(n_146),
.B1(n_241),
.B2(n_353),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_17),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_17),
.A2(n_127),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_17),
.A2(n_103),
.B1(n_127),
.B2(n_195),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_17),
.A2(n_127),
.B1(n_189),
.B2(n_224),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_18),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_18),
.A2(n_82),
.B1(n_163),
.B2(n_201),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_18),
.A2(n_201),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_18),
.A2(n_134),
.B1(n_201),
.B2(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_514),
.B(n_516),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_206),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_205),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_155),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_24),
.B(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_137),
.B2(n_138),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_65),
.C(n_105),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_27),
.A2(n_139),
.B1(n_140),
.B2(n_154),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_27),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_27),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_51),
.B1(n_58),
.B2(n_60),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_28),
.A2(n_58),
.B1(n_60),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_28),
.A2(n_240),
.B(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_28),
.A2(n_58),
.B1(n_240),
.B2(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_29),
.B(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_29),
.A2(n_436),
.B(n_437),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_37),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g413 ( 
.A(n_33),
.Y(n_413)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_40),
.Y(n_415)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_44),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_44),
.Y(n_347)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_44),
.Y(n_354)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_44),
.Y(n_392)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_48),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_48),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_48),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_48),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_52),
.B(n_59),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_54),
.Y(n_411)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_57),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_58),
.B(n_260),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_58),
.A2(n_199),
.B(n_466),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_59),
.B(n_200),
.Y(n_242)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_63),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_65),
.A2(n_66),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_65),
.A2(n_66),
.B1(n_105),
.B2(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_96),
.B(n_98),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_67),
.A2(n_253),
.B(n_261),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_67),
.A2(n_96),
.B1(n_292),
.B2(n_339),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_67),
.A2(n_261),
.B(n_339),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_67),
.A2(n_96),
.B1(n_442),
.B2(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_68),
.A2(n_97),
.B1(n_161),
.B2(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_68),
.A2(n_97),
.B1(n_161),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_68),
.A2(n_97),
.B1(n_194),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_68),
.B(n_262),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_85),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_75),
.B1(n_78),
.B2(n_82),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_73),
.Y(n_259)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_74),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_74),
.Y(n_340)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_86),
.B1(n_90),
.B2(n_93),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_84),
.Y(n_446)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_85),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_88),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_92),
.Y(n_360)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_95),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_96),
.A2(n_297),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_97),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_101),
.Y(n_266)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_123),
.B1(n_130),
.B2(n_131),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_130),
.B1(n_131),
.B2(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_107),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_107),
.A2(n_130),
.B1(n_171),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_107),
.A2(n_130),
.B1(n_387),
.B2(n_440),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_113),
.Y(n_369)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_113),
.Y(n_376)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_124),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22x1_ASAP7_75t_L g470 ( 
.A1(n_117),
.A2(n_169),
.B1(n_394),
.B2(n_471),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_119),
.Y(n_444)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_130),
.B(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_130),
.A2(n_387),
.B(n_393),
.Y(n_386)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g363 ( 
.A1(n_146),
.A2(n_349),
.A3(n_364),
.B1(n_366),
.B2(n_370),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_173),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_159),
.CI(n_173),
.CON(n_208),
.SN(n_208)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_169),
.A2(n_343),
.B(n_350),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_169),
.B(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_169),
.A2(n_350),
.B(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B(n_197),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_193),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_197),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_175),
.A2(n_193),
.B1(n_214),
.B2(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_184),
.B(n_187),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_187),
.B1(n_221),
.B2(n_226),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_176),
.A2(n_274),
.B(n_281),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_176),
.A2(n_260),
.B(n_281),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_176),
.A2(n_425),
.B1(n_426),
.B2(n_428),
.Y(n_424)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_177),
.B(n_284),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_177),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_177),
.A2(n_227),
.B1(n_358),
.B2(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_177),
.A2(n_429),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_182),
.Y(n_286)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_186),
.Y(n_309)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_186),
.Y(n_328)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g288 ( 
.A(n_190),
.Y(n_288)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_193),
.Y(n_455)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g436 ( 
.A1(n_202),
.A2(n_260),
.B(n_419),
.Y(n_436)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_243),
.B(n_513),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_208),
.B(n_209),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_208),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_218),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_215),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_218),
.B(n_473),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_233),
.C(n_239),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_219),
.B(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_220),
.B(n_228),
.Y(n_481)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_221),
.Y(n_461)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_233),
.B(n_239),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_234),
.Y(n_471)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_238),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_242),
.Y(n_437)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI311xp33_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_449),
.A3(n_489),
.B1(n_507),
.C1(n_512),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_401),
.B(n_448),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_378),
.B(n_400),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_333),
.B(n_377),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_300),
.B(n_332),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_272),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_272),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_263),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_252),
.A2(n_263),
.B1(n_264),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_259),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_260),
.A2(n_344),
.B(n_348),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_260),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_289),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_290),
.C(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_298),
.B2(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_323),
.B(n_331),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_311),
.B(n_322),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_321),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_321),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_317),
.B(n_320),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_357),
.B(n_361),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_329),
.Y(n_331)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_335),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_355),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_341),
.C(n_355),
.Y(n_379)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_354),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_363),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_363),
.Y(n_384)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_379),
.B(n_380),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_399),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_384),
.C(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_395),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_396),
.C(n_397),
.Y(n_430)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_403),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_433),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_404)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_423),
.B2(n_424),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_407),
.B(n_423),
.Y(n_485)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_410),
.A3(n_412),
.B1(n_414),
.B2(n_419),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_430),
.B(n_431),
.C(n_433),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_438),
.B2(n_447),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_434),
.B(n_439),
.C(n_441),
.Y(n_498)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_475),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_SL g507 ( 
.A1(n_450),
.A2(n_475),
.B(n_508),
.C(n_511),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_472),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_451),
.B(n_472),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.C(n_456),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_452),
.B(n_454),
.CI(n_456),
.CON(n_488),
.SN(n_488)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_464),
.C(n_470),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_460),
.Y(n_497)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_464),
.A2(n_465),
.B1(n_470),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx8_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_470),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_488),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_481),
.C(n_482),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_477),
.A2(n_478),
.B1(n_481),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_500),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_486),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_483),
.A2(n_484),
.B1(n_486),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_486),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_488),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_502),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_509),
.B(n_510),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_499),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_499),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.C(n_498),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_505),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_497),
.B1(n_498),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_498),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_504),
.Y(n_509)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx13_ASAP7_75t_L g518 ( 
.A(n_515),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_519),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);


endmodule