module real_jpeg_20415_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_25),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_0),
.A2(n_9),
.B1(n_25),
.B2(n_45),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_42),
.B1(n_49),
.B2(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_9),
.B1(n_45),
.B2(n_54),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_54),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_2),
.B(n_27),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_2),
.A2(n_9),
.B(n_14),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_42),
.B1(n_49),
.B2(n_118),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_92),
.B1(n_97),
.B2(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_74),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_30),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_2),
.A2(n_30),
.B(n_205),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_56),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_9),
.B1(n_45),
.B2(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_3),
.A2(n_42),
.B1(n_49),
.B2(n_56),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_4),
.A2(n_9),
.B1(n_45),
.B2(n_113),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_42),
.B1(n_49),
.B2(n_113),
.Y(n_193)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_6),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_42),
.B1(n_49),
.B2(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_9),
.B1(n_45),
.B2(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_45),
.Y(n_93)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_8),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_9),
.B1(n_45),
.B2(n_115),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_8),
.A2(n_42),
.B1(n_49),
.B2(n_115),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_115),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_14),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_9),
.A2(n_11),
.B1(n_33),
.B2(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_11),
.A2(n_33),
.B1(n_42),
.B2(n_49),
.Y(n_102)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_337),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_80),
.B(n_335),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_21),
.A2(n_52),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_22),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_29),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_29),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_23),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_34),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_28),
.A2(n_35),
.B1(n_117),
.B2(n_124),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_28),
.A2(n_42),
.A3(n_64),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_29),
.B(n_30),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_30),
.A2(n_62),
.B(n_63),
.C(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_31),
.A2(n_53),
.B(n_57),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_34),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_37),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_72),
.C(n_76),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_38),
.A2(n_39),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.C(n_58),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_40),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_40),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_40),
.A2(n_58),
.B1(n_59),
.B2(n_311),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_47),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_47),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_41),
.A2(n_44),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_41),
.A2(n_44),
.B1(n_173),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_41),
.A2(n_44),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_41),
.A2(n_212),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_41),
.A2(n_44),
.B1(n_100),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_41),
.A2(n_108),
.B(n_245),
.Y(n_279)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_44),
.B(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_45),
.B(n_182),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_46),
.A2(n_49),
.B(n_118),
.C(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_48),
.B(n_109),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g206 ( 
.A(n_49),
.B(n_63),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_50),
.A2(n_51),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_52),
.A2(n_57),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_52),
.A2(n_57),
.B1(n_131),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_52),
.A2(n_79),
.B(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_67),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_68),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_62),
.A2(n_68),
.B1(n_151),
.B2(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_62),
.B(n_71),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_62),
.A2(n_66),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_62),
.A2(n_68),
.B1(n_270),
.B2(n_291),
.Y(n_290)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_74),
.B(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_74),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_67),
.A2(n_75),
.B(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_67),
.A2(n_256),
.B(n_314),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_76),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_328),
.B(n_334),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_304),
.A3(n_323),
.B1(n_326),
.B2(n_327),
.C(n_340),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_283),
.B(n_303),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_261),
.B(n_282),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_153),
.B(n_236),
.C(n_260),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_136),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_86),
.B(n_136),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_121),
.B2(n_135),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_105),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_89),
.B(n_105),
.C(n_135),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_99),
.B2(n_104),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_90),
.B(n_104),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_92),
.A2(n_145),
.B1(n_162),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_92),
.A2(n_165),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_92),
.A2(n_145),
.B(n_278),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_93),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_93),
.A2(n_96),
.B(n_197),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_118),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_98),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_101),
.B(n_227),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_122),
.B(n_128),
.C(n_133),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_125),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_137),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_149),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_143),
.A2(n_144),
.B1(n_148),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_146),
.B(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_149),
.B(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_235),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_230),
.B(n_234),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_217),
.B(n_229),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_199),
.B(n_216),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_185),
.B(n_198),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_174),
.B(n_184),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_166),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_170),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_197),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_207),
.B1(n_214),
.B2(n_215),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_219),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_226),
.C(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2x2_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_258),
.B2(n_259),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_247),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_247),
.C(n_259),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_275),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_277),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_294),
.B(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_285),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_301),
.B2(n_302),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_293),
.C(n_302),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_306),
.C(n_315),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_292),
.B(n_306),
.CI(n_315),
.CON(n_325),
.SN(n_325)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_321),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_325),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);


endmodule