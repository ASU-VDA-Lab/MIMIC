module fake_jpeg_2686_n_594 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_594);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_594;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_57),
.B(n_64),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_30),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_10),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_10),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_67),
.B(n_108),
.Y(n_166)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_68),
.Y(n_191)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_70),
.B(n_44),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_79),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_86),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_88),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_93),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_115),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_100),
.Y(n_218)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_102),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_45),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_2),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_25),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_2),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_2),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_39),
.Y(n_142)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_135),
.B(n_207),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_143),
.B(n_157),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_56),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_150),
.B(n_159),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_108),
.B(n_26),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_67),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_57),
.B(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_167),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_35),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_88),
.B(n_46),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_168),
.B(n_177),
.Y(n_252)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_70),
.B(n_46),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_83),
.B(n_41),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_41),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_58),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_62),
.Y(n_194)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_71),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_74),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_202),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_66),
.B(n_44),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_119),
.B(n_53),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_78),
.B(n_53),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_92),
.B(n_54),
.C(n_52),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_2),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_79),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_257)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_80),
.Y(n_211)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_81),
.B(n_40),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_214),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_120),
.A2(n_51),
.B1(n_28),
.B2(n_40),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_38),
.B1(n_47),
.B2(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_93),
.B(n_54),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_7),
.Y(n_267)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_219),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_127),
.A2(n_24),
.B1(n_95),
.B2(n_115),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_220),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_153),
.A2(n_24),
.B1(n_51),
.B2(n_38),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_221),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_222),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_224),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_225),
.A2(n_242),
.B1(n_244),
.B2(n_257),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_226),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_205),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_230),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_266),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_235),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_129),
.B(n_3),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_240),
.A2(n_265),
.B1(n_269),
.B2(n_191),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_241),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_182),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_245),
.Y(n_338)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

BUFx24_ASAP7_75t_L g343 ( 
.A(n_248),
.Y(n_343)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_250),
.Y(n_348)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_154),
.Y(n_251)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_138),
.Y(n_254)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_258),
.Y(n_314)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_259),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_260),
.Y(n_322)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_276),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_155),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_267),
.B(n_271),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_128),
.A2(n_130),
.B1(n_152),
.B2(n_139),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_270),
.A2(n_280),
.B1(n_289),
.B2(n_292),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_166),
.B(n_149),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_272),
.B(n_279),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_131),
.B(n_186),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_274),
.B(n_275),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_196),
.B(n_140),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_146),
.B(n_145),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_278),
.Y(n_312)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_180),
.Y(n_279)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_147),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_171),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_282),
.Y(n_316)
);

CKINVDCx9p33_ASAP7_75t_R g282 ( 
.A(n_170),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_171),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_285),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_193),
.B(n_180),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_161),
.B(n_175),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_288),
.Y(n_330)
);

CKINVDCx12_ASAP7_75t_R g288 ( 
.A(n_198),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_189),
.A2(n_198),
.B1(n_193),
.B2(n_218),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_134),
.B(n_144),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_291),
.Y(n_333)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_184),
.Y(n_291)
);

CKINVDCx6p67_ASAP7_75t_R g292 ( 
.A(n_170),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_295),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_216),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_296),
.A2(n_162),
.B1(n_172),
.B2(n_228),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_210),
.A3(n_215),
.B1(n_209),
.B2(n_191),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_297),
.B(n_309),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_225),
.A2(n_148),
.B(n_195),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_303),
.A2(n_292),
.B(n_230),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_234),
.A2(n_213),
.B1(n_192),
.B2(n_181),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_304),
.A2(n_318),
.B1(n_334),
.B2(n_339),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_185),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_311),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_227),
.B(n_237),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_185),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_317),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_231),
.B(n_160),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_240),
.A2(n_160),
.B1(n_213),
.B2(n_181),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_268),
.A2(n_190),
.B1(n_192),
.B2(n_216),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_320),
.A2(n_335),
.B1(n_352),
.B2(n_243),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g323 ( 
.A(n_286),
.B(n_162),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_323),
.B(n_340),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_190),
.B1(n_148),
.B2(n_195),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_238),
.A2(n_162),
.B1(n_147),
.B2(n_172),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_263),
.B1(n_294),
.B2(n_273),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_242),
.A2(n_244),
.B(n_283),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_281),
.A2(n_284),
.B1(n_259),
.B2(n_278),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_344),
.A2(n_292),
.B(n_223),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_265),
.A2(n_289),
.B1(n_232),
.B2(n_275),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_236),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_355),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_252),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_356),
.B(n_366),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_357),
.A2(n_368),
.B(n_324),
.Y(n_413)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_300),
.A2(n_251),
.B1(n_262),
.B2(n_270),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_360),
.A2(n_367),
.B1(n_369),
.B2(n_385),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_298),
.B(n_296),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_376),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_362),
.A2(n_377),
.B1(n_380),
.B2(n_387),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_311),
.A2(n_233),
.B(n_261),
.C(n_247),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_249),
.B1(n_276),
.B2(n_226),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_248),
.B(n_224),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_306),
.A2(n_260),
.B1(n_229),
.B2(n_235),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_219),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_370),
.B(n_371),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_298),
.A2(n_245),
.B(n_293),
.C(n_280),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_310),
.B(n_241),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_374),
.B(n_379),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

INVx3_ASAP7_75t_SL g376 ( 
.A(n_341),
.Y(n_376)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_310),
.B(n_255),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_383),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_298),
.B(n_258),
.Y(n_383)
);

OAI22x1_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_351),
.B1(n_338),
.B2(n_346),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_297),
.A2(n_245),
.B1(n_293),
.B2(n_312),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_323),
.B(n_330),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_325),
.Y(n_423)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_302),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_350),
.C(n_317),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_349),
.C(n_348),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_333),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_392),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_323),
.Y(n_392)
);

INVx11_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_393),
.Y(n_432)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_346),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_307),
.A2(n_321),
.B1(n_309),
.B2(n_303),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_359),
.B1(n_392),
.B2(n_371),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_SL g397 ( 
.A1(n_359),
.A2(n_316),
.B(n_352),
.C(n_338),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_397),
.A2(n_413),
.B(n_403),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_398),
.B(n_402),
.C(n_405),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_342),
.C(n_319),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_403),
.B(n_423),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_388),
.C(n_356),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_319),
.C(n_304),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_409),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_342),
.C(n_299),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_391),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_424),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_359),
.A2(n_318),
.B1(n_314),
.B2(n_328),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_415),
.A2(n_369),
.B1(n_386),
.B2(n_361),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_373),
.C(n_366),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_418),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_331),
.B1(n_393),
.B2(n_315),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_426),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_299),
.C(n_351),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_314),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_384),
.A2(n_320),
.B1(n_328),
.B2(n_346),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_427),
.A2(n_358),
.B1(n_387),
.B2(n_372),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_395),
.A2(n_343),
.B(n_315),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_331),
.Y(n_463)
);

AO21x1_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_459),
.B(n_463),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_445),
.B1(n_453),
.B2(n_458),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_461),
.Y(n_476)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_418),
.B(n_383),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_442),
.Y(n_473)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_374),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_360),
.B1(n_364),
.B2(n_389),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_443),
.A2(n_446),
.B1(n_462),
.B2(n_401),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_357),
.B1(n_361),
.B2(n_364),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_354),
.B1(n_394),
.B2(n_368),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_353),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_451),
.Y(n_467)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_430),
.Y(n_449)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_325),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_460),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_419),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_399),
.A2(n_376),
.B1(n_380),
.B2(n_341),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_454),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_425),
.B(n_406),
.Y(n_455)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_455),
.Y(n_494)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_412),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_464),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_399),
.A2(n_376),
.B1(n_375),
.B2(n_301),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_413),
.A2(n_343),
.B(n_377),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_345),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_420),
.A2(n_322),
.B1(n_332),
.B2(n_345),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_411),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_411),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_465),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_433),
.A2(n_456),
.B(n_446),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_466),
.A2(n_468),
.B(n_483),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_456),
.A2(n_397),
.B(n_405),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_402),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_471),
.C(n_472),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_398),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_409),
.C(n_423),
.Y(n_472)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_477),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_410),
.C(n_424),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_489),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_408),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_428),
.B(n_401),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_486),
.B(n_491),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_459),
.A2(n_463),
.B(n_445),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_443),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_412),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_434),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_490),
.B(n_434),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_437),
.A2(n_401),
.B(n_422),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_441),
.B(n_431),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_438),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_473),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_496),
.B(n_500),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_494),
.A2(n_455),
.B1(n_463),
.B2(n_462),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_511),
.B1(n_513),
.B2(n_515),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_475),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_518),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_473),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_508),
.Y(n_529)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_467),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_482),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_512),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_488),
.A2(n_458),
.B1(n_453),
.B2(n_436),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_514),
.A2(n_485),
.B1(n_486),
.B2(n_476),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_435),
.B1(n_464),
.B2(n_465),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_467),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_517),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_471),
.B(n_442),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_470),
.B(n_457),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_476),
.A2(n_431),
.B1(n_454),
.B2(n_449),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_485),
.B1(n_487),
.B2(n_474),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_514),
.A2(n_501),
.B1(n_513),
.B2(n_476),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_521),
.A2(n_528),
.B1(n_531),
.B2(n_502),
.Y(n_548)
);

OAI21xp33_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_472),
.B(n_478),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_524),
.B(n_525),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_489),
.C(n_468),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_495),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_534),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_491),
.C(n_493),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_535),
.C(n_509),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_483),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_469),
.C(n_484),
.Y(n_535)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_538),
.Y(n_558)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_529),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_539),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_534),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_541),
.Y(n_564)
);

BUFx12_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_522),
.C(n_504),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_530),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_544),
.A2(n_548),
.B1(n_551),
.B2(n_552),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_502),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_547),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_536),
.Y(n_547)
);

INVx13_ASAP7_75t_L g549 ( 
.A(n_520),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_550),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_535),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_510),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_499),
.B(n_515),
.Y(n_552)
);

MAJx2_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_548),
.C(n_479),
.Y(n_560)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_553),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_525),
.C(n_532),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_559),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_547),
.A2(n_479),
.B(n_519),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_555),
.B(n_565),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_528),
.C(n_520),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_551),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_563),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_514),
.C(n_510),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_503),
.C(n_523),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_SL g566 ( 
.A(n_564),
.B(n_546),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_567),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_564),
.B(n_558),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_556),
.B(n_542),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_571),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_556),
.B(n_542),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_575),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_562),
.B(n_543),
.C(n_523),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_572),
.B(n_562),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_576),
.B(n_573),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_570),
.A2(n_543),
.B(n_557),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_577),
.A2(n_578),
.B(n_579),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_575),
.B(n_557),
.Y(n_578)
);

AOI31xp67_ASAP7_75t_L g579 ( 
.A1(n_568),
.A2(n_560),
.A3(n_511),
.B(n_507),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_578),
.Y(n_583)
);

AOI21xp33_ASAP7_75t_L g588 ( 
.A1(n_583),
.A2(n_584),
.B(n_586),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_580),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_585),
.B(n_574),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_587),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_588),
.C(n_549),
.Y(n_590)
);

NAND4xp25_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_492),
.C(n_448),
.D(n_461),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_432),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_322),
.C(n_421),
.Y(n_593)
);

AOI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_593),
.A2(n_421),
.B(n_332),
.Y(n_594)
);


endmodule