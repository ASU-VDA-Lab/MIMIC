module real_aes_4389_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_1404;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_0), .A2(n_292), .B1(n_557), .B2(n_558), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_1), .A2(n_6), .B1(n_905), .B2(n_906), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_2), .A2(n_62), .B1(n_515), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_3), .A2(n_217), .B1(n_554), .B2(n_555), .Y(n_1050) );
AOI22xp5_ASAP7_75t_L g989 ( .A1(n_4), .A2(n_225), .B1(n_622), .B2(n_650), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_5), .A2(n_168), .B1(n_547), .B2(n_548), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_7), .A2(n_288), .B1(n_576), .B2(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_8), .A2(n_362), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g598 ( .A(n_9), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g1235 ( .A(n_10), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_11), .A2(n_104), .B1(n_495), .B2(n_515), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_12), .A2(n_186), .B1(n_696), .B2(n_724), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_13), .A2(n_49), .B1(n_507), .B2(n_580), .Y(n_579) );
AOI21x1_ASAP7_75t_L g591 ( .A1(n_14), .A2(n_592), .B(n_597), .Y(n_591) );
INVx1_ASAP7_75t_L g758 ( .A(n_15), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_16), .A2(n_375), .B1(n_500), .B2(n_782), .Y(n_829) );
INVx1_ASAP7_75t_L g777 ( .A(n_17), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_18), .A2(n_342), .B1(n_457), .B2(n_709), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_19), .A2(n_36), .B1(n_582), .B2(n_705), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_20), .A2(n_106), .B1(n_500), .B2(n_694), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_21), .A2(n_117), .B1(n_513), .B2(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_22), .B(n_439), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_23), .A2(n_220), .B1(n_457), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_24), .A2(n_296), .B1(n_909), .B2(n_910), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_25), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_26), .A2(n_274), .B1(n_547), .B2(n_548), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_27), .A2(n_189), .B1(n_576), .B2(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_28), .A2(n_232), .B1(n_550), .B2(n_551), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_29), .B(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_30), .A2(n_263), .B1(n_502), .B2(n_625), .Y(n_784) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_31), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_32), .A2(n_380), .B1(n_589), .B2(n_771), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_33), .A2(n_77), .B1(n_684), .B2(n_685), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_34), .A2(n_167), .B1(n_515), .B2(n_574), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_35), .A2(n_46), .B1(n_912), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g720 ( .A(n_37), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_38), .A2(n_710), .B(n_865), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_39), .A2(n_305), .B1(n_622), .B2(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_40), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g866 ( .A(n_41), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_42), .A2(n_231), .B1(n_704), .B2(n_705), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_43), .A2(n_417), .B1(n_550), .B2(n_551), .Y(n_1003) );
XOR2x2_ASAP7_75t_L g639 ( .A(n_44), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_44), .A2(n_182), .B1(n_1128), .B2(n_1130), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_45), .A2(n_404), .B1(n_655), .B2(n_771), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_47), .A2(n_55), .B1(n_704), .B2(n_705), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_48), .A2(n_164), .B1(n_500), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g892 ( .A(n_50), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_51), .A2(n_177), .B1(n_433), .B2(n_979), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_52), .A2(n_145), .B1(n_457), .B2(n_629), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_53), .A2(n_355), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g1085 ( .A(n_54), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_56), .A2(n_156), .B1(n_625), .B2(n_831), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_57), .A2(n_183), .B1(n_488), .B2(n_495), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_58), .A2(n_201), .B1(n_615), .B2(n_861), .Y(n_888) );
OA22x2_ASAP7_75t_L g454 ( .A1(n_59), .A2(n_180), .B1(n_439), .B2(n_453), .Y(n_454) );
INVx1_ASAP7_75t_L g463 ( .A(n_59), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_60), .A2(n_345), .B1(n_574), .B2(n_786), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_61), .A2(n_71), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_63), .A2(n_65), .B1(n_547), .B2(n_548), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_64), .A2(n_336), .B1(n_622), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_66), .A2(n_401), .B1(n_477), .B2(n_775), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_67), .A2(n_290), .B1(n_488), .B2(n_502), .Y(n_974) );
INVx1_ASAP7_75t_L g1150 ( .A(n_68), .Y(n_1150) );
XOR2x2_ASAP7_75t_L g570 ( .A(n_69), .B(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_69), .A2(n_171), .B1(n_1141), .B2(n_1149), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_70), .A2(n_282), .B1(n_657), .B2(n_658), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_72), .A2(n_341), .B1(n_547), .B2(n_548), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_73), .A2(n_293), .B1(n_782), .B2(n_886), .Y(n_973) );
INVx1_ASAP7_75t_L g455 ( .A(n_74), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_75), .A2(n_114), .B1(n_650), .B2(n_886), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_76), .A2(n_295), .B1(n_550), .B2(n_551), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_78), .A2(n_209), .B1(n_642), .B2(n_643), .C(n_645), .Y(n_641) );
INVx1_ASAP7_75t_SL g1152 ( .A(n_79), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_79), .A2(n_1391), .B1(n_1411), .B2(n_1413), .Y(n_1390) );
INVx1_ASAP7_75t_L g452 ( .A(n_80), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_80), .A2(n_180), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_80), .B(n_203), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_81), .A2(n_472), .B(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g1403 ( .A1(n_82), .A2(n_169), .B1(n_433), .B2(n_1404), .Y(n_1403) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_83), .A2(n_352), .B1(n_472), .B2(n_634), .C(n_636), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_84), .A2(n_395), .B1(n_547), .B2(n_548), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_85), .A2(n_338), .B1(n_655), .B2(n_657), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_86), .A2(n_134), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_87), .A2(n_159), .B1(n_515), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_88), .A2(n_307), .B1(n_576), .B2(n_577), .Y(n_726) );
INVx1_ASAP7_75t_L g820 ( .A(n_89), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_90), .A2(n_126), .B1(n_1121), .B2(n_1125), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_91), .A2(n_207), .B1(n_618), .B2(n_692), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_92), .A2(n_170), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g727 ( .A1(n_93), .A2(n_242), .B1(n_515), .B2(n_692), .Y(n_727) );
INVx1_ASAP7_75t_L g982 ( .A(n_94), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_95), .A2(n_137), .B1(n_704), .B2(n_705), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_96), .B(n_779), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_97), .B(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_98), .A2(n_388), .B1(n_518), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g1123 ( .A(n_99), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_99), .B(n_304), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_100), .A2(n_356), .B1(n_550), .B2(n_551), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_101), .A2(n_267), .B1(n_512), .B2(n_515), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_102), .A2(n_228), .B1(n_543), .B2(n_689), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_103), .A2(n_361), .B1(n_1121), .B2(n_1138), .Y(n_1143) );
INVx1_ASAP7_75t_L g843 ( .A(n_105), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_107), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_108), .A2(n_109), .B1(n_507), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_110), .A2(n_219), .B1(n_541), .B2(n_658), .Y(n_999) );
INVx1_ASAP7_75t_L g926 ( .A(n_111), .Y(n_926) );
AO22x2_ASAP7_75t_L g1166 ( .A1(n_112), .A2(n_335), .B1(n_1121), .B2(n_1138), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_113), .A2(n_115), .B1(n_518), .B2(n_839), .C(n_841), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_116), .A2(n_654), .B(n_891), .Y(n_890) );
XNOR2x1_ASAP7_75t_L g428 ( .A(n_118), .B(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_118), .A2(n_152), .B1(n_1149), .B2(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1381 ( .A(n_119), .Y(n_1381) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_120), .A2(n_839), .B(n_996), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_121), .B(n_1061), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1127 ( .A1(n_122), .A2(n_154), .B1(n_1128), .B2(n_1130), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_123), .A2(n_172), .B1(n_615), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_124), .A2(n_202), .B1(n_655), .B2(n_658), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_125), .A2(n_161), .B1(n_856), .B2(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g842 ( .A(n_127), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_128), .A2(n_151), .B1(n_574), .B2(n_786), .Y(n_970) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_129), .B(n_1109), .Y(n_1124) );
INVx1_ASAP7_75t_SL g1129 ( .A(n_129), .Y(n_1129) );
INVx1_ASAP7_75t_L g1132 ( .A(n_129), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_130), .A2(n_291), .B1(n_457), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_131), .A2(n_195), .B1(n_1090), .B2(n_1092), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_132), .B(n_804), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_133), .A2(n_327), .B1(n_856), .B2(n_857), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_135), .A2(n_215), .B1(n_562), .B2(n_1402), .Y(n_1401) );
XNOR2x1_ASAP7_75t_L g741 ( .A(n_136), .B(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_138), .A2(n_314), .B1(n_577), .B2(n_857), .Y(n_1024) );
INVx1_ASAP7_75t_L g560 ( .A(n_139), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_140), .B(n_634), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_141), .A2(n_297), .B1(n_502), .B2(n_625), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_142), .A2(n_163), .B1(n_1121), .B2(n_1138), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_143), .A2(n_387), .B1(n_696), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_144), .A2(n_398), .B1(n_654), .B2(n_657), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_146), .A2(n_408), .B1(n_643), .B2(n_762), .C(n_763), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g1162 ( .A1(n_147), .A2(n_419), .B1(n_1121), .B2(n_1141), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_148), .A2(n_320), .B1(n_457), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_149), .A2(n_166), .B1(n_500), .B2(n_650), .Y(n_1407) );
XNOR2x1_ASAP7_75t_L g986 ( .A(n_150), .B(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_153), .A2(n_223), .B1(n_433), .B2(n_472), .Y(n_805) );
OAI22x1_ASAP7_75t_L g673 ( .A1(n_154), .A2(n_674), .B1(n_712), .B2(n_713), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_154), .B(n_690), .C(n_706), .Y(n_712) );
INVx1_ASAP7_75t_L g993 ( .A(n_155), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_157), .A2(n_198), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_158), .A2(n_405), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g1063 ( .A1(n_160), .A2(n_472), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g752 ( .A(n_162), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_165), .A2(n_193), .B1(n_577), .B2(n_1077), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_173), .A2(n_248), .B1(n_433), .B2(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_174), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g637 ( .A(n_175), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_176), .A2(n_257), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_178), .A2(n_391), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g446 ( .A(n_179), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_179), .B(n_246), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_179), .B(n_461), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_180), .B(n_319), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_181), .A2(n_256), .B1(n_509), .B2(n_615), .Y(n_783) );
INVx1_ASAP7_75t_L g733 ( .A(n_184), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_185), .A2(n_309), .B1(n_709), .B2(n_773), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_187), .A2(n_289), .B1(n_477), .B2(n_527), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_188), .A2(n_204), .B1(n_518), .B2(n_520), .C(n_524), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_190), .A2(n_269), .B1(n_509), .B2(n_615), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_191), .A2(n_344), .B1(n_509), .B2(n_615), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_192), .A2(n_351), .B1(n_912), .B2(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g1065 ( .A(n_194), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_196), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_197), .A2(n_596), .B(n_1040), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_199), .B(n_804), .Y(n_803) );
AOI21xp33_ASAP7_75t_L g1372 ( .A1(n_200), .A2(n_472), .B(n_1373), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_203), .B(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_205), .A2(n_239), .B1(n_488), .B2(n_502), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_206), .A2(n_234), .B1(n_495), .B2(n_582), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_208), .A2(n_418), .B1(n_509), .B2(n_615), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_210), .A2(n_420), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_211), .A2(n_254), .B1(n_495), .B2(n_515), .Y(n_1408) );
AO22x2_ASAP7_75t_L g1033 ( .A1(n_212), .A2(n_1034), .B1(n_1053), .B2(n_1054), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_212), .Y(n_1053) );
INVx1_ASAP7_75t_L g997 ( .A(n_213), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_214), .A2(n_278), .B1(n_682), .B2(n_685), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_216), .A2(n_340), .B1(n_625), .B2(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_218), .B(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_221), .A2(n_396), .B1(n_632), .B2(n_709), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_222), .A2(n_227), .B1(n_617), .B2(n_618), .Y(n_616) );
INVxp33_ASAP7_75t_SL g1157 ( .A(n_224), .Y(n_1157) );
AOI21xp33_ASAP7_75t_L g980 ( .A1(n_226), .A2(n_541), .B(n_981), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_229), .A2(n_399), .B1(n_1138), .B2(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_230), .A2(n_259), .B1(n_518), .B2(n_684), .Y(n_806) );
XNOR2x1_ASAP7_75t_L g881 ( .A(n_233), .B(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_235), .A2(n_414), .B1(n_509), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_236), .A2(n_409), .B1(n_919), .B2(n_920), .Y(n_918) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_237), .Y(n_1042) );
XNOR2x1_ASAP7_75t_L g767 ( .A(n_238), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g1377 ( .A(n_240), .Y(n_1377) );
INVx1_ASAP7_75t_L g1082 ( .A(n_241), .Y(n_1082) );
INVx1_ASAP7_75t_L g525 ( .A(n_243), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_244), .A2(n_390), .B1(n_488), .B2(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_245), .A2(n_421), .B1(n_472), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g450 ( .A(n_246), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_247), .A2(n_376), .B1(n_861), .B2(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_249), .B(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_250), .A2(n_416), .B1(n_580), .B2(n_696), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_251), .A2(n_384), .B1(n_688), .B2(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_252), .B(n_600), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_253), .A2(n_353), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_255), .A2(n_312), .B1(n_543), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_258), .A2(n_268), .B1(n_433), .B2(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_260), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_261), .A2(n_264), .B1(n_507), .B2(n_509), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_262), .A2(n_364), .B1(n_782), .B2(n_886), .Y(n_885) );
OR2x2_ASAP7_75t_L g975 ( .A(n_265), .B(n_976), .Y(n_975) );
INVxp67_ASAP7_75t_L g985 ( .A(n_265), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_266), .A2(n_330), .B1(n_576), .B2(n_831), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_270), .A2(n_321), .B1(n_488), .B2(n_801), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_271), .A2(n_294), .B1(n_557), .B2(n_558), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_272), .A2(n_329), .B1(n_554), .B2(n_555), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_273), .A2(n_377), .B1(n_500), .B2(n_705), .Y(n_1368) );
INVx1_ASAP7_75t_L g1383 ( .A(n_275), .Y(n_1383) );
INVx1_ASAP7_75t_L g1374 ( .A(n_276), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_277), .A2(n_392), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_279), .A2(n_280), .B1(n_580), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_281), .A2(n_357), .B1(n_472), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_283), .A2(n_317), .B1(n_600), .B2(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_284), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_285), .A2(n_325), .B1(n_488), .B2(n_502), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_286), .A2(n_358), .B1(n_696), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_287), .A2(n_397), .B1(n_617), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_298), .A2(n_413), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g921 ( .A1(n_299), .A2(n_301), .B1(n_543), .B2(n_922), .C(n_925), .Y(n_921) );
INVx1_ASAP7_75t_L g601 ( .A(n_300), .Y(n_601) );
INVx1_ASAP7_75t_L g760 ( .A(n_302), .Y(n_760) );
AOI22x1_ASAP7_75t_L g610 ( .A1(n_303), .A2(n_611), .B1(n_612), .B2(n_638), .Y(n_610) );
INVx1_ASAP7_75t_L g638 ( .A(n_303), .Y(n_638) );
AO22x1_ASAP7_75t_L g1167 ( .A1(n_303), .A2(n_311), .B1(n_1128), .B2(n_1142), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_304), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_304), .B(n_1123), .Y(n_1122) );
XNOR2x2_ASAP7_75t_L g899 ( .A(n_306), .B(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_308), .A2(n_343), .B1(n_557), .B2(n_558), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_310), .A2(n_415), .B1(n_685), .B2(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g468 ( .A(n_313), .Y(n_468) );
XOR2x2_ASAP7_75t_L g1073 ( .A(n_315), .B(n_1074), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_316), .A2(n_369), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_318), .A2(n_339), .B1(n_576), .B2(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g444 ( .A(n_319), .Y(n_444) );
INVxp67_ASAP7_75t_L g485 ( .A(n_319), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g1036 ( .A1(n_322), .A2(n_541), .B(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g646 ( .A(n_323), .Y(n_646) );
INVx1_ASAP7_75t_L g566 ( .A(n_324), .Y(n_566) );
AOI22xp5_ASAP7_75t_SL g706 ( .A1(n_326), .A2(n_381), .B1(n_707), .B2(n_710), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_328), .A2(n_346), .B1(n_554), .B2(n_555), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g1392 ( .A1(n_331), .A2(n_1393), .B1(n_1394), .B2(n_1410), .Y(n_1392) );
INVx1_ASAP7_75t_L g1410 ( .A(n_331), .Y(n_1410) );
INVx2_ASAP7_75t_L g1109 ( .A(n_332), .Y(n_1109) );
INVxp33_ASAP7_75t_SL g1236 ( .A(n_333), .Y(n_1236) );
INVx1_ASAP7_75t_L g1083 ( .A(n_334), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1396 ( .A1(n_337), .A2(n_1397), .B(n_1398), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_347), .A2(n_400), .B1(n_515), .B2(n_782), .Y(n_1365) );
AO221x2_ASAP7_75t_L g1232 ( .A1(n_348), .A2(n_349), .B1(n_1189), .B2(n_1233), .C(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1097 ( .A(n_350), .Y(n_1097) );
INVx1_ASAP7_75t_L g1086 ( .A(n_354), .Y(n_1086) );
INVx1_ASAP7_75t_L g764 ( .A(n_359), .Y(n_764) );
INVx1_ASAP7_75t_L g1038 ( .A(n_360), .Y(n_1038) );
INVx1_ASAP7_75t_L g470 ( .A(n_363), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_365), .B(n_1020), .Y(n_1019) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_366), .A2(n_775), .B(n_776), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_367), .A2(n_371), .B1(n_617), .B2(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_368), .A2(n_406), .B1(n_696), .B2(n_699), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_370), .A2(n_389), .B1(n_457), .B2(n_771), .Y(n_893) );
INVx1_ASAP7_75t_L g1056 ( .A(n_372), .Y(n_1056) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_373), .A2(n_853), .B(n_875), .Y(n_852) );
INVx1_ASAP7_75t_L g877 ( .A(n_373), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_374), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_378), .B(n_527), .Y(n_1400) );
INVx1_ASAP7_75t_L g812 ( .A(n_379), .Y(n_812) );
XNOR2x2_ASAP7_75t_L g936 ( .A(n_382), .B(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_383), .A2(n_403), .B1(n_576), .B2(n_577), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_385), .A2(n_411), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx1_ASAP7_75t_SL g809 ( .A(n_386), .Y(n_809) );
INVx1_ASAP7_75t_L g568 ( .A(n_392), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_393), .B(n_680), .Y(n_815) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_394), .Y(n_1045) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_402), .A2(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g1399 ( .A(n_407), .Y(n_1399) );
AOI21xp33_ASAP7_75t_L g818 ( .A1(n_410), .A2(n_644), .B(n_819), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_412), .Y(n_946) );
AOI31xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_1102), .A3(n_1105), .B(n_1112), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_790), .B1(n_931), .B2(n_932), .C(n_933), .Y(n_423) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_424), .Y(n_932) );
XNOR2xp5_ASAP7_75t_L g1104 ( .A(n_424), .B(n_790), .Y(n_1104) );
XNOR2x1_ASAP7_75t_L g424 ( .A(n_425), .B(n_669), .Y(n_424) );
AO22x2_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_606), .B1(n_666), .B2(n_668), .Y(n_425) );
INVx1_ASAP7_75t_L g668 ( .A(n_426), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_569), .B1(n_570), .B2(n_605), .Y(n_426) );
INVx1_ASAP7_75t_L g605 ( .A(n_427), .Y(n_605) );
XNOR2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_537), .Y(n_427) );
NAND4xp75_ASAP7_75t_L g429 ( .A(n_430), .B(n_486), .C(n_505), .D(n_517), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g430 ( .A(n_431), .B(n_469), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_455), .B1(n_456), .B2(n_468), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g1382 ( .A1(n_432), .A2(n_1383), .B(n_1384), .Y(n_1382) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g587 ( .A(n_434), .Y(n_587) );
BUFx3_ASAP7_75t_L g709 ( .A(n_434), .Y(n_709) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_447), .Y(n_434) );
AND2x4_ASAP7_75t_L g473 ( .A(n_435), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g508 ( .A(n_435), .B(n_490), .Y(n_508) );
AND2x4_ASAP7_75t_L g547 ( .A(n_435), .B(n_490), .Y(n_547) );
AND2x4_ASAP7_75t_L g654 ( .A(n_435), .B(n_474), .Y(n_654) );
AND2x4_ASAP7_75t_L g657 ( .A(n_435), .B(n_447), .Y(n_657) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_441), .Y(n_435) );
INVx2_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
AND2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g492 ( .A(n_436), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g498 ( .A(n_436), .B(n_494), .Y(n_498) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_438), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g461 ( .A(n_438), .Y(n_461) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp33_ASAP7_75t_L g445 ( .A(n_439), .B(n_446), .Y(n_445) );
NAND2xp33_ASAP7_75t_L g449 ( .A(n_439), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g453 ( .A(n_439), .Y(n_453) );
INVx1_ASAP7_75t_L g465 ( .A(n_439), .Y(n_465) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_440), .B(n_460), .C(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g466 ( .A(n_441), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g494 ( .A(n_442), .Y(n_494) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
AND2x2_ASAP7_75t_L g501 ( .A(n_447), .B(n_492), .Y(n_501) );
AND2x4_ASAP7_75t_L g513 ( .A(n_447), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g523 ( .A(n_447), .B(n_466), .Y(n_523) );
AND2x4_ASAP7_75t_L g554 ( .A(n_447), .B(n_492), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_447), .B(n_497), .Y(n_555) );
AND2x2_ASAP7_75t_L g564 ( .A(n_447), .B(n_466), .Y(n_564) );
AND2x2_ASAP7_75t_L g623 ( .A(n_447), .B(n_492), .Y(n_623) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_454), .Y(n_447) );
INVx1_ASAP7_75t_L g475 ( .A(n_448), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_450), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_452), .A2(n_465), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g474 ( .A(n_454), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g483 ( .A(n_454), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_454), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_456), .A2(n_994), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g874 ( .A(n_457), .Y(n_874) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g590 ( .A(n_458), .Y(n_590) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_458), .Y(n_684) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
AND2x4_ASAP7_75t_L g504 ( .A(n_459), .B(n_492), .Y(n_504) );
AND2x4_ASAP7_75t_L g516 ( .A(n_459), .B(n_497), .Y(n_516) );
AND2x4_ASAP7_75t_L g551 ( .A(n_459), .B(n_497), .Y(n_551) );
AND2x4_ASAP7_75t_L g558 ( .A(n_459), .B(n_492), .Y(n_558) );
AND2x4_ASAP7_75t_L g655 ( .A(n_459), .B(n_466), .Y(n_655) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AND2x2_ASAP7_75t_L g510 ( .A(n_466), .B(n_490), .Y(n_510) );
AND2x4_ASAP7_75t_L g519 ( .A(n_466), .B(n_474), .Y(n_519) );
AND2x4_ASAP7_75t_L g548 ( .A(n_466), .B(n_490), .Y(n_548) );
AND2x2_ASAP7_75t_L g644 ( .A(n_466), .B(n_474), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_476), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_471), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1084) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
BUFx3_ASAP7_75t_L g775 ( .A(n_473), .Y(n_775) );
INVx1_ASAP7_75t_L g949 ( .A(n_473), .Y(n_949) );
AND2x4_ASAP7_75t_L g490 ( .A(n_475), .B(n_491), .Y(n_490) );
BUFx4f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx5_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
BUFx2_ASAP7_75t_L g773 ( .A(n_478), .Y(n_773) );
BUFx2_ASAP7_75t_L g979 ( .A(n_478), .Y(n_979) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
AND2x2_ASAP7_75t_L g658 ( .A(n_479), .B(n_483), .Y(n_658) );
AND2x4_ASAP7_75t_L g755 ( .A(n_479), .B(n_483), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g531 ( .A(n_481), .Y(n_531) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_499), .Y(n_486) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_488), .Y(n_704) );
BUFx6f_ASAP7_75t_L g1026 ( .A(n_488), .Y(n_1026) );
INVx1_ASAP7_75t_L g1091 ( .A(n_488), .Y(n_1091) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_489), .Y(n_582) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_489), .Y(n_625) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
AND2x4_ASAP7_75t_L g496 ( .A(n_490), .B(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g550 ( .A(n_490), .B(n_514), .Y(n_550) );
AND2x4_ASAP7_75t_L g557 ( .A(n_490), .B(n_492), .Y(n_557) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g912 ( .A(n_495), .Y(n_912) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_496), .Y(n_617) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_496), .Y(n_692) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
BUFx3_ASAP7_75t_L g909 ( .A(n_500), .Y(n_909) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx8_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
BUFx2_ASAP7_75t_SL g906 ( .A(n_502), .Y(n_906) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g583 ( .A(n_503), .Y(n_583) );
INVx4_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
INVx4_ASAP7_75t_L g705 ( .A(n_503), .Y(n_705) );
INVx2_ASAP7_75t_L g801 ( .A(n_503), .Y(n_801) );
INVx4_ASAP7_75t_L g831 ( .A(n_503), .Y(n_831) );
INVx1_ASAP7_75t_L g991 ( .A(n_503), .Y(n_991) );
INVx1_ASAP7_75t_L g1079 ( .A(n_503), .Y(n_1079) );
INVx8_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx12f_ASAP7_75t_L g615 ( .A(n_508), .Y(n_615) );
INVx3_ASAP7_75t_L g698 ( .A(n_508), .Y(n_698) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx5_ASAP7_75t_L g580 ( .A(n_510), .Y(n_580) );
INVx1_ASAP7_75t_L g702 ( .A(n_510), .Y(n_702) );
BUFx3_ASAP7_75t_L g861 ( .A(n_510), .Y(n_861) );
BUFx3_ASAP7_75t_L g859 ( .A(n_512), .Y(n_859) );
BUFx12f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g577 ( .A(n_513), .Y(n_577) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_513), .Y(n_650) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_513), .Y(n_694) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_513), .Y(n_782) );
BUFx3_ASAP7_75t_L g913 ( .A(n_515), .Y(n_913) );
BUFx12f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx6_ASAP7_75t_L g619 ( .A(n_516), .Y(n_619) );
INVx2_ASAP7_75t_L g955 ( .A(n_518), .Y(n_955) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx8_ASAP7_75t_SL g562 ( .A(n_519), .Y(n_562) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
INVx2_ASAP7_75t_L g686 ( .A(n_519), .Y(n_686) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_519), .Y(n_771) );
INVx2_ASAP7_75t_L g1380 ( .A(n_519), .Y(n_1380) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g804 ( .A(n_521), .Y(n_804) );
INVx1_ASAP7_75t_L g1397 ( .A(n_521), .Y(n_1397) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g680 ( .A(n_522), .Y(n_680) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
INVx3_ASAP7_75t_L g635 ( .A(n_523), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_528), .B(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_528), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g689 ( .A(n_528), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_528), .B(n_820), .Y(n_819) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_535), .Y(n_530) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_532), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g662 ( .A(n_537), .Y(n_662) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_537), .Y(n_664) );
XOR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_568), .Y(n_537) );
NOR4xp75_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .C(n_552), .D(n_559), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g711 ( .A(n_541), .Y(n_711) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g600 ( .A(n_544), .Y(n_600) );
INVx2_ASAP7_75t_L g632 ( .A(n_544), .Y(n_632) );
INVx2_ASAP7_75t_L g688 ( .A(n_544), .Y(n_688) );
INVx2_ASAP7_75t_L g963 ( .A(n_544), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_553), .B(n_556), .Y(n_552) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_561), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_564), .Y(n_762) );
INVx2_ASAP7_75t_L g840 ( .A(n_564), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_567), .B(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_567), .B(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_567), .B(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_567), .B(n_926), .Y(n_925) );
INVx4_ASAP7_75t_L g964 ( .A(n_567), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_567), .B(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND4xp75_ASAP7_75t_SL g571 ( .A(n_572), .B(n_578), .C(n_584), .D(n_591), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
BUFx3_ASAP7_75t_L g856 ( .A(n_574), .Y(n_856) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
BUFx3_ASAP7_75t_L g903 ( .A(n_580), .Y(n_903) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g631 ( .A(n_587), .Y(n_631) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_587), .Y(n_739) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g920 ( .A(n_590), .Y(n_920) );
INVx3_ASAP7_75t_L g1402 ( .A(n_590), .Y(n_1402) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx3_ASAP7_75t_L g872 ( .A(n_596), .Y(n_872) );
INVx1_ASAP7_75t_L g1021 ( .A(n_596), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_601), .B2(n_602), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_604), .Y(n_765) );
INVx1_ASAP7_75t_L g808 ( .A(n_604), .Y(n_808) );
INVx2_ASAP7_75t_L g868 ( .A(n_604), .Y(n_868) );
BUFx6f_ASAP7_75t_L g1066 ( .A(n_604), .Y(n_1066) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_661), .B(n_663), .Y(n_606) );
AOI22x1_ASAP7_75t_SL g666 ( .A1(n_607), .A2(n_662), .B1(n_664), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g665 ( .A(n_608), .Y(n_665) );
AO22x2_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_639), .B2(n_660), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND4xp75_ASAP7_75t_L g612 ( .A(n_613), .B(n_620), .C(n_627), .D(n_633), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
BUFx3_ASAP7_75t_L g1092 ( .A(n_617), .Y(n_1092) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_618), .Y(n_1077) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g746 ( .A(n_619), .Y(n_746) );
INVx5_ASAP7_75t_L g786 ( .A(n_619), .Y(n_786) );
INVx1_ASAP7_75t_L g857 ( .A(n_619), .Y(n_857) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx4f_ASAP7_75t_L g886 ( .A(n_623), .Y(n_886) );
BUFx2_ASAP7_75t_SL g905 ( .A(n_625), .Y(n_905) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
BUFx3_ASAP7_75t_L g919 ( .A(n_629), .Y(n_919) );
BUFx3_ASAP7_75t_L g952 ( .A(n_631), .Y(n_952) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g642 ( .A(n_635), .Y(n_642) );
INVx2_ASAP7_75t_L g779 ( .A(n_635), .Y(n_779) );
INVx2_ASAP7_75t_L g924 ( .A(n_635), .Y(n_924) );
INVx3_ASAP7_75t_SL g961 ( .A(n_635), .Y(n_961) );
INVx2_ASAP7_75t_L g1061 ( .A(n_635), .Y(n_1061) );
INVx1_ASAP7_75t_L g660 ( .A(n_639), .Y(n_660) );
INVx1_ASAP7_75t_L g714 ( .A(n_639), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_639), .Y(n_715) );
NAND3x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_647), .C(n_651), .Y(n_640) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_642), .Y(n_736) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AND4x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .C(n_656), .D(n_659), .Y(n_651) );
INVx2_ASAP7_75t_L g753 ( .A(n_654), .Y(n_753) );
INVx2_ASAP7_75t_L g759 ( .A(n_655), .Y(n_759) );
INVx1_ASAP7_75t_L g757 ( .A(n_657), .Y(n_757) );
INVx2_ASAP7_75t_L g1046 ( .A(n_657), .Y(n_1046) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_716), .B2(n_788), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AO22x2_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_714), .B2(n_715), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_690), .C(n_706), .Y(n_675) );
INVx1_ASAP7_75t_L g713 ( .A(n_676), .Y(n_713) );
AND3x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .C(n_687), .Y(n_676) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_683), .A2(n_1377), .B1(n_1378), .B2(n_1381), .Y(n_1376) );
INVx4_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx3_ASAP7_75t_L g1016 ( .A(n_684), .Y(n_1016) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND4x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .C(n_695), .D(n_703), .Y(n_690) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_694), .Y(n_910) );
BUFx4f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g799 ( .A(n_698), .Y(n_799) );
INVx1_ASAP7_75t_L g972 ( .A(n_698), .Y(n_972) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_701), .Y(n_724) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g917 ( .A(n_709), .Y(n_917) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g789 ( .A(n_717), .Y(n_789) );
XNOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_740), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
XNOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_728), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .C(n_726), .D(n_727), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_735), .C(n_737), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_734), .Y(n_730) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g870 ( .A(n_739), .Y(n_870) );
INVx2_ASAP7_75t_L g1018 ( .A(n_739), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_739), .Y(n_1087) );
OAI22x1_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_766), .B1(n_767), .B2(n_787), .Y(n_740) );
INVx2_ASAP7_75t_L g787 ( .A(n_741), .Y(n_787) );
NAND4xp75_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .C(n_750), .D(n_761), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_756), .Y(n_750) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B(n_754), .Y(n_751) );
INVx4_ASAP7_75t_L g1043 ( .A(n_755), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_765), .B(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_765), .B(n_982), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_765), .B(n_997), .Y(n_996) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR2x1_ASAP7_75t_L g768 ( .A(n_769), .B(n_780), .Y(n_768) );
NAND4xp25_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .C(n_774), .D(n_778), .Y(n_769) );
INVx2_ASAP7_75t_L g994 ( .A(n_771), .Y(n_994) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_771), .Y(n_1015) );
BUFx2_ASAP7_75t_L g916 ( .A(n_775), .Y(n_916) );
NAND4xp25_ASAP7_75t_SL g780 ( .A(n_781), .B(n_783), .C(n_784), .D(n_785), .Y(n_780) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_786), .Y(n_939) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_790), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_846), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OA22x2_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_810), .B1(n_844), .B2(n_845), .Y(n_792) );
INVx1_ASAP7_75t_SL g844 ( .A(n_793), .Y(n_844) );
XOR2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_809), .Y(n_793) );
NOR2x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_798), .D(n_800), .Y(n_795) );
NAND4xp25_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .C(n_806), .D(n_807), .Y(n_802) );
INVx1_ASAP7_75t_L g1375 ( .A(n_808), .Y(n_1375) );
INVx1_ASAP7_75t_L g845 ( .A(n_810), .Y(n_845) );
XNOR2x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_826), .Y(n_810) );
XNOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
OR2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_821), .Y(n_813) );
NAND4xp25_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .C(n_817), .D(n_818), .Y(n_814) );
NAND4xp25_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .C(n_824), .D(n_825), .Y(n_821) );
BUFx3_ASAP7_75t_L g1004 ( .A(n_826), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_826), .Y(n_1005) );
XNOR2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_843), .Y(n_826) );
NAND4xp75_ASAP7_75t_L g827 ( .A(n_828), .B(n_832), .C(n_835), .D(n_838), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI22x1_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_897), .B1(n_927), .B2(n_929), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g928 ( .A(n_850), .Y(n_928) );
OA22x2_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_879), .B2(n_896), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_863), .Y(n_853) );
INVxp67_ASAP7_75t_L g878 ( .A(n_854), .Y(n_878) );
NAND4xp25_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .C(n_860), .D(n_862), .Y(n_854) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_861), .Y(n_1094) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_863), .B(n_877), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g863 ( .A(n_864), .B(n_869), .C(n_871), .D(n_873), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx3_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g957 ( .A(n_874), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_SL g896 ( .A(n_881), .Y(n_896) );
NOR2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_889), .Y(n_882) );
NAND4xp25_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .C(n_887), .D(n_888), .Y(n_883) );
NAND4xp25_ASAP7_75t_SL g889 ( .A(n_890), .B(n_893), .C(n_894), .D(n_895), .Y(n_889) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
BUFx3_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_SL g930 ( .A(n_899), .Y(n_930) );
NAND4xp75_ASAP7_75t_L g900 ( .A(n_901), .B(n_907), .C(n_914), .D(n_921), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_911), .Y(n_907) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_918), .Y(n_914) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVxp67_ASAP7_75t_SL g1103 ( .A(n_933), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_934), .A2(n_1007), .B1(n_1008), .B2(n_1101), .Y(n_933) );
INVx1_ASAP7_75t_L g1101 ( .A(n_934), .Y(n_1101) );
XNOR2x1_ASAP7_75t_SL g934 ( .A(n_935), .B(n_965), .Y(n_934) );
BUFx3_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND3xp33_ASAP7_75t_SL g937 ( .A(n_938), .B(n_940), .C(n_944), .Y(n_937) );
AND3x1_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .C(n_943), .Y(n_940) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_953), .C(n_958), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_950), .B2(n_951), .Y(n_945) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g1404 ( .A(n_949), .Y(n_1404) );
INVxp67_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_953) );
OAI21xp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_960), .B(n_962), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
AO22x2_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_1004), .B1(n_1005), .B2(n_1006), .Y(n_965) );
INVx2_ASAP7_75t_L g1006 ( .A(n_966), .Y(n_1006) );
XNOR2x1_ASAP7_75t_L g966 ( .A(n_967), .B(n_986), .Y(n_966) );
OAI22x1_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_975), .B1(n_984), .B2(n_985), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_969), .B(n_976), .Y(n_984) );
NAND4xp25_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .C(n_973), .D(n_974), .Y(n_969) );
NAND4xp25_ASAP7_75t_L g976 ( .A(n_977), .B(n_978), .C(n_980), .D(n_983), .Y(n_976) );
NAND4xp75_ASAP7_75t_L g987 ( .A(n_988), .B(n_992), .C(n_998), .D(n_1001), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_989), .B(n_990), .Y(n_988) );
OA21x2_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .B(n_995), .Y(n_992) );
AND2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1000), .Y(n_998) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
AO22x2_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1030), .B2(n_1100), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
XOR2x2_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1029), .Y(n_1011) );
NOR2x1_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1023), .Y(n_1012) );
NAND4xp25_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .C(n_1019), .D(n_1022), .Y(n_1013) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1020), .Y(n_1098) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .C(n_1027), .D(n_1028), .Y(n_1023) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1030), .Y(n_1100) );
AO22x2_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B1(n_1072), .B2(n_1073), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
XOR2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1055), .Y(n_1032) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1034), .Y(n_1054) );
NOR2x1_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1048), .Y(n_1034) );
NAND3xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1039), .C(n_1047), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1043), .B1(n_1044), .B2(n_1046), .Y(n_1040) );
CKINVDCx16_ASAP7_75t_R g1041 ( .A(n_1042), .Y(n_1041) );
OAI21xp33_ASAP7_75t_L g1398 ( .A1(n_1043), .A2(n_1399), .B(n_1400), .Y(n_1398) );
CKINVDCx9p33_ASAP7_75t_R g1044 ( .A(n_1045), .Y(n_1044) );
NAND4xp25_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .C(n_1051), .D(n_1052), .Y(n_1048) );
XNOR2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1057), .Y(n_1055) );
NOR2xp67_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1067), .Y(n_1057) );
NAND4xp25_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .C(n_1062), .D(n_1063), .Y(n_1058) );
NOR2xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1066), .Y(n_1064) );
NAND4xp25_ASAP7_75t_SL g1067 ( .A(n_1068), .B(n_1069), .C(n_1070), .D(n_1071), .Y(n_1067) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
NAND4xp75_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1080), .C(n_1088), .D(n_1095), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1078), .Y(n_1075) );
NOR2x1_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1084), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1093), .Y(n_1088) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
OAI21xp33_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1098), .B(n_1099), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_1106), .Y(n_1105) );
NAND3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1110), .C(n_1111), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1107), .B(n_1388), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1107), .B(n_1389), .Y(n_1412) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
OA21x2_ASAP7_75t_L g1414 ( .A1(n_1108), .A2(n_1129), .B(n_1415), .Y(n_1414) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
AND3x4_ASAP7_75t_L g1128 ( .A(n_1109), .B(n_1122), .C(n_1129), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1109), .B(n_1132), .Y(n_1131) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1110), .B(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1111), .Y(n_1389) );
OAI221xp5_ASAP7_75t_L g1112 ( .A1(n_1113), .A2(n_1356), .B1(n_1358), .B2(n_1385), .C(n_1390), .Y(n_1112) );
O2A1O1Ixp33_ASAP7_75t_SL g1113 ( .A1(n_1114), .A2(n_1237), .B(n_1261), .C(n_1327), .Y(n_1113) );
NAND5xp2_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1203), .C(n_1218), .D(n_1227), .E(n_1232), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1163), .B1(n_1168), .B2(n_1176), .C(n_1179), .Y(n_1115) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_1117), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1133), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1118), .B(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1118), .B(n_1281), .Y(n_1319) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1119), .B(n_1146), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1119), .B(n_1165), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_1119), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1119), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1119), .B(n_1207), .Y(n_1231) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_1119), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1119), .B(n_1146), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1119), .B(n_1253), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1119), .B(n_1165), .Y(n_1299) );
AND2x4_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1127), .Y(n_1119) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1124), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_1122), .B(n_1131), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1122), .B(n_1124), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1191 ( .A(n_1122), .B(n_1124), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1124), .B(n_1126), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1124), .B(n_1126), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1124), .B(n_1126), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1126), .B(n_1131), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1126), .B(n_1131), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_1126), .B(n_1131), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g1415 ( .A(n_1126), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1144), .Y(n_1133) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1134), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1134), .B(n_1173), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1134), .B(n_1170), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1134), .B(n_1158), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1139), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_1135), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1135), .B(n_1139), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1138), .Y(n_1151) );
BUFx2_ASAP7_75t_L g1357 ( .A(n_1138), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1139), .B(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1139), .B(n_1175), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1139), .B(n_1170), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1139), .B(n_1229), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1139), .B(n_1159), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1143), .Y(n_1139) );
INVx3_ASAP7_75t_L g1154 ( .A(n_1141), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1144), .B(n_1195), .Y(n_1202) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1145), .B(n_1174), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1158), .Y(n_1145) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1146), .Y(n_1173) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1146), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1146), .B(n_1212), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1146), .B(n_1174), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1146), .B(n_1299), .Y(n_1298) );
HB1xp67_ASAP7_75t_L g1303 ( .A(n_1146), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1146), .B(n_1165), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1153), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1150), .B1(n_1151), .B2(n_1152), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_1148), .A2(n_1151), .B1(n_1235), .B2(n_1236), .Y(n_1234) );
INVx3_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
XOR2x1_ASAP7_75t_L g1362 ( .A(n_1152), .B(n_1363), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1155), .B1(n_1156), .B2(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1154), .Y(n_1233) );
OAI311xp33_ASAP7_75t_L g1179 ( .A1(n_1158), .A2(n_1180), .A3(n_1184), .B1(n_1193), .C1(n_1199), .Y(n_1179) );
A2O1A1Ixp33_ASAP7_75t_L g1193 ( .A1(n_1158), .A2(n_1194), .B(n_1195), .C(n_1196), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1158), .B(n_1175), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1158), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1158), .B(n_1183), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1158), .B(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1158), .B(n_1257), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1158), .B(n_1175), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1158), .B(n_1226), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1158), .B(n_1174), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1158), .B(n_1283), .Y(n_1336) );
INVx3_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1159), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1159), .B(n_1207), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1162), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1163), .B(n_1198), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1163), .B(n_1186), .Y(n_1254) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
CKINVDCx6p67_ASAP7_75t_R g1178 ( .A(n_1165), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1165), .B(n_1213), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1165), .B(n_1186), .Y(n_1253) );
OR2x6_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1172), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1170), .B(n_1195), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1170), .B(n_1175), .Y(n_1276) );
AOI211xp5_ASAP7_75t_L g1332 ( .A1(n_1170), .A2(n_1173), .B(n_1174), .C(n_1333), .Y(n_1332) );
AND3x1_ASAP7_75t_L g1349 ( .A(n_1170), .B(n_1224), .C(n_1226), .Y(n_1349) );
INVx3_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1173), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1173), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1173), .B(n_1305), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1173), .B(n_1287), .Y(n_1345) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1174), .Y(n_1257) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_1176), .A2(n_1319), .B(n_1320), .Y(n_1318) );
CKINVDCx14_ASAP7_75t_R g1176 ( .A(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
NAND3xp33_ASAP7_75t_L g1227 ( .A(n_1178), .B(n_1228), .C(n_1230), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1178), .B(n_1186), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1178), .B(n_1245), .Y(n_1310) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1183), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1183), .B(n_1207), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1351 ( .A(n_1183), .B(n_1303), .Y(n_1351) );
INVx3_ASAP7_75t_L g1194 ( .A(n_1185), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1185), .B(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1185), .B(n_1221), .Y(n_1220) );
INVx5_ASAP7_75t_L g1274 ( .A(n_1185), .Y(n_1274) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_1185), .A2(n_1326), .B1(n_1338), .B2(n_1341), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1185), .B(n_1299), .Y(n_1342) );
INVx3_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1186), .B(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1186), .B(n_1245), .Y(n_1244) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1187), .B(n_1315), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1187), .B(n_1201), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1192), .Y(n_1187) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx2_ASAP7_75t_SL g1190 ( .A(n_1191), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1194), .B(n_1212), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1195), .B(n_1207), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1195), .B(n_1206), .Y(n_1284) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1195), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1195), .B(n_1229), .Y(n_1355) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI21xp33_ASAP7_75t_L g1338 ( .A1(n_1197), .A2(n_1296), .B(n_1339), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1202), .Y(n_1199) );
AOI222xp33_ASAP7_75t_L g1279 ( .A1(n_1200), .A2(n_1219), .B1(n_1251), .B2(n_1280), .C1(n_1281), .C2(n_1284), .Y(n_1279) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1202), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1210), .B1(n_1214), .B2(n_1216), .Y(n_1203) );
INVxp33_ASAP7_75t_SL g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_SL g1206 ( .A(n_1207), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1207), .B(n_1250), .Y(n_1326) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
OAI32xp33_ASAP7_75t_L g1352 ( .A1(n_1211), .A2(n_1231), .A3(n_1253), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1213), .Y(n_1225) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
AOI222xp33_ASAP7_75t_L g1328 ( .A1(n_1216), .A2(n_1310), .B1(n_1329), .B2(n_1330), .C1(n_1332), .C2(n_1335), .Y(n_1328) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1222), .B1(n_1223), .B2(n_1226), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1221), .B(n_1267), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1223), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
A2O1A1Ixp33_ASAP7_75t_L g1317 ( .A1(n_1228), .A2(n_1277), .B(n_1318), .C(n_1322), .Y(n_1317) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1228), .Y(n_1353) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1232), .Y(n_1293) );
A2O1A1Ixp33_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1239), .B(n_1243), .C(n_1246), .Y(n_1237) );
AOI21xp33_ASAP7_75t_L g1346 ( .A1(n_1238), .A2(n_1290), .B(n_1319), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
O2A1O1Ixp33_ASAP7_75t_L g1350 ( .A1(n_1241), .A2(n_1280), .B(n_1351), .C(n_1352), .Y(n_1350) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
AOI221xp5_ASAP7_75t_SL g1246 ( .A1(n_1247), .A2(n_1252), .B1(n_1254), .B2(n_1255), .C(n_1258), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1249), .Y(n_1247) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1248), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1249), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
NAND3xp33_ASAP7_75t_L g1272 ( .A(n_1250), .B(n_1273), .C(n_1274), .Y(n_1272) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1252), .A2(n_1295), .B1(n_1297), .B2(n_1300), .C(n_1306), .Y(n_1294) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1254), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1255), .B(n_1276), .Y(n_1301) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1257), .B(n_1268), .Y(n_1267) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1260), .Y(n_1270) );
NAND5xp2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1294), .C(n_1308), .D(n_1317), .E(n_1323), .Y(n_1261) );
AOI211xp5_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1264), .B(n_1271), .C(n_1285), .Y(n_1262) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_1263), .A2(n_1286), .B1(n_1288), .B2(n_1291), .C(n_1293), .Y(n_1285) );
INVxp67_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1270), .Y(n_1266) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1275), .C(n_1279), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_1273), .B(n_1289), .Y(n_1288) );
CKINVDCx14_ASAP7_75t_R g1322 ( .A(n_1274), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1274), .B(n_1325), .Y(n_1324) );
A2O1A1Ixp33_ASAP7_75t_L g1347 ( .A1(n_1274), .A2(n_1276), .B(n_1348), .C(n_1349), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .Y(n_1275) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1278), .B(n_1307), .Y(n_1306) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
O2A1O1Ixp33_ASAP7_75t_L g1343 ( .A1(n_1292), .A2(n_1313), .B(n_1344), .C(n_1346), .Y(n_1343) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx2_ASAP7_75t_L g1315 ( .A(n_1299), .Y(n_1315) );
OAI21xp33_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B(n_1304), .Y(n_1300) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1304), .Y(n_1329) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1310), .B1(n_1311), .B2(n_1313), .C(n_1316), .Y(n_1308) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1315), .Y(n_1340) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1321), .B(n_1340), .Y(n_1339) );
INVxp67_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
NAND5xp2_ASAP7_75t_SL g1327 ( .A(n_1328), .B(n_1337), .C(n_1343), .D(n_1347), .E(n_1350), .Y(n_1327) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1369), .Y(n_1363) );
AND4x1_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .C(n_1367), .D(n_1368), .Y(n_1364) );
NOR3xp33_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1376), .C(n_1382), .Y(n_1369) );
NAND2xp5_ASAP7_75t_SL g1370 ( .A(n_1371), .B(n_1372), .Y(n_1370) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .Y(n_1373) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
HB1xp67_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVxp33_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVxp67_ASAP7_75t_SL g1393 ( .A(n_1394), .Y(n_1393) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1405), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g1395 ( .A(n_1396), .B(n_1401), .C(n_1403), .Y(n_1395) );
NAND4xp25_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1407), .C(n_1408), .D(n_1409), .Y(n_1405) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
endmodule