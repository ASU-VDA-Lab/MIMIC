module fake_ibex_1457_n_1465 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1465);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1465;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1296;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1115;
wire n_998;
wire n_1395;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1361;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1369;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_183),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_29),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_131),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_123),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_75),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_201),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_122),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_89),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_66),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_18),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_132),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_76),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_164),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_86),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_160),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_249),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_188),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_171),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_45),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_103),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_210),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_48),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_192),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_111),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_112),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_94),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_102),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_245),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_182),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_168),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_107),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_173),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_77),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_99),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_17),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_191),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_57),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_180),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_133),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_5),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_118),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_256),
.B(n_228),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_159),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_7),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_71),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_200),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_155),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_44),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_78),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_68),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_152),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_232),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_218),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_75),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_61),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_127),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_154),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_63),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_69),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_167),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_84),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_52),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_195),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_172),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_80),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_46),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_213),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_80),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_33),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_10),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_4),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_96),
.Y(n_362)
);

BUFx2_ASAP7_75t_SL g363 ( 
.A(n_189),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_148),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_28),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_143),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_52),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_140),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_204),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_138),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_174),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_216),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_244),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_31),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_186),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_4),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_26),
.B(n_227),
.Y(n_377)
);

BUFx8_ASAP7_75t_SL g378 ( 
.A(n_120),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_24),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_42),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_214),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_27),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_124),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_11),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_149),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_261),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_56),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_25),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_44),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_234),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_229),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_22),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_53),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_219),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_255),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_60),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_177),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_R g398 ( 
.A(n_13),
.B(n_110),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_250),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_231),
.B(n_94),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_176),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_207),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_9),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_130),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_49),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_43),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_63),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_223),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_85),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_144),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_211),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_187),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_254),
.B(n_116),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_34),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_247),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_93),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_32),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_98),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_209),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_78),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_97),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_169),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_14),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_197),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_241),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_158),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_81),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_221),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_156),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_196),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_157),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_23),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_1),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_134),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_70),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_19),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_185),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_243),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_257),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_45),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_32),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_161),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_181),
.B(n_129),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_208),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_65),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_114),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_34),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_193),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_286),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_286),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_323),
.B(n_324),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_289),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_328),
.B(n_0),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_275),
.A2(n_117),
.B(n_115),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_289),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_347),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_289),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_318),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_291),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_378),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_291),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_3),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_302),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_318),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_283),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_291),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_332),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_330),
.B(n_262),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_320),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g471 ( 
.A(n_264),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_328),
.B(n_6),
.Y(n_473)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_275),
.A2(n_121),
.B(n_119),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_332),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_416),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_291),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_289),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_320),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_302),
.B(n_345),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_344),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_289),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_289),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_320),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_8),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_287),
.A2(n_126),
.B(n_125),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_269),
.B(n_11),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_436),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_287),
.A2(n_135),
.B(n_128),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_415),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_289),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_353),
.B(n_12),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_436),
.B(n_12),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_344),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_263),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_301),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_380),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_380),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_283),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_300),
.A2(n_372),
.B(n_352),
.Y(n_508)
);

BUFx8_ASAP7_75t_SL g509 ( 
.A(n_388),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_301),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_441),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_300),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_413),
.B(n_136),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_301),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_264),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_15),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_278),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_406),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_316),
.B(n_16),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_301),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_266),
.B(n_18),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_378),
.Y(n_523)
);

CKINVDCx6p67_ASAP7_75t_R g524 ( 
.A(n_313),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_402),
.B(n_20),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_352),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_372),
.A2(n_139),
.B(n_137),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_265),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_301),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_348),
.B(n_20),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_267),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_375),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_375),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_381),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_381),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_399),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_388),
.A2(n_421),
.B1(n_398),
.B2(n_280),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_276),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_399),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_401),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_273),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_301),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_401),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_274),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_285),
.Y(n_545)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_460),
.Y(n_546)
);

INVx8_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_451),
.B(n_327),
.Y(n_548)
);

BUFx6f_ASAP7_75t_SL g549 ( 
.A(n_496),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_506),
.B(n_404),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_524),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_517),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_480),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_296),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_506),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_496),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_469),
.A2(n_284),
.B1(n_299),
.B2(n_288),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_496),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_513),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_499),
.B(n_465),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_511),
.B(n_280),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_462),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_456),
.A2(n_359),
.B1(n_433),
.B2(n_290),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_469),
.A2(n_308),
.B1(n_310),
.B2(n_306),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_453),
.B(n_392),
.C(n_359),
.Y(n_575)
);

OA22x2_ASAP7_75t_L g576 ( 
.A1(n_456),
.A2(n_433),
.B1(n_440),
.B2(n_290),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_524),
.A2(n_440),
.B1(n_445),
.B2(n_421),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_469),
.A2(n_322),
.B1(n_326),
.B2(n_319),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_499),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_454),
.A2(n_307),
.B(n_303),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_468),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_472),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_472),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_514),
.A2(n_343),
.B1(n_357),
.B2(n_338),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_533),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_531),
.B(n_311),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_537),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

XNOR2x2_ASAP7_75t_SL g595 ( 
.A(n_509),
.B(n_361),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_476),
.B(n_445),
.C(n_271),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_541),
.B(n_315),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_490),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_268),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_512),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

BUFx4f_ASAP7_75t_L g606 ( 
.A(n_514),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_480),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_532),
.B(n_317),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_504),
.B(n_272),
.Y(n_612)
);

AND3x2_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_394),
.C(n_365),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_485),
.B(n_325),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_463),
.B(n_268),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_329),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_528),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_463),
.B(n_277),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_532),
.B(n_335),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_543),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_535),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_463),
.B(n_277),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_543),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_535),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_532),
.B(n_339),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_523),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_471),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_538),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_504),
.B(n_340),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_532),
.B(n_341),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_514),
.A2(n_298),
.B1(n_364),
.B2(n_314),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_452),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_544),
.B(n_279),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

AND3x2_ASAP7_75t_L g640 ( 
.A(n_486),
.B(n_367),
.C(n_362),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_532),
.B(n_534),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_544),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_489),
.A2(n_298),
.B1(n_364),
.B2(n_314),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_489),
.B(n_346),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_536),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_536),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_544),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_545),
.B(n_349),
.Y(n_648)
);

INVx6_ASAP7_75t_L g649 ( 
.A(n_452),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_537),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_536),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_545),
.B(n_279),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_478),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_459),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_449),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_465),
.B(n_292),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_536),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_450),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_539),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_525),
.B(n_281),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_450),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_458),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_539),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_534),
.B(n_356),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_452),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_508),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_539),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_520),
.B(n_379),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_458),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_530),
.B(n_297),
.C(n_270),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_540),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_464),
.B(n_360),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_459),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_540),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_540),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_534),
.B(n_366),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_464),
.B(n_282),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_540),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_508),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_508),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_540),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_459),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_478),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_478),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_534),
.B(n_368),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_466),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_534),
.B(n_370),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_515),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_542),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_542),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_617),
.B(n_522),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_568),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_642),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_556),
.B(n_542),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_606),
.A2(n_457),
.B1(n_483),
.B2(n_455),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_606),
.A2(n_559),
.B1(n_550),
.B2(n_555),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_571),
.Y(n_701)
);

INVx8_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_655),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_569),
.B(n_467),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_570),
.A2(n_475),
.B(n_481),
.C(n_467),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_551),
.B(n_475),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_548),
.B(n_293),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_659),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_553),
.A2(n_483),
.B1(n_484),
.B2(n_457),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_547),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_561),
.A2(n_434),
.B1(n_446),
.B2(n_425),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_591),
.B(n_448),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_662),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_428),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_584),
.B(n_429),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_671),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_560),
.A2(n_493),
.B1(n_521),
.B2(n_500),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_563),
.A2(n_493),
.B1(n_521),
.B2(n_500),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_638),
.B(n_652),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_603),
.B(n_304),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_562),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_448),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_549),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_557),
.B(n_431),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_557),
.B(n_437),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_679),
.B(n_437),
.Y(n_729)
);

O2A1O1Ixp5_ASAP7_75t_L g730 ( 
.A1(n_681),
.A2(n_373),
.B(n_386),
.C(n_385),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_309),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_670),
.B(n_481),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_498),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_644),
.B(n_294),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_561),
.B(n_503),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_672),
.B(n_566),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_661),
.B(n_614),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_567),
.A2(n_529),
.B(n_488),
.C(n_491),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_608),
.B(n_295),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_614),
.B(n_601),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_625),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_589),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_585),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_615),
.B(n_501),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_620),
.B(n_502),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_619),
.B(n_312),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_624),
.B(n_505),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_596),
.A2(n_519),
.B(n_507),
.C(n_387),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_656),
.A2(n_565),
.B1(n_636),
.B2(n_576),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_586),
.Y(n_751)
);

INVx8_ASAP7_75t_L g752 ( 
.A(n_580),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_632),
.B(n_390),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_656),
.A2(n_396),
.B1(n_407),
.B2(n_382),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_579),
.A2(n_529),
.B1(n_417),
.B2(n_420),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_588),
.B(n_336),
.C(n_333),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_631),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_633),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_616),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_616),
.B(n_395),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_587),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_588),
.B(n_305),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_580),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_554),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_643),
.B(n_337),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_592),
.B(n_397),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_648),
.A2(n_488),
.B(n_491),
.C(n_454),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_611),
.B(n_321),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_598),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_599),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_667),
.A2(n_527),
.B(n_474),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_682),
.A2(n_427),
.B1(n_432),
.B2(n_409),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_565),
.B(n_503),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_682),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_637),
.B(n_331),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_605),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_597),
.B(n_410),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_609),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_674),
.B(n_422),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_576),
.A2(n_447),
.B1(n_497),
.B2(n_474),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_630),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_653),
.B(n_424),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_613),
.A2(n_351),
.B1(n_354),
.B2(n_350),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_653),
.B(n_426),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_640),
.A2(n_358),
.B1(n_374),
.B2(n_355),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_565),
.B(n_363),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_637),
.B(n_474),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_648),
.A2(n_439),
.B(n_442),
.C(n_430),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_689),
.B(n_334),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_641),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_577),
.B(n_342),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_641),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_685),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_618),
.A2(n_444),
.B(n_443),
.C(n_400),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_650),
.B(n_376),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_582),
.A2(n_497),
.B1(n_527),
.B2(n_474),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_685),
.B(n_497),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_564),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_546),
.B(n_377),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_564),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_686),
.A2(n_527),
.B(n_518),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_369),
.Y(n_804)
);

BUFx8_ASAP7_75t_L g805 ( 
.A(n_595),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_552),
.B(n_371),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_610),
.B(n_383),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_634),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_691),
.B(n_391),
.Y(n_809)
);

BUFx5_ASAP7_75t_L g810 ( 
.A(n_552),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_692),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_693),
.A2(n_628),
.B(n_635),
.C(n_621),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_635),
.A2(n_678),
.B1(n_687),
.B2(n_665),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_666),
.B(n_408),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_612),
.B(n_278),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_665),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_678),
.B(n_411),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_690),
.B(n_412),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_690),
.B(n_419),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_581),
.B(n_403),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_583),
.B(n_414),
.C(n_405),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_590),
.B(n_418),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_SL g823 ( 
.A(n_593),
.B(n_393),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_811),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_702),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_732),
.B(n_21),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_781),
.B(n_461),
.C(n_594),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_740),
.A2(n_604),
.B(n_607),
.C(n_600),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_703),
.Y(n_829)
);

OA21x2_ASAP7_75t_L g830 ( 
.A1(n_767),
.A2(n_738),
.B(n_771),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_772),
.A2(n_600),
.B1(n_607),
.B2(n_604),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_702),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_702),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_740),
.A2(n_626),
.B(n_627),
.C(n_623),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_752),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_775),
.A2(n_626),
.B(n_623),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_749),
.A2(n_629),
.B(n_639),
.C(n_627),
.Y(n_837)
);

AO22x1_ASAP7_75t_L g838 ( 
.A1(n_805),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_760),
.A2(n_639),
.B(n_629),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_710),
.B(n_24),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_772),
.A2(n_755),
.B1(n_711),
.B2(n_700),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_749),
.A2(n_645),
.B(n_646),
.C(n_651),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_781),
.B(n_461),
.C(n_651),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_731),
.B(n_30),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_752),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_732),
.B(n_30),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_737),
.B(n_31),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_730),
.A2(n_669),
.B(n_657),
.C(n_683),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_803),
.A2(n_660),
.B(n_658),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_704),
.B(n_33),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_704),
.B(n_35),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_752),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_706),
.A2(n_664),
.B(n_660),
.C(n_683),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_763),
.B(n_37),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_722),
.A2(n_669),
.B(n_668),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_746),
.B(n_38),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_706),
.B(n_39),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_744),
.A2(n_676),
.B(n_673),
.C(n_680),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_697),
.A2(n_676),
.B(n_673),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_723),
.B(n_39),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_757),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_SL g862 ( 
.A(n_823),
.B(n_748),
.C(n_782),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_707),
.B(n_40),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_787),
.B(n_694),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_726),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_753),
.B(n_41),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_753),
.B(n_41),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_697),
.A2(n_680),
.B(n_677),
.Y(n_868)
);

OAI321xp33_ASAP7_75t_L g869 ( 
.A1(n_780),
.A2(n_494),
.A3(n_477),
.B1(n_482),
.B2(n_487),
.C(n_492),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_759),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_789),
.A2(n_654),
.B(n_574),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_789),
.A2(n_654),
.B(n_574),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_733),
.B(n_47),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_708),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_705),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_765),
.B(n_50),
.Y(n_876)
);

NOR2x1p5_ASAP7_75t_L g877 ( 
.A(n_725),
.B(n_53),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_736),
.B(n_54),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_795),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_780),
.B(n_55),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_713),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_716),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_717),
.A2(n_494),
.B1(n_482),
.B2(n_487),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_745),
.A2(n_747),
.B(n_798),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_726),
.B(n_477),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_743),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_788),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_727),
.B(n_55),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_754),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_728),
.B(n_58),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_701),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_761),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_724),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_SL g894 ( 
.A1(n_774),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_764),
.Y(n_895)
);

OR2x6_ASAP7_75t_SL g896 ( 
.A(n_797),
.B(n_62),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_715),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_729),
.A2(n_684),
.B(n_675),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_756),
.A2(n_492),
.B1(n_688),
.B2(n_684),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_770),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_754),
.B(n_67),
.C(n_68),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_808),
.A2(n_688),
.B(n_684),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_773),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_699),
.A2(n_175),
.B(n_259),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_696),
.A2(n_698),
.B1(n_790),
.B2(n_758),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_788),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_750),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_815),
.B(n_72),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_766),
.B(n_73),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_709),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_766),
.B(n_79),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_751),
.Y(n_913)
);

AO32x1_ASAP7_75t_L g914 ( 
.A1(n_816),
.A2(n_79),
.A3(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_788),
.Y(n_915)
);

NOR2x1_ASAP7_75t_L g916 ( 
.A(n_801),
.B(n_82),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_725),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_778),
.B(n_86),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_L g919 ( 
.A1(n_762),
.A2(n_88),
.B(n_89),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_L g920 ( 
.A(n_793),
.B(n_88),
.C(n_90),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_709),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_921)
);

INVx6_ASAP7_75t_L g922 ( 
.A(n_801),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_784),
.B(n_92),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_774),
.B(n_801),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_812),
.A2(n_190),
.B(n_242),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_786),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_774),
.B(n_95),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_695),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_769),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_821),
.B(n_100),
.C(n_101),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_792),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_796),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_794),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_734),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_718),
.B(n_108),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_718),
.B(n_108),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_699),
.A2(n_198),
.B(n_239),
.Y(n_938)
);

OA22x2_ASAP7_75t_L g939 ( 
.A1(n_742),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_939)
);

BUFx12f_ASAP7_75t_L g940 ( 
.A(n_768),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_721),
.B(n_113),
.Y(n_941)
);

OA22x2_ASAP7_75t_L g942 ( 
.A1(n_783),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_719),
.B(n_151),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_791),
.B(n_153),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_783),
.A2(n_162),
.B(n_163),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_785),
.A2(n_165),
.B1(n_166),
.B2(n_179),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_809),
.B(n_194),
.C(n_199),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_741),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_720),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_810),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_807),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_804),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_819),
.B(n_212),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_820),
.A2(n_222),
.B1(n_224),
.B2(n_226),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_819),
.A2(n_776),
.B1(n_739),
.B2(n_818),
.Y(n_955)
);

NAND2xp33_ASAP7_75t_L g956 ( 
.A(n_810),
.B(n_230),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_804),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_814),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_817),
.B(n_813),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_822),
.B(n_810),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_825),
.B(n_806),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_861),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_825),
.B(n_799),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_864),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_861),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_891),
.Y(n_966)
);

AO32x2_ASAP7_75t_L g967 ( 
.A1(n_911),
.A2(n_233),
.A3(n_237),
.B1(n_800),
.B2(n_802),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_835),
.B(n_832),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_835),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_897),
.A2(n_872),
.B(n_871),
.Y(n_970)
);

AO21x1_ASAP7_75t_L g971 ( 
.A1(n_905),
.A2(n_938),
.B(n_954),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_874),
.B(n_881),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_841),
.A2(n_867),
.B(n_866),
.C(n_880),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_959),
.A2(n_834),
.B(n_828),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_882),
.B(n_876),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_858),
.A2(n_853),
.B(n_843),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_855),
.A2(n_836),
.B(n_898),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_832),
.B(n_845),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_849),
.A2(n_902),
.B(n_960),
.Y(n_979)
);

NOR2x1_ASAP7_75t_R g980 ( 
.A(n_915),
.B(n_852),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_840),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_892),
.B(n_900),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_827),
.A2(n_830),
.B(n_906),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_908),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_903),
.B(n_904),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_870),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_830),
.A2(n_848),
.B(n_878),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_R g988 ( 
.A(n_907),
.B(n_924),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_925),
.A2(n_847),
.B(n_873),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_SL g990 ( 
.A(n_943),
.B(n_887),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_895),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_833),
.B(n_958),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_833),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_840),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_887),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_877),
.B(n_924),
.Y(n_996)
);

INVx4_ASAP7_75t_SL g997 ( 
.A(n_943),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_L g998 ( 
.A(n_930),
.B(n_920),
.C(n_935),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_887),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_865),
.B(n_844),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_856),
.B(n_860),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_936),
.A2(n_941),
.B(n_937),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_940),
.B(n_862),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_957),
.B(n_952),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_826),
.A2(n_846),
.B1(n_851),
.B2(n_850),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_857),
.A2(n_912),
.B(n_918),
.C(n_910),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_SL g1007 ( 
.A1(n_945),
.A2(n_921),
.B(n_889),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_924),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_913),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_854),
.B(n_879),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_839),
.A2(n_868),
.B(n_859),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_896),
.B(n_927),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_956),
.A2(n_945),
.B(n_921),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_922),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_854),
.Y(n_1015)
);

AO32x2_ASAP7_75t_L g1016 ( 
.A1(n_894),
.A2(n_883),
.A3(n_831),
.B1(n_914),
.B2(n_919),
.Y(n_1016)
);

INVx3_ASAP7_75t_SL g1017 ( 
.A(n_922),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_923),
.B(n_929),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_933),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_824),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_824),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_SL g1022 ( 
.A(n_901),
.B(n_917),
.C(n_932),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_870),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_948),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_831),
.A2(n_890),
.B(n_888),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_838),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_893),
.B(n_931),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_926),
.B(n_948),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_886),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_950),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_928),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_939),
.Y(n_1032)
);

AOI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_909),
.A2(n_939),
.B(n_899),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_SL g1034 ( 
.A1(n_955),
.A2(n_946),
.B(n_949),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_934),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_947),
.B(n_885),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_914),
.A2(n_606),
.B1(n_572),
.B2(n_579),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_864),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_864),
.B(n_732),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_861),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_864),
.B(n_732),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_841),
.A2(n_606),
.B1(n_572),
.B2(n_579),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_731),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1044)
);

NOR4xp25_ASAP7_75t_L g1045 ( 
.A(n_837),
.B(n_842),
.C(n_875),
.D(n_889),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_864),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_861),
.B(n_731),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_861),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_825),
.B(n_835),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_837),
.A2(n_842),
.B(n_740),
.C(n_863),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_864),
.B(n_829),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_861),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_825),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_832),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_837),
.A2(n_842),
.B(n_740),
.C(n_863),
.Y(n_1058)
);

NAND2x1p5_ASAP7_75t_L g1059 ( 
.A(n_825),
.B(n_835),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_864),
.B(n_732),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_837),
.A2(n_842),
.B(n_740),
.C(n_863),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_864),
.B(n_732),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_825),
.B(n_835),
.Y(n_1064)
);

NOR4xp25_ASAP7_75t_L g1065 ( 
.A(n_837),
.B(n_842),
.C(n_875),
.D(n_889),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_864),
.B(n_732),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_837),
.A2(n_842),
.B(n_740),
.C(n_863),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_861),
.A2(n_711),
.B1(n_735),
.B2(n_712),
.Y(n_1068)
);

AOI31xp67_ASAP7_75t_L g1069 ( 
.A1(n_942),
.A2(n_944),
.A3(n_951),
.B(n_953),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_864),
.B(n_732),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_841),
.A2(n_606),
.B1(n_572),
.B2(n_579),
.Y(n_1072)
);

CKINVDCx11_ASAP7_75t_R g1073 ( 
.A(n_861),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_864),
.B(n_732),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_864),
.B(n_732),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_SL g1078 ( 
.A(n_825),
.B(n_835),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_861),
.B(n_731),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_837),
.A2(n_842),
.B(n_740),
.C(n_863),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_861),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_861),
.B(n_643),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_864),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_SL g1086 ( 
.A(n_825),
.B(n_835),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_SL g1087 ( 
.A(n_861),
.B(n_631),
.C(n_757),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_861),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1089)
);

BUFx8_ASAP7_75t_L g1090 ( 
.A(n_915),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_861),
.B(n_643),
.Y(n_1091)
);

INVx3_ASAP7_75t_SL g1092 ( 
.A(n_825),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_864),
.Y(n_1093)
);

NOR4xp25_ASAP7_75t_L g1094 ( 
.A(n_837),
.B(n_842),
.C(n_875),
.D(n_889),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_861),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_864),
.B(n_732),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_864),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_864),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_864),
.B(n_732),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_825),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_861),
.B(n_712),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_852),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_825),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_864),
.B(n_732),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_861),
.B(n_731),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_861),
.B(n_712),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_884),
.A2(n_738),
.B(n_767),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_825),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_864),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_864),
.A2(n_775),
.B(n_771),
.Y(n_1113)
);

AND3x4_ASAP7_75t_L g1114 ( 
.A(n_916),
.B(n_596),
.C(n_595),
.Y(n_1114)
);

AOI211x1_ASAP7_75t_L g1115 ( 
.A1(n_864),
.A2(n_749),
.B(n_897),
.C(n_911),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_864),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_971),
.A2(n_1013),
.A3(n_1006),
.B(n_1005),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_964),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1005),
.A2(n_1058),
.A3(n_1062),
.B(n_1052),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1067),
.A2(n_1081),
.A3(n_970),
.B(n_979),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1044),
.A2(n_1054),
.B(n_1048),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_962),
.A2(n_1088),
.B1(n_1060),
.B2(n_1066),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_1084),
.B(n_1076),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1038),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1083),
.B(n_1091),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_977),
.A2(n_1032),
.A3(n_1037),
.B(n_1089),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1046),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1049),
.A2(n_1077),
.B(n_1070),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1056),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1099),
.A2(n_1113),
.B(n_1112),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1070),
.A2(n_1079),
.B(n_1077),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1085),
.B(n_1093),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1097),
.B(n_1098),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_981),
.A2(n_973),
.B(n_997),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1090),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1059),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_1072),
.B1(n_1022),
.B2(n_1012),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1111),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1116),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1092),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1053),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1078),
.B(n_1051),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1059),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1105),
.A2(n_1109),
.B(n_1011),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1040),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_974),
.B(n_1002),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_987),
.A2(n_983),
.B(n_974),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_1037),
.B(n_1042),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1151)
);

INVxp33_ASAP7_75t_L g1152 ( 
.A(n_1050),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_989),
.A2(n_976),
.B(n_1025),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1053),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1101),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1096),
.B(n_1100),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1106),
.B(n_1043),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1115),
.B(n_985),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_984),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1072),
.A2(n_1015),
.B1(n_994),
.B2(n_985),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_1007),
.A2(n_997),
.B(n_990),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1104),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1082),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_965),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_966),
.B(n_972),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1047),
.B(n_1080),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1090),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1064),
.B(n_997),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1086),
.B(n_995),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_995),
.B(n_969),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1055),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1004),
.B(n_1095),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_1033),
.A2(n_1034),
.B(n_1010),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_1087),
.B(n_1008),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1068),
.B(n_1107),
.Y(n_1175)
);

BUFx5_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1009),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_998),
.A2(n_1065),
.B(n_1094),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1045),
.A2(n_1065),
.B(n_1094),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_994),
.A2(n_1015),
.B(n_996),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_991),
.B(n_1110),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1045),
.B(n_998),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1028),
.B(n_1057),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1001),
.A2(n_1018),
.B(n_975),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1103),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_993),
.B(n_982),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_992),
.B(n_1003),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1036),
.A2(n_1108),
.B(n_1102),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1057),
.Y(n_1189)
);

CKINVDCx8_ASAP7_75t_R g1190 ( 
.A(n_999),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1017),
.B(n_1000),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1073),
.B(n_1000),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1020),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1021),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_968),
.A2(n_978),
.B(n_986),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1035),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_986),
.A2(n_1023),
.B(n_1031),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_980),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1026),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1035),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1030),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_963),
.B(n_1069),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1035),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1114),
.A2(n_988),
.B(n_1024),
.Y(n_1205)
);

CKINVDCx11_ASAP7_75t_R g1206 ( 
.A(n_961),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_967),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1016),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_962),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_971),
.A2(n_1013),
.A3(n_1006),
.B(n_1005),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1056),
.B(n_887),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_964),
.B(n_1038),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1214)
);

BUFx4f_ASAP7_75t_SL g1215 ( 
.A(n_1056),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1090),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_964),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_964),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1059),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1101),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1178),
.B(n_1142),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1134),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1144),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1134),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1168),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1158),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1158),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1164),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1154),
.B(n_1156),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1144),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1157),
.B(n_1166),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1176),
.Y(n_1232)
);

OAI21xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1186),
.A2(n_1135),
.B(n_1138),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1178),
.B(n_1182),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1126),
.A2(n_1138),
.B1(n_1175),
.B2(n_1143),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1168),
.B(n_1148),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1146),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1176),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1160),
.A2(n_1151),
.B1(n_1143),
.B2(n_1214),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1182),
.B(n_1179),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1122),
.A2(n_1131),
.B(n_1124),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1120),
.B(n_1151),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1133),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1179),
.B(n_1120),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1213),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1212),
.B(n_1214),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1148),
.B(n_1220),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1164),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1215),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1212),
.B(n_1159),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1177),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1207),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1119),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1119),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1117),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1117),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1155),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1210),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1165),
.B(n_1189),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1121),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1126),
.B(n_1123),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1170),
.Y(n_1264)
);

BUFx2_ASAP7_75t_SL g1265 ( 
.A(n_1201),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1163),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1253),
.B(n_1149),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1246),
.B(n_1240),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1232),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1252),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1253),
.B(n_1149),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1246),
.B(n_1129),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1239),
.B(n_1160),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1229),
.B(n_1132),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1259),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1238),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1244),
.B(n_1221),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1252),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1259),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1263),
.A2(n_1175),
.B1(n_1173),
.B2(n_1150),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1237),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1261),
.B(n_1153),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1266),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1266),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1247),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1254),
.B(n_1153),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1258),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1239),
.B(n_1184),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1235),
.A2(n_1161),
.B1(n_1183),
.B2(n_1206),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1248),
.Y(n_1290)
);

OAI33xp33_ASAP7_75t_L g1291 ( 
.A1(n_1228),
.A2(n_1172),
.A3(n_1218),
.B1(n_1139),
.B2(n_1125),
.B3(n_1118),
.Y(n_1291)
);

INVx4_ASAP7_75t_R g1292 ( 
.A(n_1264),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1234),
.B(n_1180),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1229),
.B(n_1208),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1226),
.B(n_1184),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1250),
.B(n_1127),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1227),
.B(n_1165),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1250),
.B(n_1127),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1223),
.B(n_1174),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1247),
.B(n_1236),
.Y(n_1300)
);

OAI321xp33_ASAP7_75t_L g1301 ( 
.A1(n_1234),
.A2(n_1170),
.A3(n_1188),
.B1(n_1217),
.B2(n_1128),
.C(n_1140),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1269),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1281),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1272),
.B(n_1255),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1270),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1300),
.B(n_1285),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1270),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1287),
.B(n_1258),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1272),
.B(n_1241),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1268),
.B(n_1256),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1296),
.B(n_1241),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1301),
.B(n_1233),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1278),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1296),
.B(n_1241),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1278),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1298),
.B(n_1262),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1268),
.B(n_1256),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1298),
.B(n_1257),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1294),
.B(n_1257),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1274),
.B(n_1262),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1274),
.B(n_1262),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1277),
.B(n_1260),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1279),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1287),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1290),
.B(n_1209),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1300),
.B(n_1247),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1277),
.B(n_1260),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1300),
.B(n_1247),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1305),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1311),
.B(n_1267),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1310),
.B(n_1293),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1305),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1310),
.B(n_1293),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1311),
.B(n_1267),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1307),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1317),
.B(n_1282),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1300),
.Y(n_1337)
);

NAND4xp25_ASAP7_75t_L g1338 ( 
.A(n_1312),
.B(n_1289),
.C(n_1280),
.D(n_1273),
.Y(n_1338)
);

AND2x4_ASAP7_75t_SL g1339 ( 
.A(n_1324),
.B(n_1279),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1311),
.B(n_1314),
.Y(n_1340)
);

NAND2x1_ASAP7_75t_L g1341 ( 
.A(n_1324),
.B(n_1292),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1303),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_R g1343 ( 
.A(n_1324),
.B(n_1136),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1314),
.B(n_1267),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1324),
.B(n_1292),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1317),
.B(n_1318),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1325),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1314),
.B(n_1271),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1306),
.B(n_1285),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1309),
.B(n_1271),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1307),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1309),
.B(n_1271),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1309),
.B(n_1286),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_SL g1354 ( 
.A(n_1341),
.B(n_1209),
.C(n_1199),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1329),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1331),
.B(n_1290),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1331),
.B(n_1320),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1329),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1332),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1340),
.B(n_1304),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1333),
.B(n_1320),
.Y(n_1361)
);

INVxp67_ASAP7_75t_SL g1362 ( 
.A(n_1343),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1340),
.B(n_1312),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1353),
.B(n_1320),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1339),
.A2(n_1302),
.B1(n_1265),
.B2(n_1284),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1347),
.B(n_1338),
.Y(n_1366)
);

NAND4xp25_ASAP7_75t_L g1367 ( 
.A(n_1333),
.B(n_1273),
.C(n_1288),
.D(n_1198),
.Y(n_1367)
);

NAND2x1_ASAP7_75t_L g1368 ( 
.A(n_1337),
.B(n_1302),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1353),
.B(n_1350),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1342),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1339),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_SL g1372 ( 
.A(n_1346),
.B(n_1136),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1341),
.A2(n_1291),
.B1(n_1318),
.B2(n_1231),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1355),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1358),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1370),
.Y(n_1376)
);

O2A1O1Ixp5_ASAP7_75t_SL g1377 ( 
.A1(n_1359),
.A2(n_1299),
.B(n_1351),
.C(n_1332),
.Y(n_1377)
);

AOI211xp5_ASAP7_75t_L g1378 ( 
.A1(n_1354),
.A2(n_1205),
.B(n_1192),
.C(n_1346),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1369),
.B(n_1350),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1369),
.B(n_1330),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1360),
.Y(n_1381)
);

AOI32xp33_ASAP7_75t_L g1382 ( 
.A1(n_1372),
.A2(n_1352),
.A3(n_1344),
.B1(n_1330),
.B2(n_1348),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1366),
.A2(n_1349),
.B1(n_1337),
.B2(n_1336),
.Y(n_1383)
);

NAND2xp33_ASAP7_75t_SL g1384 ( 
.A(n_1368),
.B(n_1345),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1360),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1366),
.A2(n_1367),
.B1(n_1356),
.B2(n_1362),
.C(n_1373),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1363),
.A2(n_1345),
.B(n_1233),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1371),
.A2(n_1337),
.B1(n_1336),
.B2(n_1349),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1357),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1352),
.Y(n_1390)
);

OAI32xp33_ASAP7_75t_L g1391 ( 
.A1(n_1371),
.A2(n_1308),
.A3(n_1284),
.B1(n_1283),
.B2(n_1323),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_1334),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1364),
.B(n_1334),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1386),
.B(n_1365),
.C(n_1288),
.Y(n_1394)
);

OAI211xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1378),
.A2(n_1206),
.B(n_1130),
.C(n_1180),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1384),
.A2(n_1275),
.B(n_1283),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1374),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1383),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1381),
.B(n_1344),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1382),
.A2(n_1291),
.B1(n_1348),
.B2(n_1335),
.C(n_1351),
.Y(n_1400)
);

AOI222xp33_ASAP7_75t_L g1401 ( 
.A1(n_1384),
.A2(n_1231),
.B1(n_1243),
.B2(n_1245),
.C1(n_1275),
.C2(n_1171),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1388),
.A2(n_1349),
.B1(n_1306),
.B2(n_1321),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1390),
.B(n_1370),
.Y(n_1403)
);

OAI21xp33_ASAP7_75t_L g1404 ( 
.A1(n_1385),
.A2(n_1304),
.B(n_1319),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1391),
.A2(n_1387),
.B1(n_1379),
.B2(n_1393),
.Y(n_1405)
);

AOI211xp5_ASAP7_75t_L g1406 ( 
.A1(n_1389),
.A2(n_1199),
.B(n_1216),
.C(n_1167),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1405),
.A2(n_1379),
.B(n_1393),
.C(n_1216),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1398),
.B(n_1390),
.Y(n_1409)
);

AO21x1_ASAP7_75t_L g1410 ( 
.A1(n_1396),
.A2(n_1375),
.B(n_1308),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1397),
.Y(n_1411)
);

OAI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1401),
.A2(n_1392),
.B1(n_1376),
.B2(n_1265),
.C(n_1147),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1395),
.B(n_1167),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1394),
.A2(n_1376),
.B1(n_1306),
.B2(n_1321),
.Y(n_1414)
);

OAI21xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1402),
.A2(n_1377),
.B(n_1276),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1404),
.A2(n_1236),
.B1(n_1224),
.B2(n_1222),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1399),
.A2(n_1306),
.B1(n_1321),
.B2(n_1326),
.Y(n_1417)
);

AOI222xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1406),
.A2(n_1185),
.B1(n_1249),
.B2(n_1152),
.C1(n_1215),
.C2(n_1171),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1403),
.A2(n_1328),
.B1(n_1326),
.B2(n_1316),
.Y(n_1419)
);

OAI211xp5_ASAP7_75t_L g1420 ( 
.A1(n_1405),
.A2(n_1190),
.B(n_1141),
.C(n_1201),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1409),
.B(n_1313),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1411),
.Y(n_1422)
);

AOI211xp5_ASAP7_75t_L g1423 ( 
.A1(n_1420),
.A2(n_1301),
.B(n_1187),
.C(n_1200),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1410),
.B(n_1407),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1415),
.B(n_1418),
.C(n_1412),
.Y(n_1425)
);

NAND4xp25_ASAP7_75t_L g1426 ( 
.A(n_1413),
.B(n_1187),
.C(n_1225),
.D(n_1191),
.Y(n_1426)
);

NOR3xp33_ASAP7_75t_L g1427 ( 
.A(n_1408),
.B(n_1202),
.C(n_1162),
.Y(n_1427)
);

OAI311xp33_ASAP7_75t_L g1428 ( 
.A1(n_1414),
.A2(n_1242),
.A3(n_1297),
.B1(n_1327),
.C1(n_1322),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1417),
.B(n_1342),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1416),
.A2(n_1188),
.B(n_1308),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1416),
.A2(n_1230),
.B(n_1223),
.C(n_1202),
.Y(n_1431)
);

NOR3xp33_ASAP7_75t_L g1432 ( 
.A(n_1425),
.B(n_1162),
.C(n_1196),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_L g1433 ( 
.A(n_1424),
.B(n_1211),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1426),
.B(n_1211),
.Y(n_1434)
);

NOR3xp33_ASAP7_75t_L g1435 ( 
.A(n_1427),
.B(n_1145),
.C(n_1137),
.Y(n_1435)
);

AND5x1_ASAP7_75t_L g1436 ( 
.A(n_1423),
.B(n_1419),
.C(n_1203),
.D(n_1195),
.E(n_1197),
.Y(n_1436)
);

NOR3xp33_ASAP7_75t_L g1437 ( 
.A(n_1431),
.B(n_1145),
.C(n_1137),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1422),
.B(n_1211),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1421),
.B(n_1429),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_SL g1440 ( 
.A(n_1430),
.B(n_1169),
.C(n_1428),
.Y(n_1440)
);

NOR3xp33_ASAP7_75t_L g1441 ( 
.A(n_1425),
.B(n_1219),
.C(n_1204),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1434),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1440),
.A2(n_1152),
.B1(n_1251),
.B2(n_1194),
.C(n_1193),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1432),
.B(n_1313),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1441),
.B(n_1433),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_SL g1446 ( 
.A(n_1439),
.B(n_1435),
.C(n_1437),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1438),
.B(n_1181),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1436),
.B(n_1315),
.Y(n_1448)
);

NAND4xp25_ASAP7_75t_SL g1449 ( 
.A(n_1433),
.B(n_1297),
.C(n_1295),
.D(n_1251),
.Y(n_1449)
);

XOR2xp5_ASAP7_75t_L g1450 ( 
.A(n_1434),
.B(n_1169),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1448),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1444),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1442),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1443),
.Y(n_1454)
);

XNOR2x1_ASAP7_75t_L g1455 ( 
.A(n_1450),
.B(n_1181),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1453),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1451),
.A2(n_1445),
.B(n_1447),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1452),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1456),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_SL g1460 ( 
.A1(n_1459),
.A2(n_1457),
.B(n_1458),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1459),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1460),
.A2(n_1446),
.B(n_1454),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1462),
.A2(n_1461),
.B(n_1455),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1463),
.B(n_1457),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1464),
.A2(n_1455),
.B(n_1449),
.Y(n_1465)
);


endmodule