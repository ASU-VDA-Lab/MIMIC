module fake_netlist_1_4354_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_6), .B(n_4), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_10), .B(n_0), .Y(n_16) );
O2A1O1Ixp33_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_0), .B(n_1), .C(n_2), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_14), .Y(n_18) );
AOI21x1_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_10), .B(n_12), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_18), .B(n_15), .Y(n_20) );
NAND2x1p5_ASAP7_75t_L g21 ( .A(n_19), .B(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NAND2x1_ASAP7_75t_L g23 ( .A(n_20), .B(n_12), .Y(n_23) );
NOR2xp67_ASAP7_75t_L g24 ( .A(n_22), .B(n_1), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_23), .B(n_17), .Y(n_25) );
NOR2xp33_ASAP7_75t_SL g26 ( .A(n_24), .B(n_25), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_21), .B1(n_12), .B2(n_5), .Y(n_27) );
INVxp67_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
NAND2x1p5_ASAP7_75t_L g29 ( .A(n_27), .B(n_2), .Y(n_29) );
NOR2x1_ASAP7_75t_L g30 ( .A(n_26), .B(n_3), .Y(n_30) );
BUFx6f_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
OAI22x1_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_32) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVxp67_ASAP7_75t_SL g34 ( .A(n_33), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_29), .B1(n_32), .B2(n_31), .Y(n_35) );
endmodule