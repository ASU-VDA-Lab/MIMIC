module real_jpeg_4005_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_53),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_1),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_1),
.B(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_3),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_3),
.B(n_303),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_3),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_4),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_4),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_5),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_5),
.B(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_7),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_7),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_7),
.B(n_300),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_8),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_8),
.B(n_349),
.Y(n_348)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_11),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_11),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_12),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_12),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_12),
.B(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_14),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_14),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_14),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_14),
.B(n_351),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_15),
.Y(n_141)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_15),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_16),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

AND2x6_ASAP7_75t_SL g140 ( 
.A(n_16),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_16),
.B(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_314),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_257),
.B(n_313),
.Y(n_19)
);

AOI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_210),
.B(n_256),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_162),
.B(n_209),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_131),
.B(n_161),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_96),
.B(n_130),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_71),
.B(n_95),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_47),
.B(n_70),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_40),
.B(n_46),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_36),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_31),
.Y(n_329)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_32),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_32),
.Y(n_288)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_45),
.Y(n_157)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_45),
.Y(n_220)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_45),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_60),
.C(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_55),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_63),
.Y(n_202)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_94),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_94),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_77),
.C(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_116),
.C(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_83),
.Y(n_237)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_84),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_88),
.Y(n_337)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_90),
.Y(n_242)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_90),
.Y(n_271)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_115),
.C(n_118),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_103),
.C(n_107),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_126),
.C(n_128),
.Y(n_159)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_120),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_125),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_125),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_126),
.Y(n_129)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_160),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_144),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_143),
.C(n_208),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_184),
.C(n_185),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_153),
.C(n_158),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_159),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_207),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_207),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_182),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_165),
.B(n_166),
.C(n_182),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_179),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_230),
.C(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_172),
.C(n_177),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_187),
.C(n_206),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_195),
.B1(n_205),
.B2(n_206),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_190),
.B(n_194),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_190),
.Y(n_194)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_194),
.B(n_214),
.C(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_201),
.C(n_203),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_201),
.Y(n_204)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_255),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_255),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_228),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_227),
.C(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_224),
.B2(n_226),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_216),
.B(n_219),
.C(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_221),
.Y(n_308)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_228),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_233),
.C(n_246),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_246),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_239),
.C(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_251),
.C(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_254),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_311),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_311),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_292),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_261),
.B(n_292),
.C(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_274),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_275),
.C(n_278),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_263),
.B(n_268),
.C(n_272),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_283),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_289),
.C(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_290),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_297),
.B1(n_309),
.B2(n_310),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_310),
.C(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_307),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_302),
.C(n_307),
.Y(n_345)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_358),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_356),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_356),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_342),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_331),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_328),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_341),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_355),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_353),
.B2(n_354),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);


endmodule