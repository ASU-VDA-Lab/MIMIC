module fake_jpeg_6191_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_33),
.B1(n_23),
.B2(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_1),
.C(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_21),
.B1(n_12),
.B2(n_24),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_51),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_29),
.C(n_18),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.C(n_32),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_31),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_45),
.Y(n_60)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_20),
.B(n_19),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.C(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_12),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_52),
.B1(n_44),
.B2(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

OR2x6_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_88),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_41),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_87),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_69),
.C(n_66),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_72),
.B(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_21),
.B1(n_24),
.B2(n_14),
.C(n_30),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_88),
.B(n_69),
.C(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_69),
.B1(n_83),
.B2(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_33),
.B1(n_41),
.B2(n_23),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_111),
.B(n_18),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_94),
.B1(n_91),
.B2(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_33),
.B1(n_16),
.B2(n_19),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_91),
.C(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_109),
.B1(n_103),
.B2(n_102),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_109),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_110),
.C(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_105),
.C(n_16),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_117),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_6),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_123),
.B1(n_119),
.B2(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_11),
.B1(n_7),
.B2(n_5),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_134),
.B1(n_133),
.B2(n_5),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_5),
.Y(n_137)
);


endmodule