module real_jpeg_29930_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_25),
.B1(n_31),
.B2(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_36),
.B1(n_40),
.B2(n_69),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_2),
.A2(n_25),
.B1(n_31),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_25),
.B1(n_31),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_5),
.A2(n_36),
.B1(n_40),
.B2(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_25),
.B1(n_31),
.B2(n_39),
.Y(n_91)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_31),
.A3(n_40),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_36),
.B1(n_40),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_10),
.A2(n_22),
.B(n_65),
.C(n_66),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_25),
.B1(n_31),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_36),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_22),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_13),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_31),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_13),
.B(n_31),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_13),
.B(n_77),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_34),
.B1(n_43),
.B2(n_128),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_70),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_18),
.B(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.C(n_60),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_19),
.A2(n_20),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_33),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.A3(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_26),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_23),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_25),
.A2(n_31),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_29),
.B(n_53),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_29),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_41),
.B2(n_44),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_34),
.A2(n_38),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_34),
.A2(n_41),
.B1(n_121),
.B2(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_35),
.A2(n_42),
.B1(n_45),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_35),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_36),
.B(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_36),
.B(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_42),
.Y(n_116)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_47),
.A2(n_60),
.B1(n_61),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_47),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_53),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_53),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_86),
.B2(n_87),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_139),
.B(n_145),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_117),
.B(n_138),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_113),
.C(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_125),
.B(n_137),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_130),
.B(n_136),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_140),
.B(n_141),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);


endmodule