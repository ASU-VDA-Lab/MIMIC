module fake_jpeg_1546_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_80),
.B(n_122),
.Y(n_151)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g205 ( 
.A(n_89),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_127),
.Y(n_181)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

CKINVDCx6p67_ASAP7_75t_R g182 ( 
.A(n_104),
.Y(n_182)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_37),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_45),
.Y(n_137)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_56),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_8),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

BUFx4f_ASAP7_75t_L g127 ( 
.A(n_21),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_25),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_137),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_56),
.B1(n_60),
.B2(n_58),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_144),
.A2(n_33),
.B1(n_43),
.B2(n_42),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_145),
.B(n_155),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_56),
.B1(n_59),
.B2(n_26),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_161),
.B1(n_166),
.B2(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_60),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_153),
.B(n_0),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_58),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_24),
.B1(n_55),
.B2(n_54),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_172),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_63),
.A2(n_59),
.B1(n_51),
.B2(n_26),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_65),
.A2(n_59),
.B1(n_51),
.B2(n_26),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_22),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_167),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_109),
.A2(n_22),
.B1(n_51),
.B2(n_25),
.Y(n_169)
);

NAND2x1_ASAP7_75t_L g172 ( 
.A(n_92),
.B(n_22),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_21),
.B1(n_25),
.B2(n_55),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_180),
.A2(n_196),
.B1(n_202),
.B2(n_30),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_54),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_194),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_185),
.B(n_0),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_76),
.A2(n_21),
.B1(n_53),
.B2(n_19),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_116),
.B(n_33),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_53),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_127),
.A2(n_52),
.B1(n_48),
.B2(n_43),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_69),
.A2(n_93),
.B1(n_82),
.B2(n_106),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_118),
.A2(n_42),
.B1(n_52),
.B2(n_48),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_73),
.B(n_38),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_19),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_212),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_214),
.Y(n_305)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_135),
.B(n_128),
.C(n_125),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_216),
.B(n_221),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_217),
.A2(n_232),
.B1(n_247),
.B2(n_267),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_89),
.B1(n_101),
.B2(n_94),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_218),
.A2(n_225),
.B1(n_231),
.B2(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_162),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_219),
.B(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_220),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_151),
.B(n_103),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_224),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_97),
.B1(n_91),
.B2(n_90),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_150),
.B1(n_196),
.B2(n_84),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_168),
.B(n_38),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_172),
.B(n_24),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_242),
.B(n_244),
.Y(n_331)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_154),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_190),
.A2(n_88),
.B1(n_30),
.B2(n_3),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_130),
.B(n_138),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_249),
.A2(n_253),
.B(n_260),
.Y(n_310)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_10),
.Y(n_255)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_142),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_262),
.Y(n_330)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_142),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_164),
.Y(n_263)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_200),
.A2(n_6),
.B1(n_1),
.B2(n_4),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_265),
.A2(n_169),
.B(n_184),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_149),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_270),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_186),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_268),
.B(n_269),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_132),
.B(n_146),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_170),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_209),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_271),
.B(n_272),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_140),
.B(n_5),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_190),
.A2(n_5),
.B(n_11),
.C(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_166),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_147),
.B(n_11),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_277),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_180),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_203),
.B1(n_148),
.B2(n_178),
.Y(n_316)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g278 ( 
.A(n_134),
.Y(n_278)
);

CKINVDCx12_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_171),
.B(n_17),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_280),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_281),
.Y(n_291)
);

CKINVDCx6p67_ASAP7_75t_R g282 ( 
.A(n_161),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_17),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_284),
.Y(n_344)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_286),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_296),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_157),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_177),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_298),
.B(n_304),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_210),
.B1(n_163),
.B2(n_159),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_303),
.A2(n_225),
.B1(n_217),
.B2(n_233),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_198),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_254),
.A2(n_192),
.B1(n_187),
.B2(n_141),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_306),
.A2(n_332),
.B(n_345),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_245),
.A2(n_173),
.B1(n_187),
.B2(n_148),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_307),
.A2(n_322),
.B1(n_320),
.B2(n_295),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_230),
.B(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_337),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_324),
.B1(n_227),
.B2(n_239),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_282),
.A2(n_173),
.B1(n_178),
.B2(n_176),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_218),
.A2(n_176),
.B1(n_188),
.B2(n_199),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_237),
.A2(n_197),
.B1(n_131),
.B2(n_210),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_159),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_231),
.A2(n_197),
.B1(n_131),
.B2(n_163),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_293),
.A2(n_213),
.B1(n_229),
.B2(n_267),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_349),
.A2(n_352),
.B1(n_342),
.B2(n_312),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_287),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_350),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_308),
.A2(n_293),
.B1(n_251),
.B2(n_292),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_354),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_288),
.A2(n_213),
.B1(n_229),
.B2(n_265),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_343),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_353),
.B(n_359),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_337),
.A2(n_217),
.B(n_270),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_326),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_361),
.B(n_317),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_216),
.C(n_223),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_365),
.Y(n_410)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_364),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_296),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_326),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_390),
.Y(n_422)
);

AO21x2_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_329),
.B(n_327),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_304),
.B(n_222),
.C(n_214),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_385),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_331),
.B(n_284),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_369),
.B(n_317),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_330),
.B(n_215),
.CI(n_238),
.CON(n_370),
.SN(n_370)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_323),
.B(n_306),
.C(n_338),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_372),
.A2(n_316),
.B1(n_324),
.B2(n_333),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_266),
.B(n_243),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_382),
.B(n_347),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_288),
.A2(n_240),
.B1(n_246),
.B2(n_252),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_375),
.A2(n_378),
.B1(n_332),
.B2(n_318),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_309),
.B(n_224),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_376),
.B(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_314),
.B(n_248),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_303),
.A2(n_281),
.B1(n_273),
.B2(n_259),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_264),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_380),
.B(n_384),
.Y(n_421)
);

INVx11_ASAP7_75t_SL g381 ( 
.A(n_297),
.Y(n_381)
);

BUFx12f_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_290),
.A2(n_236),
.B(n_261),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_310),
.B(n_250),
.Y(n_384)
);

XOR2x2_ASAP7_75t_L g385 ( 
.A(n_298),
.B(n_278),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_290),
.B(n_256),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_388),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_280),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_294),
.B(n_278),
.C(n_280),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_327),
.Y(n_413)
);

AOI32xp33_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_12),
.A3(n_15),
.B1(n_334),
.B2(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_302),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_339),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_392),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_318),
.A2(n_315),
.B(n_345),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_347),
.B(n_313),
.Y(n_414)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_302),
.Y(n_394)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_291),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

INVx3_ASAP7_75t_SL g398 ( 
.A(n_357),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_398),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_400),
.B(n_430),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_401),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_420),
.B1(n_423),
.B2(n_361),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_405),
.A2(n_432),
.B1(n_375),
.B2(n_378),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_339),
.B(n_323),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_408),
.A2(n_411),
.B(n_407),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_315),
.B(n_329),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_385),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_414),
.A2(n_428),
.B(n_363),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_369),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_351),
.A2(n_373),
.B1(n_348),
.B2(n_367),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_425),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_382),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_348),
.A2(n_313),
.B(n_319),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_395),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_352),
.A2(n_312),
.B1(n_342),
.B2(n_328),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_431),
.A2(n_433),
.B(n_393),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_349),
.A2(n_328),
.B1(n_305),
.B2(n_289),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_299),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_359),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_399),
.B(n_402),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_439),
.B(n_447),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_441),
.A2(n_451),
.B1(n_455),
.B2(n_456),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_424),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_442),
.B(n_444),
.Y(n_497)
);

AO22x1_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_354),
.B1(n_351),
.B2(n_385),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_446),
.B(n_465),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_388),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_368),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_457),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_405),
.A2(n_351),
.B1(n_354),
.B2(n_362),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_425),
.A2(n_374),
.B(n_386),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_453),
.A2(n_459),
.B(n_462),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_420),
.A2(n_351),
.B1(n_365),
.B2(n_387),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_397),
.A2(n_371),
.B1(n_390),
.B2(n_386),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_366),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_458),
.B(n_463),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_460),
.A2(n_471),
.B1(n_473),
.B2(n_435),
.Y(n_507)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_414),
.A2(n_363),
.B(n_389),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_411),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_472),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_434),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_418),
.Y(n_466)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_466),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_410),
.B(n_371),
.C(n_383),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_413),
.C(n_419),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_401),
.A2(n_358),
.B(n_364),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_410),
.B(n_355),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_412),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_407),
.B(n_353),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_405),
.A2(n_370),
.B1(n_360),
.B2(n_357),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_412),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_506),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_492),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_451),
.A2(n_397),
.B1(n_432),
.B2(n_405),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_478),
.A2(n_482),
.B1(n_507),
.B2(n_471),
.Y(n_512)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_438),
.A2(n_405),
.B1(n_422),
.B2(n_423),
.Y(n_482)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_485),
.Y(n_508)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_486),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_455),
.A2(n_433),
.B1(n_431),
.B2(n_423),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_487),
.A2(n_490),
.B1(n_438),
.B2(n_473),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_441),
.A2(n_408),
.B1(n_428),
.B2(n_400),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_468),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_496),
.B(n_416),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_439),
.B(n_409),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_502),
.B(n_305),
.Y(n_534)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_443),
.Y(n_503)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_505),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_403),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_509),
.A2(n_505),
.B1(n_503),
.B2(n_481),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_458),
.C(n_454),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_510),
.B(n_516),
.C(n_536),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_512),
.A2(n_533),
.B1(n_501),
.B2(n_494),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_513),
.Y(n_541)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_446),
.CI(n_445),
.CON(n_514),
.SN(n_514)
);

FAx1_ASAP7_75t_SL g542 ( 
.A(n_514),
.B(n_490),
.CI(n_499),
.CON(n_542),
.SN(n_542)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_497),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_515),
.B(n_518),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_454),
.C(n_448),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_480),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_483),
.A2(n_456),
.B1(n_465),
.B2(n_440),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_521),
.A2(n_525),
.B1(n_538),
.B2(n_479),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_491),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_529),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_492),
.B(n_463),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_484),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_482),
.A2(n_459),
.B1(n_462),
.B2(n_453),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_446),
.Y(n_526)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

OAI21x1_ASAP7_75t_SL g561 ( 
.A1(n_527),
.A2(n_532),
.B(n_415),
.Y(n_561)
);

INVx11_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_528),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_499),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_489),
.A2(n_437),
.B(n_426),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_478),
.A2(n_437),
.B1(n_396),
.B2(n_426),
.Y(n_533)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_534),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_484),
.B(n_436),
.C(n_394),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_370),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_537),
.B(n_500),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_504),
.A2(n_436),
.B1(n_398),
.B2(n_470),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_539),
.B(n_555),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_540),
.A2(n_550),
.B1(n_556),
.B2(n_559),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_545),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_513),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_517),
.B(n_489),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_553),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_547),
.A2(n_526),
.B1(n_530),
.B2(n_532),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_477),
.Y(n_549)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_549),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_509),
.A2(n_501),
.B1(n_476),
.B2(n_493),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_538),
.Y(n_551)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_551),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_486),
.Y(n_554)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_498),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_531),
.A2(n_485),
.B1(n_476),
.B2(n_495),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_520),
.B(n_510),
.C(n_536),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_558),
.B(n_561),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_531),
.A2(n_470),
.B1(n_427),
.B2(n_415),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_560),
.Y(n_566)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_562),
.B(n_511),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_516),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_564),
.B(n_570),
.Y(n_591)
);

XNOR2x1_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_526),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_567),
.B(n_572),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_539),
.B(n_520),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_558),
.B(n_524),
.Y(n_572)
);

INVx6_ASAP7_75t_L g573 ( 
.A(n_548),
.Y(n_573)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_573),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_557),
.B(n_533),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_578),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_557),
.B(n_537),
.C(n_508),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_580),
.C(n_552),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_523),
.C(n_519),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_549),
.B(n_514),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_582),
.B(n_583),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_544),
.A2(n_523),
.B1(n_519),
.B2(n_511),
.Y(n_583)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_584),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_568),
.A2(n_541),
.B(n_552),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_592),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_596),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_550),
.Y(n_587)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_576),
.A2(n_542),
.B(n_554),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_590),
.B(n_593),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_582),
.A2(n_540),
.B(n_542),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_556),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_543),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_595),
.B(n_409),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_553),
.C(n_563),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_565),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_598),
.B(n_601),
.Y(n_610)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_573),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_575),
.B(n_563),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_560),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_595),
.A2(n_579),
.B(n_571),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_603),
.A2(n_608),
.B(n_611),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_572),
.C(n_564),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_607),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_569),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_SL g608 ( 
.A(n_591),
.B(n_567),
.Y(n_608)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_609),
.Y(n_624)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_514),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_569),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_613),
.Y(n_625)
);

MAJx2_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_570),
.C(n_566),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_615),
.A2(n_600),
.B1(n_588),
.B2(n_585),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_596),
.C(n_587),
.Y(n_617)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_617),
.Y(n_630)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_618),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_616),
.B(n_597),
.Y(n_619)
);

AOI21xp33_ASAP7_75t_L g631 ( 
.A1(n_619),
.A2(n_627),
.B(n_614),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_611),
.B(n_590),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_621),
.B(n_623),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_614),
.A2(n_589),
.B1(n_587),
.B2(n_593),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_622),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_610),
.B(n_391),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_604),
.B(n_592),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_626),
.A2(n_604),
.B(n_619),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_629),
.A2(n_631),
.B(n_627),
.Y(n_637)
);

NAND4xp25_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_615),
.C(n_528),
.D(n_379),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_632),
.B(n_617),
.C(n_625),
.Y(n_635)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_635),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_630),
.B(n_624),
.C(n_622),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_637),
.C(n_638),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_628),
.Y(n_638)
);

OAI321xp33_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_633),
.A3(n_634),
.B1(n_427),
.B2(n_289),
.C(n_301),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_634),
.C(n_639),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_299),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_301),
.Y(n_644)
);


endmodule