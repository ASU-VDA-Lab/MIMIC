module fake_netlist_1_732_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_6), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_7), .B(n_5), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_0), .B(n_8), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_2), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
BUFx4f_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_15), .Y(n_21) );
INVx5_ASAP7_75t_L g22 ( .A(n_10), .Y(n_22) );
NOR2xp67_ASAP7_75t_L g23 ( .A(n_13), .B(n_2), .Y(n_23) );
CKINVDCx6p67_ASAP7_75t_R g24 ( .A(n_22), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_10), .Y(n_25) );
BUFx12f_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
AND4x1_ASAP7_75t_L g28 ( .A(n_25), .B(n_17), .C(n_16), .D(n_18), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_25), .B(n_23), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_24), .B(n_20), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OAI31xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_19), .A3(n_27), .B(n_21), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_30), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B1(n_20), .B2(n_16), .Y(n_34) );
OAI21xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_29), .B(n_28), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_33), .B(n_30), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_33), .Y(n_37) );
NOR3xp33_ASAP7_75t_SL g38 ( .A(n_35), .B(n_14), .C(n_11), .Y(n_38) );
AND2x2_ASAP7_75t_L g39 ( .A(n_37), .B(n_26), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_38), .B1(n_36), .B2(n_9), .Y(n_41) );
endmodule