module real_jpeg_25967_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_4),
.A2(n_25),
.B(n_45),
.C(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_24),
.B(n_79),
.C(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_4),
.A2(n_38),
.B1(n_82),
.B2(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_4),
.B(n_33),
.C(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_4),
.B(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_29),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_4),
.B(n_65),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_21),
.B1(n_25),
.B2(n_38),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_21),
.B1(n_25),
.B2(n_35),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_8),
.A2(n_21),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_55),
.B1(n_82),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_10),
.Y(n_86)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_11),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_11),
.B(n_140),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_114),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_73),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_16),
.B(n_73),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_56),
.C(n_60),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_17),
.B(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_26),
.C(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_21),
.A2(n_25),
.B1(n_45),
.B2(n_49),
.Y(n_52)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_23),
.A2(n_25),
.B(n_38),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_24),
.B1(n_93),
.B2(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_27),
.B(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_30),
.A2(n_37),
.B(n_39),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_32),
.A2(n_33),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_33),
.B(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_36),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_37),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_46),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_39),
.B(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_43),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_47),
.B1(n_66),
.B2(n_67),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_47),
.B(n_124),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_51),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_56),
.B(n_60),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_57),
.A2(n_59),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_57),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_59),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_64),
.B(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_63),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_65),
.B(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_69),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_71),
.B(n_131),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_88),
.B2(n_89),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_101),
.B1(n_102),
.B2(n_112),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_174),
.B(n_178),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_160),
.B(n_173),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_142),
.B(n_159),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_134),
.B2(n_141),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_128),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_133),
.C(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_148),
.B(n_158),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_154),
.B(n_157),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_162),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_168),
.C(n_170),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_176),
.Y(n_178)
);


endmodule