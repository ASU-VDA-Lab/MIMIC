module fake_jpeg_13663_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_15),
.B1(n_13),
.B2(n_2),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_31),
.B1(n_53),
.B2(n_49),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_60),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_62),
.B(n_73),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_1),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_82),
.B(n_105),
.Y(n_146)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_39),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_90),
.Y(n_152)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_9),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_6),
.Y(n_112)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_100),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_6),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_23),
.B1(n_31),
.B2(n_29),
.Y(n_153)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_104),
.Y(n_140)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_38),
.B(n_4),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_5),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_107),
.B(n_26),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_42),
.B(n_5),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_41),
.B(n_8),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_174),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_33),
.B1(n_52),
.B2(n_50),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_113),
.A2(n_116),
.B1(n_131),
.B2(n_143),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_53),
.B1(n_49),
.B2(n_44),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_114),
.A2(n_137),
.B1(n_153),
.B2(n_119),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_33),
.B1(n_52),
.B2(n_50),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_133),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_129),
.B(n_162),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_32),
.B1(n_48),
.B2(n_45),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_132),
.A2(n_152),
.B1(n_158),
.B2(n_123),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_54),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_55),
.A2(n_29),
.B1(n_44),
.B2(n_37),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_54),
.B1(n_48),
.B2(n_45),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_22),
.B(n_34),
.C(n_27),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_144),
.A2(n_139),
.B(n_117),
.C(n_126),
.Y(n_197)
);

AO22x2_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_40),
.B1(n_34),
.B2(n_8),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_139),
.B(n_144),
.C(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_40),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_21),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_57),
.B(n_21),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_58),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_65),
.B(n_26),
.Y(n_171)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_63),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_56),
.A2(n_37),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_173),
.A2(n_127),
.B1(n_150),
.B2(n_142),
.Y(n_226)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_75),
.B1(n_86),
.B2(n_67),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_182),
.A2(n_184),
.B1(n_186),
.B2(n_217),
.Y(n_251)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_72),
.B1(n_80),
.B2(n_98),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_106),
.B1(n_66),
.B2(n_68),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_187),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_56),
.B1(n_171),
.B2(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_191),
.B1(n_206),
.B2(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_190),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_124),
.A2(n_156),
.B(n_121),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_127),
.B(n_161),
.Y(n_230)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_194),
.B(n_199),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_112),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_209),
.Y(n_262)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_138),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_203),
.B(n_208),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_133),
.B(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_132),
.B1(n_130),
.B2(n_147),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_147),
.A2(n_111),
.B1(n_157),
.B2(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_136),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_122),
.B(n_136),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_222),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_123),
.A2(n_145),
.B1(n_142),
.B2(n_154),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_163),
.B1(n_170),
.B2(n_222),
.Y(n_242)
);

OR2x4_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_215),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_125),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_111),
.B(n_157),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_208),
.B1(n_195),
.B2(n_204),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_145),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_150),
.C(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_175),
.C(n_211),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_225),
.B(n_227),
.Y(n_259)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_221),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_230),
.B(n_265),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_238),
.A2(n_247),
.B1(n_251),
.B2(n_256),
.Y(n_285)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_135),
.A3(n_154),
.B1(n_163),
.B2(n_161),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_246),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_195),
.B1(n_204),
.B2(n_191),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_243),
.A2(n_234),
.B1(n_268),
.B2(n_232),
.Y(n_272)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_197),
.A3(n_219),
.B1(n_214),
.B2(n_212),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_179),
.A2(n_218),
.B1(n_192),
.B2(n_180),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_193),
.B(n_224),
.C(n_176),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_247),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_180),
.A2(n_188),
.B1(n_185),
.B2(n_194),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_259),
.A2(n_236),
.B1(n_244),
.B2(n_250),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_264),
.C(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_187),
.Y(n_264)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_178),
.A3(n_181),
.B1(n_201),
.B2(n_177),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_210),
.B(n_183),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_267),
.B(n_266),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_270),
.B(n_284),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_283),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_274),
.B1(n_228),
.B2(n_240),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_234),
.A2(n_243),
.B1(n_232),
.B2(n_238),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_246),
.A2(n_231),
.B(n_259),
.C(n_249),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_275),
.A2(n_287),
.B(n_276),
.C(n_296),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_295),
.C(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_280),
.B(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_286),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_255),
.B1(n_263),
.B2(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_254),
.B1(n_228),
.B2(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_253),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_291),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_300),
.B1(n_254),
.B2(n_266),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_250),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_270),
.B(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_235),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_299),
.C(n_284),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_235),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_239),
.B(n_242),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_313),
.B(n_317),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_309),
.B1(n_312),
.B2(n_319),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_308),
.A2(n_318),
.B1(n_324),
.B2(n_314),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_285),
.A2(n_241),
.B1(n_236),
.B2(n_244),
.Y(n_309)
);

AOI22x1_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_281),
.B1(n_275),
.B2(n_272),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_293),
.B1(n_294),
.B2(n_277),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_298),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_282),
.B1(n_269),
.B2(n_276),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_315),
.A2(n_299),
.B(n_283),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_269),
.B(n_287),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_282),
.B1(n_280),
.B2(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_286),
.B1(n_280),
.B2(n_290),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_291),
.B1(n_297),
.B2(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_288),
.Y(n_329)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_289),
.C(n_278),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_331),
.C(n_336),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_304),
.B(n_277),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_343),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_334),
.A2(n_309),
.B1(n_304),
.B2(n_305),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_322),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_301),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_312),
.C(n_314),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_303),
.Y(n_338)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_340),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_320),
.Y(n_339)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_310),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_317),
.B1(n_320),
.B2(n_307),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_346),
.A2(n_356),
.B1(n_362),
.B2(n_342),
.Y(n_373)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_357),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_321),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_321),
.Y(n_354)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_302),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_337),
.A2(n_315),
.B1(n_302),
.B2(n_325),
.Y(n_356)
);

OAI22x1_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_315),
.B1(n_325),
.B2(n_328),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_329),
.A2(n_339),
.B1(n_330),
.B2(n_345),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_344),
.B(n_340),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_365),
.A2(n_358),
.B(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_369),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_330),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_338),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_375),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_342),
.B1(n_334),
.B2(n_315),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_372),
.A2(n_373),
.B1(n_344),
.B2(n_349),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_331),
.C(n_336),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_350),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_347),
.B(n_341),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_374),
.B(n_359),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_379),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_361),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_381),
.C(n_383),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_370),
.B(n_358),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_363),
.A2(n_353),
.B1(n_361),
.B2(n_360),
.Y(n_382)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_385),
.A2(n_372),
.B1(n_364),
.B2(n_365),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_373),
.B1(n_364),
.B2(n_363),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_390),
.B1(n_362),
.B2(n_356),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_343),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_385),
.A2(n_369),
.B1(n_366),
.B2(n_367),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_394),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_391),
.A2(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_396),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_384),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_341),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_397),
.A2(n_398),
.B(n_394),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_360),
.B1(n_353),
.B2(n_371),
.Y(n_398)
);

FAx1_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_392),
.CI(n_381),
.CON(n_399),
.SN(n_399)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_392),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_404),
.B(n_401),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_386),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_402),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_407),
.Y(n_408)
);

AOI322xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_403),
.A3(n_398),
.B1(n_389),
.B2(n_399),
.C1(n_393),
.C2(n_376),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_399),
.C(n_380),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_315),
.Y(n_411)
);


endmodule