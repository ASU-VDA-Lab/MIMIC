module fake_jpeg_15510_n_335 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_44),
.B(n_45),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_62),
.Y(n_76)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_6),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_61),
.B(n_63),
.Y(n_118)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_13),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_13),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_37),
.B(n_31),
.Y(n_113)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_92),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_78),
.B(n_84),
.Y(n_127)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_21),
.B1(n_23),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_87),
.B1(n_100),
.B2(n_101),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_21),
.B1(n_18),
.B2(n_33),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_21),
.B1(n_32),
.B2(n_28),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_101)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_27),
.C(n_38),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_27),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_117),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_39),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_106),
.A2(n_112),
.B1(n_114),
.B2(n_36),
.Y(n_147)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_47),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_24),
.B1(n_39),
.B2(n_20),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_69),
.B(n_59),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_48),
.A2(n_37),
.B1(n_22),
.B2(n_12),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_44),
.A2(n_11),
.B(n_12),
.C(n_10),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_124),
.B(n_148),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_128),
.A2(n_134),
.B1(n_152),
.B2(n_155),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_58),
.B1(n_65),
.B2(n_62),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_160),
.B1(n_136),
.B2(n_96),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_45),
.Y(n_130)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_43),
.Y(n_132)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g133 ( 
.A1(n_87),
.A2(n_51),
.B1(n_50),
.B2(n_27),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_137),
.B1(n_107),
.B2(n_99),
.Y(n_167)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_67),
.B1(n_53),
.B2(n_38),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_38),
.B1(n_36),
.B2(n_20),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_4),
.B(n_133),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_145),
.Y(n_199)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_156),
.B1(n_161),
.B2(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_10),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_12),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_11),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_157),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_36),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_0),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_137),
.CI(n_150),
.CON(n_197),
.SN(n_197)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_116),
.B(n_27),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_104),
.C(n_27),
.Y(n_165)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_86),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_159),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_164),
.A2(n_167),
.B1(n_183),
.B2(n_172),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_187),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_107),
.B1(n_90),
.B2(n_82),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_126),
.B1(n_146),
.B2(n_128),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_90),
.B1(n_103),
.B2(n_95),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_172),
.A2(n_176),
.B1(n_181),
.B2(n_186),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_95),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_182),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_93),
.B1(n_75),
.B2(n_91),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_93),
.B1(n_75),
.B2(n_3),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_178)
);

XOR2x2_ASAP7_75t_SL g225 ( 
.A(n_178),
.B(n_200),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_0),
.C(n_3),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_4),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_133),
.B1(n_129),
.B2(n_136),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_135),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_129),
.A2(n_134),
.B1(n_161),
.B2(n_126),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_190),
.B1(n_185),
.B2(n_164),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_129),
.A2(n_138),
.B1(n_155),
.B2(n_152),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_119),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_197),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_121),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_196),
.C(n_169),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_143),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_214),
.B1(n_221),
.B2(n_234),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_151),
.B(n_120),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_206),
.A2(n_219),
.B(n_225),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_207),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_215),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_189),
.B1(n_174),
.B2(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_173),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_176),
.B1(n_197),
.B2(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_175),
.B(n_182),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_175),
.B(n_195),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_229),
.B1(n_207),
.B2(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_181),
.B1(n_190),
.B2(n_167),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_240),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_178),
.Y(n_242)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_177),
.B(n_180),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_262),
.B(n_258),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_213),
.B1(n_232),
.B2(n_225),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_255),
.B1(n_240),
.B2(n_243),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_236),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_239),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_211),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_233),
.B1(n_212),
.B2(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_263),
.A2(n_261),
.B1(n_251),
.B2(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_256),
.C(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_270),
.C(n_277),
.Y(n_293)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_250),
.A3(n_242),
.B1(n_252),
.B2(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_273),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_241),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_248),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_241),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_270),
.B(n_263),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_251),
.B1(n_247),
.B2(n_249),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_276),
.B1(n_265),
.B2(n_274),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_249),
.B(n_265),
.C(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_297),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_278),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_280),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_272),
.C(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_301),
.B(n_306),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_268),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_304),
.C(n_286),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_308),
.B(n_285),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_287),
.B(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_276),
.B1(n_275),
.B2(n_280),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_296),
.B1(n_292),
.B2(n_294),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_317),
.B(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_298),
.C(n_293),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_292),
.C(n_294),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_296),
.B(n_289),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_310),
.Y(n_325)
);

NAND4xp25_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_299),
.C(n_290),
.D(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_326),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_320),
.B(n_308),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_317),
.B(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_297),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_322),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_307),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.C(n_325),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_328),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_314),
.Y(n_335)
);


endmodule