module fake_jpeg_24017_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_76),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_51),
.B(n_52),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_28),
.B1(n_31),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_65),
.B1(n_66),
.B2(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_31),
.B1(n_23),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_35),
.B1(n_18),
.B2(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_35),
.B1(n_18),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_32),
.B1(n_29),
.B2(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_84),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_88),
.B(n_95),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_29),
.B1(n_49),
.B2(n_34),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_97),
.Y(n_128)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_64),
.B1(n_54),
.B2(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_101),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_17),
.B1(n_34),
.B2(n_26),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_102),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_17),
.B1(n_34),
.B2(n_26),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_22),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_17),
.B1(n_34),
.B2(n_26),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_22),
.B1(n_39),
.B2(n_42),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_73),
.Y(n_126)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_116),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_17),
.B1(n_5),
.B2(n_10),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_79),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_118),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_126),
.A2(n_138),
.B1(n_152),
.B2(n_146),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_69),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_139),
.B(n_141),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_54),
.B1(n_64),
.B2(n_52),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_140),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_136),
.Y(n_159)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_82),
.A2(n_61),
.B1(n_72),
.B2(n_51),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_66),
.B(n_53),
.C(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_68),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_42),
.B(n_39),
.C(n_80),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_94),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_84),
.B1(n_92),
.B2(n_105),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_81),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_63),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_56),
.B(n_42),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_115),
.C(n_110),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_54),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_112),
.B(n_87),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_164),
.B(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_158),
.B(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_172),
.B1(n_139),
.B2(n_126),
.Y(n_190)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_169),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_143),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_115),
.B1(n_93),
.B2(n_91),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_185),
.B1(n_133),
.B2(n_147),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_171),
.B(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_112),
.B1(n_83),
.B2(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_83),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_117),
.B(n_118),
.C(n_108),
.D(n_116),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.C(n_125),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_123),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_141),
.B(n_152),
.C(n_138),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_192),
.B1(n_161),
.B2(n_141),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_195),
.B1(n_175),
.B2(n_130),
.Y(n_230)
);

CKINVDCx12_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_124),
.B1(n_127),
.B2(n_130),
.Y(n_195)
);

OR2x2_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_142),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_197),
.B(n_153),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_150),
.B(n_140),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_8),
.CI(n_13),
.CON(n_236),
.SN(n_236)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.Y(n_220)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_178),
.B(n_158),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_178),
.B(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_211),
.B1(n_185),
.B2(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_230),
.B1(n_238),
.B2(n_210),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_228),
.B1(n_229),
.B2(n_196),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_240),
.B1(n_194),
.B2(n_215),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_164),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_227),
.C(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_181),
.B1(n_173),
.B2(n_171),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_233),
.B1(n_188),
.B2(n_209),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_226),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_179),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_164),
.B(n_168),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_141),
.B1(n_177),
.B2(n_156),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_167),
.A3(n_141),
.B1(n_125),
.B2(n_155),
.C1(n_134),
.C2(n_119),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_151),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_99),
.B1(n_120),
.B2(n_144),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_199),
.B(n_188),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_10),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_198),
.C(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_254),
.B1(n_256),
.B2(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_186),
.C(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_260),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_218),
.A2(n_186),
.B1(n_207),
.B2(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_259),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_202),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_213),
.C(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_202),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_200),
.B(n_1),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_265),
.A2(n_268),
.B1(n_270),
.B2(n_273),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_228),
.B1(n_217),
.B2(n_223),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_236),
.B1(n_191),
.B2(n_219),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_243),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_275),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_239),
.B1(n_205),
.B2(n_219),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_193),
.B1(n_203),
.B2(n_206),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_227),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_236),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_249),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_203),
.B1(n_120),
.B2(n_200),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_258),
.B(n_255),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_244),
.B1(n_248),
.B2(n_262),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_275),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_254),
.C(n_252),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_293),
.C(n_276),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_242),
.B(n_10),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_294),
.B(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_0),
.C(n_1),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_264),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_291),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_274),
.B(n_270),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.C(n_287),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_304),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_266),
.B1(n_269),
.B2(n_265),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_277),
.C(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_301),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_292),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_287),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_282),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_284),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_296),
.B1(n_285),
.B2(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_6),
.B(n_8),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

AOI31xp67_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_313),
.A3(n_6),
.B(n_4),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_316),
.B(n_6),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

OAI221xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_325),
.B1(n_323),
.B2(n_321),
.C(n_318),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_3),
.B(n_4),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_3),
.Y(n_329)
);


endmodule