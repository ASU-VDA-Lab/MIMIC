module fake_jpeg_19568_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_19),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_18),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_47),
.C(n_41),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_30),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_90),
.B1(n_93),
.B2(n_45),
.Y(n_106)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_19),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_91),
.C(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_35),
.B(n_20),
.C(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_95),
.Y(n_112)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_23),
.B1(n_33),
.B2(n_45),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_47),
.C(n_37),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_23),
.B1(n_33),
.B2(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_23),
.B1(n_40),
.B2(n_47),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_50),
.B1(n_68),
.B2(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_127),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_110),
.B1(n_118),
.B2(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_91),
.B1(n_77),
.B2(n_86),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_83),
.B1(n_76),
.B2(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_49),
.B1(n_40),
.B2(n_47),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_46),
.C(n_39),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_46),
.C(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_124),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_40),
.B1(n_63),
.B2(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_64),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_31),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_43),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_71),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_133),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_46),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_143),
.B(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_138),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_12),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_89),
.B1(n_87),
.B2(n_94),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_152),
.Y(n_160)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_89),
.B1(n_94),
.B2(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_82),
.B1(n_50),
.B2(n_37),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_99),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_39),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_96),
.B1(n_37),
.B2(n_39),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_43),
.B1(n_85),
.B2(n_26),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_34),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_70),
.B1(n_34),
.B2(n_41),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_122),
.B1(n_115),
.B2(n_105),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_115),
.B1(n_108),
.B2(n_123),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_28),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_171),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_116),
.C(n_117),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_169),
.C(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_126),
.B1(n_121),
.B2(n_100),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_174),
.B1(n_182),
.B2(n_184),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_101),
.B(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_186),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_101),
.C(n_41),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_43),
.C(n_123),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_120),
.B1(n_43),
.B2(n_32),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_172),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_26),
.C(n_17),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_180),
.B(n_156),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_31),
.B1(n_17),
.B2(n_25),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_36),
.B1(n_21),
.B2(n_18),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_132),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_138),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_21),
.B(n_18),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_36),
.C(n_28),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_137),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_195),
.B(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

OR2x4_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_145),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_172),
.B(n_159),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_131),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_140),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_141),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_180),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_135),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_149),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_218),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_130),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_170),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_230),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_232),
.B(n_243),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_159),
.B(n_172),
.C(n_177),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_200),
.B1(n_197),
.B2(n_192),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_195),
.B1(n_218),
.B2(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_193),
.B1(n_191),
.B2(n_190),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_163),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_186),
.B(n_184),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_189),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_203),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_256),
.B1(n_260),
.B2(n_233),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_201),
.B1(n_214),
.B2(n_196),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_201),
.B1(n_210),
.B2(n_198),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_253),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_198),
.B1(n_191),
.B2(n_202),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_225),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_208),
.B1(n_171),
.B2(n_155),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_188),
.C(n_28),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_259),
.C(n_262),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_188),
.C(n_21),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_226),
.C(n_237),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_10),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_275),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_225),
.B(n_235),
.C(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_224),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_234),
.C(n_221),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_239),
.B(n_236),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_281),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_241),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_221),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_267),
.B1(n_236),
.B2(n_264),
.C(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_255),
.B1(n_235),
.B2(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_282),
.Y(n_306)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_236),
.B(n_265),
.C(n_246),
.D(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_222),
.B1(n_236),
.B2(n_234),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_222),
.B1(n_258),
.B2(n_266),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_293),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_299),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_11),
.C(n_5),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_270),
.C(n_273),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_289),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_275),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_12),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_298),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_12),
.C(n_5),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_16),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_13),
.B(n_6),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_15),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_285),
.B1(n_297),
.B2(n_291),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_305),
.B1(n_307),
.B2(n_304),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_290),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_300),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_300),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_326),
.A2(n_327),
.B(n_312),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_306),
.B(n_310),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_331),
.B(n_324),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_7),
.B(n_8),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_326),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_328),
.C(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_7),
.C(n_8),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_14),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_14),
.B(n_1),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_1),
.Y(n_338)
);


endmodule