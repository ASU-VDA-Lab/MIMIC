module real_aes_2607_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_0), .B(n_212), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_1), .A2(n_220), .B(n_225), .Y(n_219) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_2), .A2(n_58), .B1(n_93), .B2(n_97), .Y(n_96) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_3), .B(n_227), .Y(n_266) );
INVx1_ASAP7_75t_L g193 ( .A(n_4), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_5), .B(n_227), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_6), .A2(n_55), .B1(n_152), .B2(n_155), .Y(n_151) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_7), .A2(n_22), .B1(n_93), .B2(n_94), .Y(n_92) );
NAND2xp33_ASAP7_75t_L g309 ( .A(n_8), .B(n_229), .Y(n_309) );
INVx2_ASAP7_75t_L g209 ( .A(n_9), .Y(n_209) );
AOI221x1_ASAP7_75t_L g251 ( .A1(n_10), .A2(n_16), .B1(n_212), .B2(n_220), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_11), .B(n_212), .Y(n_305) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_12), .A2(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_13), .B(n_231), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_14), .B(n_227), .Y(n_240) );
AO21x1_ASAP7_75t_L g261 ( .A1(n_15), .A2(n_212), .B(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_16), .A2(n_81), .B1(n_82), .B2(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_16), .Y(n_523) );
NAND2x1_ASAP7_75t_L g283 ( .A(n_17), .B(n_227), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_18), .A2(n_35), .B1(n_136), .B2(n_140), .Y(n_135) );
NAND2x1_ASAP7_75t_L g316 ( .A(n_19), .B(n_229), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_20), .A2(n_38), .B1(n_144), .B2(n_146), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g85 ( .A1(n_21), .A2(n_48), .B1(n_86), .B2(n_107), .Y(n_85) );
OAI221xp5_ASAP7_75t_L g185 ( .A1(n_22), .A2(n_58), .B1(n_63), .B2(n_186), .C(n_188), .Y(n_185) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_23), .A2(n_68), .B(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g233 ( .A(n_23), .B(n_68), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_24), .B(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_26), .B(n_227), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_27), .B(n_229), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_28), .A2(n_56), .B1(n_160), .B2(n_162), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_29), .A2(n_220), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_SL g102 ( .A(n_30), .Y(n_102) );
INVx1_ASAP7_75t_L g195 ( .A(n_31), .Y(n_195) );
AND2x2_ASAP7_75t_L g218 ( .A(n_31), .B(n_193), .Y(n_218) );
AND2x2_ASAP7_75t_L g221 ( .A(n_31), .B(n_222), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_32), .A2(n_65), .B1(n_175), .B2(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_32), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_32), .B(n_212), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_33), .A2(n_39), .B1(n_128), .B2(n_131), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_34), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_36), .B(n_229), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_37), .A2(n_74), .B1(n_172), .B2(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_37), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_40), .A2(n_220), .B(n_315), .Y(n_314) );
AO22x2_ASAP7_75t_L g105 ( .A1(n_41), .A2(n_63), .B1(n_93), .B2(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_42), .B(n_123), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_43), .A2(n_60), .B1(n_112), .B2(n_116), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_44), .B(n_229), .Y(n_284) );
INVx1_ASAP7_75t_L g215 ( .A(n_45), .Y(n_215) );
INVx1_ASAP7_75t_L g224 ( .A(n_45), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_46), .A2(n_54), .B1(n_180), .B2(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_46), .Y(n_181) );
INVx1_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_49), .A2(n_81), .B1(n_82), .B2(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_49), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_50), .B(n_227), .Y(n_254) );
INVx1_ASAP7_75t_L g541 ( .A(n_50), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_51), .A2(n_220), .B(n_282), .Y(n_281) );
AO21x1_ASAP7_75t_L g263 ( .A1(n_52), .A2(n_220), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_53), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g180 ( .A(n_54), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_57), .B(n_212), .Y(n_318) );
INVxp33_ASAP7_75t_L g190 ( .A(n_58), .Y(n_190) );
AND2x2_ASAP7_75t_L g277 ( .A(n_59), .B(n_232), .Y(n_277) );
INVx1_ASAP7_75t_L g217 ( .A(n_61), .Y(n_217) );
INVx1_ASAP7_75t_L g222 ( .A(n_61), .Y(n_222) );
AND2x2_ASAP7_75t_L g320 ( .A(n_62), .B(n_206), .Y(n_320) );
INVxp67_ASAP7_75t_L g189 ( .A(n_63), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g80 ( .A1(n_64), .A2(n_81), .B1(n_82), .B2(n_166), .Y(n_80) );
INVx1_ASAP7_75t_L g166 ( .A(n_64), .Y(n_166) );
INVx1_ASAP7_75t_L g175 ( .A(n_65), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_65), .B(n_212), .Y(n_242) );
AND2x2_ASAP7_75t_L g205 ( .A(n_66), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g262 ( .A(n_67), .B(n_236), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_69), .B(n_229), .Y(n_241) );
AND2x2_ASAP7_75t_L g286 ( .A(n_70), .B(n_206), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_71), .B(n_227), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_72), .A2(n_220), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_73), .B(n_229), .Y(n_253) );
INVx1_ASAP7_75t_L g172 ( .A(n_74), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_75), .B(n_227), .Y(n_226) );
BUFx2_ASAP7_75t_SL g187 ( .A(n_76), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_77), .A2(n_220), .B(n_307), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_182), .B1(n_196), .B2(n_516), .C(n_521), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_167), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_121), .C(n_150), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_111), .Y(n_84) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx8_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
AND2x2_ASAP7_75t_L g114 ( .A(n_90), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g125 ( .A(n_90), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g154 ( .A(n_90), .B(n_139), .Y(n_154) );
AND2x4_ASAP7_75t_L g90 ( .A(n_91), .B(n_95), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g110 ( .A(n_92), .B(n_96), .Y(n_110) );
INVx1_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
AND2x4_ASAP7_75t_L g130 ( .A(n_92), .B(n_95), .Y(n_130) );
INVx2_ASAP7_75t_L g94 ( .A(n_93), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
OAI22x1_ASAP7_75t_L g100 ( .A1(n_93), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_93), .Y(n_101) );
INVx1_ASAP7_75t_L g106 ( .A(n_93), .Y(n_106) );
INVxp67_ASAP7_75t_L g134 ( .A(n_95), .Y(n_134) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g119 ( .A(n_96), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g118 ( .A(n_98), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g158 ( .A(n_98), .B(n_130), .Y(n_158) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_104), .Y(n_98) );
AND2x2_ASAP7_75t_L g115 ( .A(n_99), .B(n_105), .Y(n_115) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g126 ( .A(n_100), .B(n_105), .Y(n_126) );
AND2x2_ASAP7_75t_L g139 ( .A(n_100), .B(n_104), .Y(n_139) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_100), .Y(n_142) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g141 ( .A(n_110), .B(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g164 ( .A(n_110), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g129 ( .A(n_115), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g161 ( .A(n_115), .B(n_119), .Y(n_161) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx8_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g145 ( .A(n_119), .B(n_139), .Y(n_145) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_127), .C(n_135), .D(n_143), .Y(n_121) );
INVx4_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx6_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g133 ( .A(n_126), .B(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g147 ( .A(n_126), .B(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g138 ( .A(n_130), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx6_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx12f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_159), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx5_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B1(n_178), .B2(n_179), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B1(n_174), .B2(n_177), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_174), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
AND3x1_ASAP7_75t_SL g184 ( .A(n_185), .B(n_191), .C(n_194), .Y(n_184) );
INVxp67_ASAP7_75t_L g529 ( .A(n_185), .Y(n_529) );
CKINVDCx8_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_191), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_191), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_SL g534 ( .A(n_192), .B(n_194), .Y(n_534) );
AND2x2_ASAP7_75t_L g539 ( .A(n_192), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g223 ( .A(n_193), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_194), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1p5_ASAP7_75t_L g518 ( .A(n_195), .B(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
NOR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_403), .Y(n_198) );
AO211x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_245), .B(n_296), .C(n_371), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVxp67_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND3x2_ASAP7_75t_L g452 ( .A(n_202), .B(n_333), .C(n_349), .Y(n_452) );
AND2x4_ASAP7_75t_L g455 ( .A(n_202), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_234), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_203), .B(n_311), .Y(n_310) );
INVx4_ASAP7_75t_L g364 ( .A(n_203), .Y(n_364) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_203), .B(n_358), .Y(n_449) );
AND2x2_ASAP7_75t_L g492 ( .A(n_203), .B(n_312), .Y(n_492) );
INVx5_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g341 ( .A(n_204), .Y(n_341) );
AND2x2_ASAP7_75t_L g360 ( .A(n_204), .B(n_302), .Y(n_360) );
AND2x2_ASAP7_75t_L g378 ( .A(n_204), .B(n_312), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_204), .B(n_311), .Y(n_438) );
NOR2x1_ASAP7_75t_SL g465 ( .A(n_204), .B(n_234), .Y(n_465) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_210), .Y(n_204) );
INVx3_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_208), .Y(n_303) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_209), .B(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g236 ( .A(n_209), .B(n_233), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_219), .B(n_231), .Y(n_210) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_218), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
AND2x6_ASAP7_75t_L g229 ( .A(n_214), .B(n_222), .Y(n_229) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g227 ( .A(n_216), .B(n_224), .Y(n_227) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx5_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
AND2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx2_ASAP7_75t_L g520 ( .A(n_222), .Y(n_520) );
AND2x4_ASAP7_75t_L g517 ( .A(n_223), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g540 ( .A(n_224), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_228), .B(n_230), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_230), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_230), .A2(n_253), .B(n_254), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_265), .B(n_266), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_273), .B(n_274), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_230), .A2(n_283), .B(n_284), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_230), .A2(n_308), .B(n_309), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_230), .A2(n_316), .B(n_317), .Y(n_315) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_231), .A2(n_251), .B(n_255), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_231), .Y(n_319) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_231), .A2(n_251), .B(n_255), .Y(n_324) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_234), .B(n_302), .Y(n_301) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_237), .B(n_243), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_235), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_235), .A2(n_237), .B(n_243), .Y(n_337) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_236), .B(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_236), .A2(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_278), .B(n_287), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_247), .A2(n_347), .B1(n_351), .B2(n_352), .Y(n_346) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_256), .Y(n_247) );
AND2x2_ASAP7_75t_L g407 ( .A(n_248), .B(n_293), .Y(n_407) );
BUFx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g340 ( .A(n_249), .B(n_323), .Y(n_340) );
AND2x2_ASAP7_75t_L g412 ( .A(n_249), .B(n_295), .Y(n_412) );
AND2x2_ASAP7_75t_L g431 ( .A(n_249), .B(n_397), .Y(n_431) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_250), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_256), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g391 ( .A(n_257), .B(n_290), .Y(n_391) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_269), .Y(n_257) );
AND2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g328 ( .A(n_258), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_258), .B(n_324), .Y(n_388) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g481 ( .A(n_259), .Y(n_481) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g323 ( .A(n_260), .Y(n_323) );
OAI21x1_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_263), .B(n_267), .Y(n_260) );
INVx1_ASAP7_75t_L g268 ( .A(n_262), .Y(n_268) );
INVx2_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_269), .Y(n_429) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_276), .B(n_277), .Y(n_269) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_270), .A2(n_276), .B(n_277), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_271), .B(n_275), .Y(n_270) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_276), .A2(n_280), .B(n_286), .Y(n_279) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_280), .B(n_286), .Y(n_292) );
INVx2_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_278), .B(n_457), .Y(n_483) );
AND2x2_ASAP7_75t_L g502 ( .A(n_278), .B(n_492), .Y(n_502) );
BUFx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_279), .B(n_329), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .Y(n_280) );
AND2x2_ASAP7_75t_SL g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g369 ( .A(n_288), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_288), .B(n_339), .Y(n_374) );
INVx1_ASAP7_75t_SL g501 ( .A(n_288), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_289), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
AND2x2_ASAP7_75t_L g513 ( .A(n_290), .B(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g389 ( .A(n_291), .B(n_294), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_291), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g443 ( .A(n_291), .B(n_295), .Y(n_443) );
AND2x2_ASAP7_75t_L g474 ( .A(n_291), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g339 ( .A(n_292), .B(n_295), .Y(n_339) );
INVxp67_ASAP7_75t_L g356 ( .A(n_292), .Y(n_356) );
BUFx3_ASAP7_75t_L g397 ( .A(n_292), .Y(n_397) );
AND2x2_ASAP7_75t_L g417 ( .A(n_293), .B(n_418), .Y(n_417) );
NAND2xp33_ASAP7_75t_L g430 ( .A(n_293), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_294), .B(n_323), .Y(n_386) );
AND2x2_ASAP7_75t_L g475 ( .A(n_294), .B(n_324), .Y(n_475) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g402 ( .A(n_295), .B(n_324), .Y(n_402) );
OR3x1_ASAP7_75t_L g296 ( .A(n_297), .B(n_346), .C(n_361), .Y(n_296) );
OAI321xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_310), .A3(n_321), .B1(n_326), .B2(n_330), .C(n_338), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_301), .Y(n_377) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_301), .Y(n_395) );
OR2x2_ASAP7_75t_L g399 ( .A(n_301), .B(n_310), .Y(n_399) );
BUFx3_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
AND2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_336), .Y(n_350) );
INVx1_ASAP7_75t_L g367 ( .A(n_302), .Y(n_367) );
INVx2_ASAP7_75t_L g383 ( .A(n_302), .Y(n_383) );
OR2x2_ASAP7_75t_L g422 ( .A(n_302), .B(n_311), .Y(n_422) );
INVx2_ASAP7_75t_L g410 ( .A(n_310), .Y(n_410) );
AND2x2_ASAP7_75t_L g334 ( .A(n_311), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
AND2x4_ASAP7_75t_L g358 ( .A(n_311), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_311), .B(n_335), .Y(n_381) );
AND2x2_ASAP7_75t_L g488 ( .A(n_311), .B(n_383), .Y(n_488) );
INVx4_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_312), .Y(n_447) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B(n_320), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g375 ( .A(n_321), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_325), .Y(n_321) );
AND2x2_ASAP7_75t_L g462 ( .A(n_322), .B(n_389), .Y(n_462) );
INVx1_ASAP7_75t_SL g479 ( .A(n_322), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_322), .B(n_455), .Y(n_508) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OR2x2_ASAP7_75t_L g351 ( .A(n_323), .B(n_324), .Y(n_351) );
AND2x2_ASAP7_75t_L g444 ( .A(n_325), .B(n_340), .Y(n_444) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_329), .B(n_340), .Y(n_467) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_331), .A2(n_480), .B1(n_485), .B2(n_487), .Y(n_484) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g409 ( .A(n_332), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g504 ( .A(n_332), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g460 ( .A(n_333), .B(n_378), .Y(n_460) );
AND2x4_ASAP7_75t_L g414 ( .A(n_334), .B(n_360), .Y(n_414) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_336), .Y(n_512) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g345 ( .A(n_337), .Y(n_345) );
INVx1_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .C(n_341), .D(n_342), .Y(n_338) );
AND2x2_ASAP7_75t_L g496 ( .A(n_339), .B(n_481), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_339), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_340), .B(n_416), .Y(n_415) );
OAI322xp33_ASAP7_75t_L g423 ( .A1(n_340), .A2(n_424), .A3(n_428), .B1(n_430), .B2(n_432), .C1(n_434), .C2(n_439), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_340), .B(n_389), .Y(n_439) );
INVx1_ASAP7_75t_L g507 ( .A(n_340), .Y(n_507) );
INVx2_ASAP7_75t_L g353 ( .A(n_341), .Y(n_353) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_344), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_345), .B(n_364), .Y(n_421) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_348), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
AND2x2_ASAP7_75t_L g466 ( .A(n_349), .B(n_377), .Y(n_466) );
AOI31xp33_ASAP7_75t_L g352 ( .A1(n_350), .A2(n_353), .A3(n_354), .B(n_357), .Y(n_352) );
AND2x2_ASAP7_75t_L g363 ( .A(n_350), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g491 ( .A(n_350), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_350), .B(n_378), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_350), .Y(n_499) );
INVx1_ASAP7_75t_SL g457 ( .A(n_351), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_351), .B(n_479), .C(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_358), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g427 ( .A(n_358), .Y(n_427) );
AOI322xp5_ASAP7_75t_L g509 ( .A1(n_358), .A2(n_388), .A3(n_391), .B1(n_510), .B2(n_511), .C1(n_513), .C2(n_515), .Y(n_509) );
AND2x2_ASAP7_75t_L g515 ( .A(n_358), .B(n_364), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_368), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_364), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g510 ( .A(n_364), .B(n_397), .Y(n_510) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
AND2x2_ASAP7_75t_L g464 ( .A(n_367), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g511 ( .A(n_367), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_376), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g433 ( .A(n_378), .B(n_383), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B(n_390), .C(n_392), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_380), .A2(n_406), .B1(n_408), .B2(n_411), .C(n_413), .Y(n_405) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
OR2x2_ASAP7_75t_L g445 ( .A(n_382), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g490 ( .A(n_385), .Y(n_490) );
INVx1_ASAP7_75t_L g514 ( .A(n_386), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AND2x2_ASAP7_75t_L g396 ( .A(n_388), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_388), .B(n_458), .Y(n_470) );
INVx1_ASAP7_75t_L g450 ( .A(n_389), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_398), .B2(n_400), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_SL g458 ( .A(n_397), .Y(n_458) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND4xp75_ASAP7_75t_L g403 ( .A(n_404), .B(n_440), .C(n_468), .D(n_493), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_405), .B(n_423), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_412), .B(n_481), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_417), .B2(n_419), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_416), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
OR2x2_ASAP7_75t_L g471 ( .A(n_422), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g477 ( .A1(n_433), .A2(n_478), .B(n_480), .Y(n_477) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_453), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_448), .B2(n_450), .C(n_451), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_443), .A2(n_490), .B(n_491), .Y(n_489) );
INVx3_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
OAI322xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .A3(n_458), .B1(n_459), .B2(n_461), .C1(n_463), .C2(n_467), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g476 ( .A(n_464), .Y(n_476) );
INVx1_ASAP7_75t_L g472 ( .A(n_465), .Y(n_472) );
AND2x2_ASAP7_75t_L g487 ( .A(n_465), .B(n_488), .Y(n_487) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_482), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_473), .B2(n_476), .C(n_477), .Y(n_469) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
OAI211xp5_ASAP7_75t_SL g482 ( .A1(n_476), .A2(n_483), .B(n_484), .C(n_489), .Y(n_482) );
INVx2_ASAP7_75t_SL g505 ( .A(n_492), .Y(n_505) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B1(n_499), .B2(n_500), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
OAI211xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_508), .C(n_509), .Y(n_503) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_518), .Y(n_537) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI222xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B1(n_530), .B2(n_532), .C1(n_535), .C2(n_541), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
endmodule