module real_aes_18144_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g102 ( .A(n_0), .B(n_103), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_1), .A2(n_4), .B1(n_242), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_2), .A2(n_40), .B1(n_137), .B2(n_139), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_3), .A2(n_22), .B1(n_139), .B2(n_182), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_5), .A2(n_15), .B1(n_164), .B2(n_233), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_6), .A2(n_57), .B1(n_184), .B2(n_209), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_7), .A2(n_16), .B1(n_137), .B2(n_168), .Y(n_599) );
INVx1_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_9), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_10), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_11), .A2(n_17), .B1(n_166), .B2(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g110 ( .A(n_12), .B(n_36), .Y(n_110) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_14), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_18), .A2(n_96), .B1(n_164), .B2(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_19), .A2(n_37), .B1(n_200), .B2(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_20), .B(n_165), .Y(n_197) );
OAI21x1_ASAP7_75t_L g153 ( .A1(n_21), .A2(n_54), .B(n_154), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_23), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_24), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_25), .B(n_143), .Y(n_507) );
INVx4_ASAP7_75t_R g562 ( .A(n_26), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_27), .A2(n_44), .B1(n_145), .B2(n_147), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_28), .A2(n_50), .B1(n_147), .B2(n_164), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_29), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_30), .B(n_200), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_31), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_32), .B(n_139), .Y(n_514) );
INVx1_ASAP7_75t_L g523 ( .A(n_33), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_SL g580 ( .A1(n_34), .A2(n_137), .B(n_149), .C(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_35), .A2(n_51), .B1(n_137), .B2(n_147), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_38), .A2(n_82), .B1(n_137), .B2(n_181), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_39), .A2(n_43), .B1(n_137), .B2(n_168), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_41), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_42), .A2(n_56), .B1(n_164), .B2(n_219), .Y(n_244) );
INVx1_ASAP7_75t_L g511 ( .A(n_45), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_46), .B(n_137), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_47), .Y(n_532) );
INVx2_ASAP7_75t_L g116 ( .A(n_48), .Y(n_116) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
BUFx3_ASAP7_75t_L g119 ( .A(n_49), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_52), .A2(n_121), .B1(n_828), .B2(n_829), .Y(n_120) );
INVx1_ASAP7_75t_L g828 ( .A(n_52), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_53), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_55), .A2(n_84), .B1(n_137), .B2(n_147), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_58), .A2(n_71), .B1(n_145), .B2(n_219), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_59), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_60), .A2(n_73), .B1(n_137), .B2(n_168), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_61), .A2(n_94), .B1(n_164), .B2(n_166), .Y(n_163) );
AND2x4_ASAP7_75t_L g133 ( .A(n_62), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g154 ( .A(n_63), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_64), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_65), .A2(n_87), .B1(n_145), .B2(n_147), .Y(n_519) );
AO22x1_ASAP7_75t_L g549 ( .A1(n_66), .A2(n_72), .B1(n_230), .B2(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g134 ( .A(n_67), .Y(n_134) );
AND2x2_ASAP7_75t_L g583 ( .A(n_68), .B(n_151), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_69), .B(n_184), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_70), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_74), .B(n_139), .Y(n_533) );
INVx2_ASAP7_75t_L g143 ( .A(n_75), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_76), .B(n_151), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_77), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_78), .A2(n_95), .B1(n_147), .B2(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_79), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_80), .B(n_161), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_81), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_83), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_85), .A2(n_122), .B1(n_840), .B2(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_85), .Y(n_840) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_86), .B(n_151), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_88), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_89), .B(n_151), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_90), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g482 ( .A(n_90), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g201 ( .A(n_91), .B(n_165), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_92), .A2(n_170), .B(n_184), .C(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g564 ( .A(n_93), .B(n_565), .Y(n_564) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_97), .B(n_146), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_111), .B(n_855), .Y(n_98) );
CKINVDCx6p67_ASAP7_75t_R g99 ( .A(n_100), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx2_ASAP7_75t_SL g865 ( .A(n_102), .Y(n_865) );
INVx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx3_ASAP7_75t_L g866 ( .A(n_105), .Y(n_866) );
AND2x6_ASAP7_75t_SL g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_108), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_109), .B(n_118), .Y(n_117) );
AND3x2_ASAP7_75t_L g836 ( .A(n_109), .B(n_837), .C(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_110), .B(n_119), .Y(n_854) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_120), .B(n_830), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x6_ASAP7_75t_SL g114 ( .A(n_115), .B(n_117), .Y(n_114) );
BUFx3_ASAP7_75t_L g846 ( .A(n_115), .Y(n_846) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_116), .B(n_852), .Y(n_851) );
INVx3_ASAP7_75t_L g863 ( .A(n_116), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_116), .B(n_866), .Y(n_870) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g829 ( .A(n_121), .Y(n_829) );
OA22x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_478), .B1(n_483), .B2(n_485), .Y(n_121) );
INVx2_ASAP7_75t_L g841 ( .A(n_122), .Y(n_841) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_374), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_326), .Y(n_123) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_273), .C(n_311), .Y(n_124) );
AOI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_204), .B1(n_224), .B2(n_252), .C(n_258), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_126), .A2(n_451), .B1(n_454), .B2(n_455), .Y(n_450) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_175), .Y(n_127) );
INVx1_ASAP7_75t_L g365 ( .A(n_128), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_157), .Y(n_128) );
INVx1_ASAP7_75t_L g317 ( .A(n_129), .Y(n_317) );
AND2x4_ASAP7_75t_L g360 ( .A(n_129), .B(n_281), .Y(n_360) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g288 ( .A(n_130), .B(n_191), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_130), .B(n_257), .Y(n_348) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g256 ( .A(n_131), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g272 ( .A(n_131), .B(n_177), .Y(n_272) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_131), .Y(n_279) );
INVx1_ASAP7_75t_L g335 ( .A(n_131), .Y(n_335) );
AO31x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_135), .A3(n_150), .B(n_155), .Y(n_131) );
INVx2_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_132), .A2(n_159), .A3(n_206), .B(n_212), .Y(n_205) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_132), .A2(n_178), .A3(n_228), .B(n_235), .Y(n_227) );
AO31x2_ASAP7_75t_L g597 ( .A1(n_132), .A2(n_223), .A3(n_598), .B(n_601), .Y(n_597) );
BUFx10_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
BUFx10_ASAP7_75t_L g498 ( .A(n_133), .Y(n_498) );
INVx1_ASAP7_75t_L g553 ( .A(n_133), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B1(n_144), .B2(n_148), .Y(n_135) );
INVx1_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
INVx4_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g219 ( .A(n_137), .Y(n_219) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_138), .Y(n_139) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
INVx2_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
INVx1_ASAP7_75t_L g231 ( .A(n_138), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx1_ASAP7_75t_L g243 ( .A(n_138), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_139), .B(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_140), .A2(n_148), .B1(n_218), .B2(n_220), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_140), .A2(n_148), .B1(n_229), .B2(n_232), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_140), .A2(n_148), .B1(n_241), .B2(n_244), .Y(n_240) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g497 ( .A(n_141), .Y(n_497) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g535 ( .A(n_142), .Y(n_535) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx8_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
INVx1_ASAP7_75t_L g510 ( .A(n_143), .Y(n_510) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_146), .A2(n_234), .B1(n_562), .B2(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_147), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g521 ( .A(n_147), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_148), .A2(n_163), .B1(n_167), .B2(n_169), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_148), .A2(n_180), .B1(n_183), .B2(n_185), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_148), .A2(n_199), .B(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_148), .A2(n_169), .B1(n_207), .B2(n_211), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_148), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_148), .A2(n_185), .B1(n_519), .B2(n_520), .Y(n_518) );
OAI22x1_ASAP7_75t_L g598 ( .A1(n_148), .A2(n_185), .B1(n_599), .B2(n_600), .Y(n_598) );
INVx6_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_168), .B(n_196), .C(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_149), .A2(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_149), .B(n_549), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_149), .A2(n_545), .B(n_549), .C(n_552), .Y(n_611) );
AO31x2_ASAP7_75t_L g493 ( .A1(n_150), .A2(n_494), .A3(n_498), .B(n_499), .Y(n_493) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_151), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_152), .B(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_152), .B(n_174), .Y(n_173) );
BUFx3_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx2_ASAP7_75t_SL g193 ( .A(n_152), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_152), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g515 ( .A(n_152), .B(n_498), .Y(n_515) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
INVx3_ASAP7_75t_L g255 ( .A(n_157), .Y(n_255) );
AND2x2_ASAP7_75t_L g270 ( .A(n_157), .B(n_191), .Y(n_270) );
INVx2_ASAP7_75t_L g276 ( .A(n_157), .Y(n_276) );
AND2x4_ASAP7_75t_L g338 ( .A(n_157), .B(n_177), .Y(n_338) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_157), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_157), .B(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g287 ( .A(n_158), .B(n_177), .Y(n_287) );
AND2x2_ASAP7_75t_L g315 ( .A(n_158), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g394 ( .A(n_158), .Y(n_394) );
AO31x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .A3(n_171), .B(n_173), .Y(n_158) );
AO31x2_ASAP7_75t_L g517 ( .A1(n_159), .A2(n_186), .A3(n_518), .B(n_522), .Y(n_517) );
AOI21x1_ASAP7_75t_L g572 ( .A1(n_159), .A2(n_573), .B(n_583), .Y(n_572) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_160), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_160), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g565 ( .A(n_160), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_160), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
INVx2_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_161), .A2(n_547), .B(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_165), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_168), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_171), .A2(n_215), .A3(n_240), .B(n_245), .Y(n_239) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_172), .A2(n_557), .B(n_560), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
INVx1_ASAP7_75t_L g350 ( .A(n_176), .Y(n_350) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_176), .B(n_270), .Y(n_378) );
BUFx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x2_ASAP7_75t_L g280 ( .A(n_177), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g316 ( .A(n_177), .Y(n_316) );
INVx1_ASAP7_75t_L g392 ( .A(n_177), .Y(n_392) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .A3(n_186), .B(n_188), .Y(n_177) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_182), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_185), .B(n_561), .Y(n_560) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_186), .A2(n_215), .A3(n_217), .B(n_221), .Y(n_214) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_SL g202 ( .A(n_187), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_189), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
AND2x4_ASAP7_75t_L g331 ( .A(n_191), .B(n_316), .Y(n_331) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g353 ( .A(n_192), .Y(n_353) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_203), .Y(n_192) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_193), .A2(n_194), .B(n_203), .Y(n_257) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_198), .B(n_202), .Y(n_194) );
AND2x4_ASAP7_75t_L g225 ( .A(n_204), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
INVx4_ASAP7_75t_SL g249 ( .A(n_205), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_205), .B(n_251), .Y(n_261) );
BUFx2_ASAP7_75t_L g325 ( .A(n_205), .Y(n_325) );
AND2x2_ASAP7_75t_L g369 ( .A(n_205), .B(n_227), .Y(n_369) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_210), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g247 ( .A(n_214), .Y(n_247) );
OR2x2_ASAP7_75t_L g285 ( .A(n_214), .B(n_227), .Y(n_285) );
INVx2_ASAP7_75t_L g296 ( .A(n_214), .Y(n_296) );
AND2x4_ASAP7_75t_L g299 ( .A(n_214), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_214), .Y(n_340) );
INVx1_ASAP7_75t_L g381 ( .A(n_214), .Y(n_381) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_215), .A2(n_556), .B(n_564), .Y(n_555) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_223), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_237), .Y(n_224) );
INVx2_ASAP7_75t_L g474 ( .A(n_225), .Y(n_474) );
AND2x4_ASAP7_75t_L g435 ( .A(n_226), .B(n_238), .Y(n_435) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g251 ( .A(n_227), .Y(n_251) );
INVx2_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
INVx1_ASAP7_75t_L g356 ( .A(n_227), .Y(n_356) );
AND2x2_ASAP7_75t_L g382 ( .A(n_227), .B(n_307), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_227), .B(n_295), .Y(n_386) );
OAI21xp33_ASAP7_75t_SL g506 ( .A1(n_230), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_248), .Y(n_237) );
INVx3_ASAP7_75t_L g363 ( .A(n_238), .Y(n_363) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_247), .Y(n_238) );
INVx2_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
INVx2_ASAP7_75t_L g307 ( .A(n_239), .Y(n_307) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_243), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_247), .B(n_249), .Y(n_308) );
AND2x2_ASAP7_75t_L g336 ( .A(n_247), .B(n_307), .Y(n_336) );
INVx1_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_248), .B(n_372), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_248), .B(n_336), .Y(n_447) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g265 ( .A(n_249), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_249), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g355 ( .A(n_249), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_249), .Y(n_432) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_252), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_254), .B(n_288), .Y(n_323) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g346 ( .A(n_255), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g445 ( .A(n_255), .B(n_256), .Y(n_445) );
AND2x2_ASAP7_75t_L g318 ( .A(n_256), .B(n_287), .Y(n_318) );
AND2x4_ASAP7_75t_L g337 ( .A(n_256), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g388 ( .A(n_256), .B(n_315), .Y(n_388) );
INVx1_ASAP7_75t_L g281 ( .A(n_257), .Y(n_281) );
AOI31xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .A3(n_263), .B(n_268), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_260), .B(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_260), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_260), .A2(n_262), .B(n_292), .Y(n_472) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g449 ( .A(n_264), .B(n_285), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_266), .Y(n_411) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
OR2x2_ASAP7_75t_L g321 ( .A(n_267), .B(n_296), .Y(n_321) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2x1p5_ASAP7_75t_L g310 ( .A(n_272), .B(n_276), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_282), .B1(n_286), .B2(n_289), .C(n_301), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g390 ( .A(n_279), .B(n_293), .Y(n_390) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OR2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g407 ( .A(n_283), .B(n_299), .Y(n_407) );
AND2x4_ASAP7_75t_L g324 ( .A(n_284), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g343 ( .A(n_285), .B(n_306), .Y(n_343) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x4_ASAP7_75t_SL g359 ( .A(n_287), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g400 ( .A(n_287), .Y(n_400) );
INVx2_ASAP7_75t_L g409 ( .A(n_287), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_287), .B(n_353), .Y(n_423) );
INVx1_ASAP7_75t_L g401 ( .A(n_288), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_297), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_291), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_292), .B(n_299), .Y(n_333) );
AND2x2_ASAP7_75t_L g354 ( .A(n_292), .B(n_355), .Y(n_354) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_292), .B(n_324), .Y(n_462) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B(n_309), .Y(n_301) );
NAND2x1_ASAP7_75t_L g463 ( .A(n_303), .B(n_407), .Y(n_463) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_304), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx4_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
AND2x2_ASAP7_75t_L g442 ( .A(n_306), .B(n_347), .Y(n_442) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g339 ( .A(n_307), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_353), .Y(n_352) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_310), .B(n_423), .Y(n_422) );
AOI322xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .A3(n_317), .B1(n_318), .B2(n_319), .C1(n_322), .C2(n_324), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g405 ( .A(n_315), .B(n_353), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_315), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g429 ( .A(n_315), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g434 ( .A(n_315), .B(n_419), .Y(n_434) );
INVx1_ASAP7_75t_L g443 ( .A(n_315), .Y(n_443) );
OR2x2_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g456 ( .A(n_317), .Y(n_456) );
AND2x2_ASAP7_75t_L g459 ( .A(n_318), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_321), .B(n_335), .C(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g437 ( .A(n_321), .Y(n_437) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND3xp33_ASAP7_75t_SL g326 ( .A(n_327), .B(n_341), .C(n_351), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_332), .B1(n_334), .B2(n_336), .C1(n_337), .C2(n_339), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22x1_ASAP7_75t_L g473 ( .A1(n_330), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g334 ( .A(n_331), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_331), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g427 ( .A(n_331), .B(n_393), .Y(n_427) );
AND2x4_ASAP7_75t_L g457 ( .A(n_331), .B(n_394), .Y(n_457) );
AND2x2_ASAP7_75t_L g438 ( .A(n_332), .B(n_405), .Y(n_438) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g430 ( .A(n_335), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_336), .B(n_369), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_336), .B(n_355), .Y(n_453) );
INVx1_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
INVx2_ASAP7_75t_L g417 ( .A(n_339), .Y(n_417) );
INVx1_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AOI221xp5_ASAP7_75t_SL g433 ( .A1(n_346), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_433) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g419 ( .A(n_348), .Y(n_419) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_348), .Y(n_471) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_350), .B(n_456), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_357), .B2(n_368), .C(n_370), .Y(n_351) );
OR2x2_ASAP7_75t_L g408 ( .A(n_353), .B(n_409), .Y(n_408) );
AOI32xp33_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_369), .A3(n_390), .B1(n_391), .B2(n_395), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_355), .B(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B1(n_364), .B2(n_366), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_360), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g431 ( .A(n_363), .B(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g424 ( .A(n_367), .B(n_369), .Y(n_424) );
AND2x2_ASAP7_75t_L g477 ( .A(n_367), .B(n_382), .Y(n_477) );
AND2x2_ASAP7_75t_L g436 ( .A(n_368), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_369), .B(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_375), .B(n_439), .Y(n_374) );
NAND4xp75_ASAP7_75t_L g375 ( .A(n_376), .B(n_402), .C(n_420), .D(n_433), .Y(n_375) );
AOI211x1_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_383), .C(n_397), .Y(n_376) );
INVxp67_ASAP7_75t_L g475 ( .A(n_377), .Y(n_475) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
BUFx2_ASAP7_75t_L g396 ( .A(n_392), .Y(n_396) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g468 ( .A(n_396), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .C(n_401), .Y(n_397) );
INVx2_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_412), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_408), .B2(n_410), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_417), .B2(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B(n_425), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_432), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g452 ( .A(n_435), .Y(n_452) );
NAND4xp75_ASAP7_75t_SL g439 ( .A(n_440), .B(n_450), .C(n_458), .D(n_466), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NOR2xp67_ASAP7_75t_SL g458 ( .A(n_459), .B(n_461), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_464), .Y(n_461) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AOI21x1_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_472), .B(n_473), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx8_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx12f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
BUFx8_ASAP7_75t_SL g484 ( .A(n_481), .Y(n_484) );
AND2x2_ASAP7_75t_L g853 ( .A(n_481), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g838 ( .A(n_482), .Y(n_838) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_718), .Y(n_485) );
NOR4xp25_ASAP7_75t_L g486 ( .A(n_487), .B(n_618), .C(n_660), .D(n_692), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_524), .B(n_566), .C(n_603), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
INVx2_ASAP7_75t_L g631 ( .A(n_491), .Y(n_631) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g710 ( .A(n_492), .B(n_503), .Y(n_710) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_493), .B(n_517), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_493), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g617 ( .A(n_493), .Y(n_617) );
OR2x2_ASAP7_75t_L g680 ( .A(n_493), .B(n_517), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_497), .A2(n_513), .B(n_514), .Y(n_512) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_497), .A2(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g614 ( .A(n_502), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g626 ( .A(n_502), .Y(n_626) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_502), .Y(n_804) );
OR2x2_ASAP7_75t_L g817 ( .A(n_502), .B(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_516), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_503), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g590 ( .A(n_503), .Y(n_590) );
AND2x2_ASAP7_75t_L g637 ( .A(n_503), .B(n_638), .Y(n_637) );
NAND2x1p5_ASAP7_75t_SL g656 ( .A(n_503), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_503), .B(n_591), .Y(n_706) );
INVx1_ASAP7_75t_L g795 ( .A(n_503), .Y(n_795) );
AND2x2_ASAP7_75t_L g824 ( .A(n_503), .B(n_517), .Y(n_824) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_512), .B(n_515), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_517), .B(n_617), .Y(n_639) );
INVx1_ASAP7_75t_L g659 ( .A(n_517), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_517), .B(n_593), .Y(n_711) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_541), .Y(n_525) );
OR2x2_ASAP7_75t_L g608 ( .A(n_526), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g715 ( .A(n_526), .B(n_664), .Y(n_715) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g624 ( .A(n_527), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_527), .B(n_644), .Y(n_643) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_527), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g587 ( .A(n_528), .Y(n_587) );
BUFx3_ASAP7_75t_L g635 ( .A(n_528), .Y(n_635) );
AND2x2_ASAP7_75t_L g671 ( .A(n_528), .B(n_652), .Y(n_671) );
AND2x2_ASAP7_75t_L g751 ( .A(n_528), .B(n_597), .Y(n_751) );
AND2x2_ASAP7_75t_L g764 ( .A(n_528), .B(n_555), .Y(n_764) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_536), .B(n_539), .Y(n_530) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g704 ( .A(n_541), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_541), .B(n_634), .Y(n_712) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_554), .Y(n_541) );
AND2x2_ASAP7_75t_L g623 ( .A(n_542), .B(n_555), .Y(n_623) );
INVx1_ASAP7_75t_L g731 ( .A(n_542), .Y(n_731) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g585 ( .A(n_543), .B(n_555), .Y(n_585) );
AND2x2_ASAP7_75t_L g648 ( .A(n_543), .B(n_554), .Y(n_648) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_548), .B(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_553), .A2(n_574), .B(n_580), .Y(n_573) );
AND2x2_ASAP7_75t_L g606 ( .A(n_554), .B(n_597), .Y(n_606) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g664 ( .A(n_555), .B(n_597), .Y(n_664) );
INVx1_ASAP7_75t_L g675 ( .A(n_555), .Y(n_675) );
AND2x2_ASAP7_75t_L g738 ( .A(n_555), .B(n_587), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_584), .B1(n_588), .B2(n_594), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_567), .A2(n_637), .B1(n_640), .B2(n_642), .Y(n_636) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
OR2x2_ASAP7_75t_L g716 ( .A(n_569), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g822 ( .A(n_569), .Y(n_822) );
INVx1_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
OR2x2_ASAP7_75t_L g744 ( .A(n_570), .B(n_639), .Y(n_744) );
OR2x2_ASAP7_75t_L g615 ( .A(n_571), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_571), .B(n_590), .Y(n_691) );
AND2x2_ASAP7_75t_L g708 ( .A(n_571), .B(n_635), .Y(n_708) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_571), .Y(n_725) );
INVxp67_ASAP7_75t_L g773 ( .A(n_571), .Y(n_773) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g593 ( .A(n_572), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B(n_579), .Y(n_574) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_585), .Y(n_683) );
INVx3_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
AND2x2_ASAP7_75t_L g701 ( .A(n_585), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g801 ( .A(n_585), .B(n_763), .Y(n_801) );
INVx1_ASAP7_75t_L g595 ( .A(n_586), .Y(n_595) );
OR2x2_ASAP7_75t_L g778 ( .A(n_586), .B(n_753), .Y(n_778) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g702 ( .A(n_587), .B(n_612), .Y(n_702) );
AND2x2_ASAP7_75t_L g723 ( .A(n_587), .B(n_648), .Y(n_723) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_589), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g724 ( .A(n_589), .Y(n_724) );
AND2x2_ASAP7_75t_L g766 ( .A(n_589), .B(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g667 ( .A(n_590), .Y(n_667) );
AND2x2_ASAP7_75t_L g698 ( .A(n_590), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_590), .B(n_657), .Y(n_717) );
AND2x2_ASAP7_75t_L g666 ( .A(n_592), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g782 ( .A(n_592), .Y(n_782) );
AND2x2_ASAP7_75t_L g805 ( .A(n_592), .B(n_795), .Y(n_805) );
INVx1_ASAP7_75t_L g818 ( .A(n_592), .Y(n_818) );
INVx2_ASAP7_75t_L g657 ( .A(n_593), .Y(n_657) );
OR2x2_ASAP7_75t_L g753 ( .A(n_593), .B(n_617), .Y(n_753) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_596), .B(n_634), .Y(n_641) );
INVx2_ASAP7_75t_L g612 ( .A(n_597), .Y(n_612) );
INVx2_ASAP7_75t_L g652 ( .A(n_597), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_597), .B(n_610), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_613), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_606), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g747 ( .A(n_609), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx2_ASAP7_75t_L g653 ( .A(n_610), .Y(n_653) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g627 ( .A(n_615), .Y(n_627) );
INVxp67_ASAP7_75t_L g798 ( .A(n_615), .Y(n_798) );
OR2x2_ASAP7_75t_L g700 ( .A(n_616), .B(n_657), .Y(n_700) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_628), .C(n_636), .D(n_645), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_625), .C(n_627), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_621), .A2(n_815), .B(n_817), .C(n_819), .Y(n_814) );
OR2x6_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_623), .B(n_671), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_623), .B(n_727), .C(n_729), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_623), .B(n_702), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_623), .A2(n_728), .B1(n_820), .B2(n_823), .C(n_825), .Y(n_819) );
INVx1_ASAP7_75t_L g810 ( .A(n_624), .Y(n_810) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_629), .A2(n_637), .B1(n_672), .B2(n_746), .C(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_631), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g696 ( .A(n_632), .Y(n_696) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_634), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g811 ( .A(n_634), .B(n_662), .Y(n_811) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g647 ( .A(n_635), .Y(n_647) );
AND3x1_ASAP7_75t_L g820 ( .A(n_635), .B(n_821), .C(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g690 ( .A(n_639), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g760 ( .A(n_642), .Y(n_760) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g736 ( .A(n_644), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g763 ( .A(n_644), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B(n_654), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_647), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g728 ( .A(n_648), .Y(n_728) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g684 ( .A(n_652), .Y(n_684) );
OR2x2_ASAP7_75t_L g663 ( .A(n_653), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g776 ( .A(n_653), .Y(n_776) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_655), .B(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
OR2x2_ASAP7_75t_L g732 ( .A(n_656), .B(n_680), .Y(n_732) );
INVx2_ASAP7_75t_L g821 ( .A(n_656), .Y(n_821) );
INVx1_ASAP7_75t_L g695 ( .A(n_657), .Y(n_695) );
NOR4xp25_ASAP7_75t_L g825 ( .A(n_657), .B(n_688), .C(n_826), .D(n_827), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_658), .Y(n_827) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx3_ASAP7_75t_L g813 ( .A(n_659), .Y(n_813) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_665), .B(n_668), .C(n_676), .Y(n_660) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g800 ( .A(n_663), .Y(n_800) );
INVx2_ASAP7_75t_L g785 ( .A(n_664), .Y(n_785) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_666), .A2(n_669), .B(n_672), .Y(n_668) );
OR2x2_ASAP7_75t_L g752 ( .A(n_667), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g770 ( .A(n_667), .B(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g686 ( .A(n_671), .Y(n_686) );
AND2x4_ASAP7_75t_SL g775 ( .A(n_671), .B(n_776), .Y(n_775) );
INVx3_ASAP7_75t_R g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_674), .Y(n_741) );
INVx1_ASAP7_75t_L g748 ( .A(n_675), .Y(n_748) );
AOI32xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_682), .A3(n_684), .B1(n_685), .B2(n_689), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_679), .B(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_679), .Y(n_740) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g757 ( .A(n_680), .B(n_695), .Y(n_757) );
INVx2_ASAP7_75t_L g771 ( .A(n_680), .Y(n_771) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_688), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .B(n_697), .C(n_713), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B(n_703), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g754 ( .A(n_702), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_702), .B(n_789), .Y(n_788) );
OAI32xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .A3(n_707), .B1(n_709), .B2(n_712), .Y(n_703) );
INVx1_ASAP7_75t_L g789 ( .A(n_704), .Y(n_789) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g781 ( .A(n_706), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_790), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_745), .C(n_758), .D(n_786), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g720 ( .A(n_721), .B(n_733), .Y(n_720) );
OAI32xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .A3(n_725), .B1(n_726), .B2(n_732), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g772 ( .A(n_724), .B(n_773), .Y(n_772) );
OAI32xp33_ASAP7_75t_L g777 ( .A1(n_724), .A2(n_778), .A3(n_779), .B1(n_781), .B2(n_783), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_725), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_727), .B(n_792), .Y(n_791) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g784 ( .A(n_730), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g816 ( .A(n_730), .Y(n_816) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g780 ( .A(n_731), .Y(n_780) );
OAI22x1_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_739), .B1(n_741), .B2(n_742), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_743), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2x1_ASAP7_75t_L g809 ( .A(n_747), .B(n_810), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_754), .B2(n_755), .Y(n_749) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_751), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g826 ( .A(n_751), .Y(n_826) );
INVx2_ASAP7_75t_L g767 ( .A(n_753), .Y(n_767) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR3xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_768), .C(n_777), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B(n_765), .Y(n_759) );
NAND2xp33_ASAP7_75t_L g787 ( .A(n_761), .B(n_788), .Y(n_787) );
INVx2_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x4_ASAP7_75t_L g823 ( .A(n_767), .B(n_824), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_772), .B(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x4_ASAP7_75t_L g794 ( .A(n_771), .B(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_773), .Y(n_793) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND3xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_796), .C(n_808), .Y(n_790) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx1_ASAP7_75t_L g799 ( .A(n_795), .Y(n_799) );
AOI222xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_800), .B1(n_801), .B2(n_802), .C1(n_805), .C2(n_806), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
O2A1O1Ixp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_811), .B(n_812), .C(n_814), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_845), .B(n_847), .Y(n_830) );
INVxp67_ASAP7_75t_L g867 ( .A(n_831), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_839), .B(n_842), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx3_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2x1_ASAP7_75t_R g843 ( .A(n_835), .B(n_844), .Y(n_843) );
INVx4_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_840), .A2(n_856), .B1(n_867), .B2(n_868), .Y(n_855) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
INVx6_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx10_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
OR2x6_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
OR2x4_ASAP7_75t_L g869 ( .A(n_864), .B(n_870), .Y(n_869) );
BUFx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx4_ASAP7_75t_SL g868 ( .A(n_869), .Y(n_868) );
endmodule