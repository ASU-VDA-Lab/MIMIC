module fake_jpeg_3072_n_191 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_55),
.B1(n_61),
.B2(n_63),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_62),
.B(n_44),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_63),
.B1(n_61),
.B2(n_47),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_60),
.B(n_57),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_47),
.B(n_45),
.C(n_54),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_49),
.B1(n_51),
.B2(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_67),
.B1(n_62),
.B2(n_56),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_82),
.B1(n_73),
.B2(n_53),
.Y(n_105)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_120),
.B1(n_99),
.B2(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_112),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_49),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_1),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_2),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_2),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_112),
.B(n_103),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_3),
.B(n_6),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_126),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_132),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_86),
.B1(n_90),
.B2(n_95),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_117),
.A3(n_110),
.B1(n_21),
.B2(n_23),
.C(n_42),
.Y(n_141)
);

OAI321xp33_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_15),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_117),
.CON(n_143),
.SN(n_143)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_149),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_41),
.B(n_40),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_131),
.CI(n_125),
.CON(n_150),
.SN(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_156),
.B(n_128),
.C(n_121),
.D(n_32),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_6),
.B(n_7),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_8),
.B(n_9),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_156),
.B1(n_151),
.B2(n_152),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_39),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_138),
.B1(n_128),
.B2(n_121),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_170),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_26),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_155),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_153),
.B1(n_148),
.B2(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_175),
.B(n_176),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_146),
.C(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_24),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_163),
.A3(n_150),
.B1(n_159),
.B2(n_165),
.C(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_180),
.B1(n_18),
.B2(n_15),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_174),
.B(n_13),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_177),
.B1(n_175),
.B2(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_187),
.B(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_11),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_16),
.B(n_17),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_18),
.Y(n_191)
);


endmodule