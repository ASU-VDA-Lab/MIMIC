module fake_jpeg_1715_n_199 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_9),
.B(n_27),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_0),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_58),
.B1(n_55),
.B2(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_58),
.B1(n_64),
.B2(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_46),
.B1(n_61),
.B2(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_46),
.B1(n_61),
.B2(n_51),
.Y(n_80)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_93),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_58),
.B1(n_74),
.B2(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_77),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_94),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_68),
.C(n_71),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_80),
.B1(n_65),
.B2(n_72),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_72),
.B1(n_65),
.B2(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_47),
.B2(n_53),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_55),
.B1(n_52),
.B2(n_62),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_0),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_75),
.B1(n_76),
.B2(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_114),
.B1(n_119),
.B2(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_118),
.B(n_7),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_49),
.B1(n_63),
.B2(n_45),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_63),
.B(n_50),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_57),
.B1(n_50),
.B2(n_45),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_132),
.C(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_126),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_53),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_54),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_139),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_54),
.B1(n_2),
.B2(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_134),
.B1(n_137),
.B2(n_13),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_54),
.B(n_4),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_138),
.B(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_42),
.C(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_12),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_5),
.Y(n_136)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_39),
.B(n_38),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_5),
.B(n_6),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_6),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_12),
.B(n_13),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_140),
.Y(n_160)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_37),
.C(n_36),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_132),
.C(n_130),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_126),
.B(n_138),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_137),
.B1(n_18),
.B2(n_19),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_137),
.C(n_35),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_137),
.C(n_34),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_173),
.B1(n_156),
.B2(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_179),
.B1(n_163),
.B2(n_170),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_144),
.A3(n_148),
.B1(n_155),
.B2(n_158),
.C1(n_152),
.C2(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_152),
.A3(n_154),
.B1(n_159),
.B2(n_145),
.C1(n_22),
.C2(n_26),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_23),
.A3(n_24),
.B1(n_26),
.B2(n_30),
.C(n_31),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_169),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_166),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_178),
.C(n_181),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_183),
.B(n_174),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_189),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_173),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_33),
.Y(n_199)
);


endmodule