module fake_jpeg_2958_n_114 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_26),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_20),
.Y(n_24)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_20),
.B1(n_18),
.B2(n_13),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_25),
.B1(n_27),
.B2(n_17),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_18),
.C(n_16),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_42),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_21),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_33),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_15),
.B1(n_17),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_51),
.B1(n_21),
.B2(n_38),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_39),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_61),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_39),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_49),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_37),
.C(n_33),
.Y(n_81)
);

XOR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_53),
.C(n_46),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_16),
.A3(n_14),
.B1(n_48),
.B2(n_44),
.C1(n_33),
.C2(n_37),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_72),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_61),
.B1(n_58),
.B2(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_82),
.B1(n_79),
.B2(n_70),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_79),
.B(n_81),
.Y(n_86)
);

AOI21x1_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_44),
.B(n_48),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_35),
.B1(n_31),
.B2(n_16),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_65),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_93),
.C(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_35),
.B1(n_31),
.B2(n_14),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_66),
.C(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_92),
.B1(n_90),
.B2(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.C(n_98),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_89),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_14),
.C(n_4),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_14),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_1),
.C(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_92),
.B(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_96),
.B1(n_4),
.B2(n_6),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_6),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_10),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_107),
.B(n_105),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_111),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_3),
.B1(n_106),
.B2(n_112),
.C(n_111),
.Y(n_114)
);


endmodule