module fake_jpeg_21677_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_7),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_4),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_38)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_39),
.A3(n_49),
.B1(n_26),
.B2(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_15),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_35),
.B1(n_26),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_54),
.Y(n_85)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_32),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_73),
.B(n_12),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_37),
.C(n_27),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_69),
.C(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_70),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_14),
.B1(n_34),
.B2(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_5),
.Y(n_68)
);

NOR2xp67_ASAP7_75t_R g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_14),
.C(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_5),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_6),
.B(n_9),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_14),
.C(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_62),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_67),
.B(n_63),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_10),
.B(n_12),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_79),
.C(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_99),
.B(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_55),
.B1(n_60),
.B2(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_86),
.B1(n_82),
.B2(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_52),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_78),
.C(n_87),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_81),
.B1(n_93),
.B2(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_80),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_98),
.C(n_89),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_95),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_103),
.B(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_122),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_114),
.Y(n_122)
);

AOI31xp33_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_100),
.A3(n_104),
.B(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_108),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_116),
.B(n_119),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_126),
.B(n_76),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_122),
.C(n_114),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_128),
.B(n_76),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_52),
.Y(n_130)
);


endmodule