module fake_jpeg_2884_n_187 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_32),
.B(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_54),
.Y(n_61)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_12),
.B(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_51),
.Y(n_68)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_16),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_39),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_24),
.B1(n_25),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_24),
.B1(n_25),
.B2(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_30),
.A2(n_15),
.B1(n_16),
.B2(n_5),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_15),
.B1(n_16),
.B2(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_32),
.A2(n_16),
.B1(n_4),
.B2(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_3),
.B1(n_40),
.B2(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_31),
.B(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_21),
.B1(n_24),
.B2(n_36),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_96),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_50),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_71),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_122)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_70),
.B(n_82),
.C(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_75),
.B1(n_79),
.B2(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_121),
.B1(n_102),
.B2(n_59),
.Y(n_145)
);

NAND2xp67_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_123),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_90),
.B(n_63),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_79),
.B1(n_90),
.B2(n_78),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_67),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_59),
.B1(n_78),
.B2(n_86),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_133),
.B1(n_112),
.B2(n_101),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_59),
.B1(n_78),
.B2(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_143),
.Y(n_154)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_96),
.A3(n_91),
.B1(n_99),
.B2(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_137),
.C(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_111),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_147),
.A3(n_119),
.B1(n_118),
.B2(n_125),
.C1(n_128),
.C2(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_99),
.B1(n_89),
.B2(n_80),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_156),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_123),
.C(n_122),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_142),
.B(n_136),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_163),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_136),
.B(n_134),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_153),
.B1(n_147),
.B2(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_169),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_153),
.B1(n_132),
.B2(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_159),
.A3(n_151),
.B(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_170),
.B1(n_121),
.B2(n_123),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_179),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_170),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_138),
.B(n_125),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_129),
.B(n_130),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_180),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_177),
.CI(n_129),
.CON(n_187),
.SN(n_187)
);


endmodule