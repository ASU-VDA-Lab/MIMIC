module fake_jpeg_29499_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_11),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_26),
.B1(n_6),
.B2(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

AO221x1_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_22),
.C(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_25),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.C(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_6),
.B(n_7),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_8),
.Y(n_37)
);


endmodule