module fake_netlist_1_1463_n_694 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_694);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_694;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_57), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_65), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_61), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_43), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_52), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_31), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_0), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_3), .Y(n_86) );
BUFx10_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_69), .Y(n_89) );
INVx1_ASAP7_75t_SL g90 ( .A(n_42), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_15), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_50), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_23), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_35), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_4), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_70), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_49), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_59), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_27), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_53), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_21), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_26), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_68), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_0), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_58), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_14), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_39), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_96), .B(n_1), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_96), .B(n_1), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_114), .Y(n_128) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_79), .A2(n_28), .B(n_75), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_93), .B(n_2), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_89), .B(n_3), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_80), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_102), .B(n_5), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_79), .B(n_6), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_77), .B(n_7), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_83), .B(n_9), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_78), .B(n_9), .Y(n_145) );
BUFx8_ASAP7_75t_L g146 ( .A(n_109), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_106), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_85), .B(n_10), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_98), .B(n_11), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_104), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_92), .B(n_11), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_85), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_86), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_113), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_86), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_126), .B(n_88), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
CKINVDCx6p67_ASAP7_75t_R g174 ( .A(n_152), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_128), .B(n_124), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_128), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_126), .B(n_107), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_127), .B(n_107), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_152), .B(n_123), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_162), .B(n_163), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_166), .B(n_110), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_130), .A2(n_117), .B1(n_88), .B2(n_120), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_127), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_136), .A2(n_112), .B1(n_117), .B2(n_111), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_127), .B(n_120), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_152), .B(n_91), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_127), .B(n_120), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_130), .A2(n_120), .B1(n_119), .B2(n_116), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_133), .B(n_120), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_125), .B(n_87), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_146), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_133), .B(n_138), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_136), .A2(n_87), .B1(n_99), .B2(n_100), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_138), .B(n_108), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_144), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_134), .B(n_87), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_153), .B(n_164), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_148), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_148), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_157), .Y(n_227) );
AND2x6_ASAP7_75t_L g228 ( .A(n_134), .B(n_90), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_218), .B(n_160), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_216), .B(n_209), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_189), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g232 ( .A(n_213), .B(n_146), .C(n_160), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_216), .B(n_146), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_178), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_185), .B(n_164), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_178), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_205), .A2(n_132), .B1(n_159), .B2(n_158), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_216), .B(n_161), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_169), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_209), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_206), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_161), .B1(n_159), .B2(n_158), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_187), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_206), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_169), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_218), .B(n_154), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_168), .A2(n_153), .B1(n_156), .B2(n_154), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_185), .B(n_151), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_205), .B(n_156), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_206), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_173), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_193), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_216), .B(n_140), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_173), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_212), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_187), .Y(n_263) );
NOR2xp67_ASAP7_75t_L g264 ( .A(n_213), .B(n_145), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_212), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_186), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_188), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_186), .Y(n_269) );
CKINVDCx11_ASAP7_75t_R g270 ( .A(n_193), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_167), .B(n_151), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_195), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_198), .B(n_155), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_179), .B(n_137), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_174), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_174), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_179), .A2(n_141), .B1(n_150), .B2(n_149), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_182), .B(n_101), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_188), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_195), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_172), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_188), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_168), .A2(n_139), .B1(n_150), .B2(n_149), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_198), .B(n_84), .Y(n_286) );
BUFx8_ASAP7_75t_L g287 ( .A(n_175), .Y(n_287) );
BUFx4f_ASAP7_75t_SL g288 ( .A(n_174), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_168), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_183), .B(n_118), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_195), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_179), .B(n_97), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_168), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_188), .Y(n_294) );
OR2x6_ASAP7_75t_L g295 ( .A(n_289), .B(n_167), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
AND2x2_ASAP7_75t_SL g297 ( .A(n_292), .B(n_167), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_253), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_282), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_276), .B(n_167), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_261), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_231), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_248), .B(n_179), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_251), .B(n_175), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_276), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_248), .B(n_181), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_234), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_240), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_261), .Y(n_315) );
AOI21x1_ASAP7_75t_L g316 ( .A1(n_280), .A2(n_226), .B(n_225), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_253), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_253), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_234), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_253), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_280), .A2(n_170), .B(n_172), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_232), .B(n_203), .C(n_191), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_254), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_262), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_230), .A2(n_271), .B1(n_251), .B2(n_257), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_277), .B(n_191), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_291), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_235), .B(n_224), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_271), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_256), .A2(n_228), .B1(n_168), .B2(n_191), .Y(n_332) );
AOI22x1_ASAP7_75t_L g333 ( .A1(n_242), .A2(n_188), .B1(n_191), .B2(n_172), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_248), .B(n_181), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_252), .B(n_228), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_271), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_235), .B(n_181), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_264), .A2(n_228), .B1(n_168), .B2(n_181), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_237), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_237), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_293), .B(n_202), .Y(n_342) );
AOI21xp5_ASAP7_75t_SL g343 ( .A1(n_242), .A2(n_170), .B(n_202), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_263), .A2(n_228), .B1(n_168), .B2(n_203), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_287), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_300), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_326), .A2(n_256), .B1(n_287), .B2(n_244), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_271), .B1(n_260), .B2(n_269), .Y(n_349) );
OAI21xp33_ASAP7_75t_SL g350 ( .A1(n_303), .A2(n_260), .B(n_250), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_306), .A2(n_270), .B1(n_244), .B2(n_287), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_340), .A2(n_270), .B1(n_228), .B2(n_292), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_329), .A2(n_229), .B1(n_239), .B2(n_238), .C(n_279), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_306), .A2(n_229), .B1(n_292), .B2(n_228), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_337), .B(n_229), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_306), .A2(n_334), .B1(n_310), .B2(n_297), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_228), .B1(n_275), .B2(n_291), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_298), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_314), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_340), .A2(n_233), .B1(n_274), .B2(n_249), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_334), .A2(n_297), .B1(n_308), .B2(n_313), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_334), .A2(n_228), .B1(n_275), .B2(n_236), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_330), .B(n_275), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_341), .A2(n_241), .B1(n_286), .B2(n_273), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_302), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_302), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_330), .B(n_246), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_336), .B(n_246), .Y(n_376) );
AO22x1_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_345), .B1(n_319), .B2(n_307), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_255), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_350), .A2(n_323), .B(n_335), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_338), .B(n_344), .C(n_336), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_332), .B1(n_304), .B2(n_315), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_305), .B1(n_315), .B2(n_304), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_355), .A2(n_307), .B1(n_312), .B2(n_309), .Y(n_384) );
AOI33xp33_ASAP7_75t_L g385 ( .A1(n_348), .A2(n_190), .A3(n_202), .B1(n_285), .B2(n_272), .B3(n_268), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_202), .B1(n_278), .B2(n_172), .C1(n_190), .C2(n_322), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_352), .A2(n_357), .B1(n_363), .B2(n_368), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_365), .A2(n_307), .B1(n_350), .B2(n_370), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_225), .B1(n_220), .B2(n_226), .C(n_222), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_347), .B(n_311), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_370), .A2(n_312), .B1(n_295), .B2(n_290), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_367), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_352), .A2(n_266), .B1(n_269), .B2(n_255), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_331), .B1(n_328), .B2(n_312), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_321), .B(n_294), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_371), .A2(n_343), .B(n_243), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_362), .A2(n_294), .B(n_284), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_351), .A2(n_259), .B1(n_258), .B2(n_247), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_381), .A2(n_358), .B1(n_359), .B2(n_360), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_381), .A2(n_365), .B1(n_374), .B2(n_376), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_388), .B(n_364), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_382), .A2(n_358), .B1(n_222), .B2(n_247), .C(n_373), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_389), .A2(n_247), .B1(n_375), .B2(n_373), .C(n_372), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_377), .A2(n_97), .B(n_99), .C(n_100), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_388), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_396), .A2(n_376), .B1(n_374), .B2(n_364), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_401), .A2(n_375), .B1(n_372), .B2(n_361), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_378), .B(n_369), .Y(n_415) );
AO22x1_ASAP7_75t_L g416 ( .A1(n_383), .A2(n_369), .B1(n_364), .B2(n_367), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_378), .B(n_369), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_393), .A2(n_327), .A3(n_301), .B(n_183), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_403), .B(n_266), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_390), .B(n_118), .C(n_157), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_316), .B(n_343), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_384), .B(n_301), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_394), .A2(n_200), .A3(n_196), .B1(n_197), .B2(n_199), .B3(n_208), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_396), .A2(n_361), .B1(n_327), .B2(n_295), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_401), .A2(n_398), .B1(n_391), .B2(n_386), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_387), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_380), .A2(n_361), .B1(n_295), .B2(n_170), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_361), .B1(n_333), .B2(n_295), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_377), .A2(n_392), .B(n_400), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_397), .B(n_367), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_400), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_404), .A2(n_367), .B1(n_342), .B2(n_325), .Y(n_436) );
INVx5_ASAP7_75t_SL g437 ( .A(n_392), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
AO21x1_ASAP7_75t_SL g439 ( .A1(n_395), .A2(n_367), .B(n_318), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_245), .B1(n_283), .B2(n_293), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_413), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_415), .B(n_385), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_415), .B(n_402), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_342), .A3(n_245), .B(n_298), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_402), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_402), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_411), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_13), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_450) );
OAI222xp33_ASAP7_75t_L g451 ( .A1(n_405), .A2(n_13), .B1(n_16), .B2(n_17), .C1(n_18), .C2(n_284), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_407), .B(n_402), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_418), .B(n_399), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_420), .B(n_367), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_433), .B(n_399), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_410), .B(n_427), .C(n_431), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_437), .A2(n_399), .B1(n_325), .B2(n_320), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_433), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_419), .A2(n_157), .B1(n_298), .B2(n_188), .C(n_399), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_438), .B(n_157), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_438), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_432), .B(n_325), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_422), .B(n_207), .C(n_196), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_434), .B(n_19), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_416), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_432), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_437), .B(n_325), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_434), .B(n_20), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_432), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_437), .B(n_320), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_437), .B(n_320), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_408), .A2(n_207), .B1(n_197), .B2(n_199), .C(n_200), .Y(n_478) );
OAI33xp33_ASAP7_75t_L g479 ( .A1(n_421), .A2(n_208), .A3(n_211), .B1(n_214), .B2(n_219), .B3(n_215), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_409), .B(n_320), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_414), .B(n_201), .C(n_217), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_424), .B(n_207), .C(n_211), .D(n_214), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_423), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_436), .Y(n_487) );
BUFx2_ASAP7_75t_SL g488 ( .A(n_439), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
OAI33xp33_ASAP7_75t_L g490 ( .A1(n_429), .A2(n_176), .A3(n_227), .B1(n_223), .B2(n_219), .B3(n_215), .Y(n_490) );
NAND5xp2_ASAP7_75t_SL g491 ( .A(n_430), .B(n_22), .C(n_24), .D(n_25), .E(n_29), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_457), .A2(n_425), .B1(n_440), .B2(n_267), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_460), .B(n_318), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_443), .B(n_318), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_488), .B(n_318), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_488), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_317), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_457), .B(n_180), .C(n_227), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_447), .B(n_317), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
AND2x4_ASAP7_75t_SL g504 ( .A(n_489), .B(n_317), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_447), .B(n_30), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_445), .B(n_317), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_452), .B(n_32), .Y(n_507) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_489), .A2(n_180), .B(n_171), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_450), .B(n_180), .C(n_227), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
AND2x4_ASAP7_75t_SL g511 ( .A(n_489), .B(n_296), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_299), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_471), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_484), .A2(n_296), .B(n_299), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_459), .A2(n_177), .B(n_171), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_454), .B(n_33), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
AND3x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_34), .C(n_37), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_451), .A2(n_192), .A3(n_223), .B(n_219), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_442), .B(n_299), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_454), .B(n_458), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_485), .B(n_184), .C(n_223), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_454), .B(n_299), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_467), .B(n_296), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_458), .B(n_474), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_482), .B(n_38), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_476), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_467), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_469), .B(n_40), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_441), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_441), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g537 ( .A(n_469), .B(n_267), .Y(n_537) );
AOI31xp33_ASAP7_75t_L g538 ( .A1(n_475), .A2(n_41), .A3(n_44), .B(n_48), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_476), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_449), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_487), .A2(n_267), .B1(n_265), .B2(n_262), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_462), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_473), .B(n_51), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_484), .A2(n_267), .B(n_265), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_462), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_453), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_475), .A2(n_194), .B(n_192), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_455), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_464), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_533), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_514), .B(n_455), .Y(n_552) );
AND3x1_ASAP7_75t_L g553 ( .A(n_500), .B(n_444), .C(n_473), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_498), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_533), .Y(n_555) );
OAI21xp5_ASAP7_75t_SL g556 ( .A1(n_538), .A2(n_461), .B(n_455), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_513), .B(n_483), .Y(n_557) );
NOR2x1p5_ASAP7_75t_L g558 ( .A(n_518), .B(n_472), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_502), .B(n_483), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_495), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_510), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_502), .B(n_486), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_537), .B(n_455), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_527), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_516), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_547), .B(n_486), .Y(n_567) );
OR2x6_ASAP7_75t_L g568 ( .A(n_523), .B(n_480), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_547), .B(n_464), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_539), .B(n_480), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_531), .B(n_466), .Y(n_571) );
AOI32xp33_ASAP7_75t_L g572 ( .A1(n_537), .A2(n_468), .A3(n_491), .B1(n_477), .B2(n_481), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_494), .B(n_479), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_528), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_504), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_494), .B(n_54), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_500), .B(n_490), .C(n_491), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_519), .B(n_67), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_529), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_519), .B(n_478), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_549), .B(n_71), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_534), .B(n_73), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_535), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_505), .B(n_76), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_536), .B(n_171), .Y(n_587) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_523), .B(n_267), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_540), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_507), .B(n_176), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_492), .B(n_201), .C(n_221), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_546), .B(n_176), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_543), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_544), .B(n_265), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_497), .A2(n_265), .B1(n_262), .B2(n_207), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_504), .B(n_177), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_550), .B(n_177), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_522), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_506), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_550), .B(n_184), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_565), .B(n_496), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_554), .B(n_530), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_560), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_561), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
XNOR2x2_ASAP7_75t_L g608 ( .A(n_575), .B(n_525), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_551), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_553), .A2(n_492), .B1(n_524), .B2(n_518), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_566), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_552), .B(n_499), .Y(n_613) );
OAI32xp33_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_525), .A3(n_493), .B1(n_501), .B2(n_512), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_557), .B(n_526), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_555), .B(n_497), .Y(n_616) );
NAND2x1_ASAP7_75t_L g617 ( .A(n_568), .B(n_497), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_574), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_579), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_559), .B(n_511), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_568), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_589), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_591), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_583), .B(n_511), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_555), .B(n_518), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_563), .B(n_520), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_585), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_581), .B(n_517), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_567), .B(n_520), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_581), .B(n_515), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_569), .B(n_541), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_601), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_558), .B(n_524), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_600), .B(n_548), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_571), .B(n_509), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_594), .B(n_509), .Y(n_639) );
AOI211xp5_ASAP7_75t_SL g640 ( .A1(n_556), .A2(n_545), .B(n_521), .C(n_508), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_580), .A2(n_184), .B1(n_192), .B2(n_194), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_564), .A2(n_265), .B(n_262), .C(n_210), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_597), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_572), .A2(n_194), .B(n_210), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_599), .Y(n_645) );
XOR2x2_ASAP7_75t_L g646 ( .A(n_588), .B(n_262), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_568), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_564), .B(n_210), .Y(n_648) );
OAI31xp33_ASAP7_75t_SL g649 ( .A1(n_592), .A2(n_215), .A3(n_201), .B(n_217), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_587), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_578), .A2(n_201), .B1(n_217), .B2(n_221), .C1(n_595), .C2(n_576), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_593), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_597), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_577), .A2(n_201), .B(n_217), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_578), .B(n_201), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_595), .A2(n_217), .B(n_221), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_598), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_602), .B(n_217), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_586), .Y(n_659) );
NAND4xp25_ASAP7_75t_SL g660 ( .A(n_582), .B(n_221), .C(n_590), .D(n_596), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g661 ( .A1(n_654), .A2(n_625), .B(n_614), .C(n_660), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_659), .Y(n_662) );
AOI21xp33_ASAP7_75t_SL g663 ( .A1(n_634), .A2(n_610), .B(n_649), .Y(n_663) );
OAI22x1_ASAP7_75t_L g664 ( .A1(n_621), .A2(n_604), .B1(n_608), .B2(n_636), .Y(n_664) );
NOR4xp25_ASAP7_75t_L g665 ( .A(n_611), .B(n_627), .C(n_639), .D(n_633), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_637), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_640), .A2(n_656), .B(n_638), .Y(n_667) );
NAND4xp25_ASAP7_75t_SL g668 ( .A(n_651), .B(n_627), .C(n_630), .D(n_656), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_617), .B(n_621), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_643), .A2(n_637), .B(n_653), .C(n_611), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g672 ( .A(n_642), .B(n_630), .C(n_644), .Y(n_672) );
AOI32xp33_ASAP7_75t_L g673 ( .A1(n_603), .A2(n_643), .A3(n_647), .B1(n_653), .B2(n_620), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_669), .A2(n_609), .A3(n_622), .B1(n_605), .B2(n_606), .C1(n_607), .C2(n_619), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_662), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_665), .A2(n_612), .B1(n_618), .B2(n_623), .C(n_624), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_666), .A2(n_647), .A3(n_613), .B1(n_615), .B2(n_635), .C1(n_620), .C2(n_652), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_671), .A2(n_626), .B1(n_631), .B2(n_616), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_672), .A2(n_615), .A3(n_650), .B1(n_657), .B2(n_645), .C1(n_655), .C2(n_641), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_670), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_664), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_675), .B(n_668), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_681), .A2(n_667), .B1(n_661), .B2(n_663), .Y(n_683) );
AND4x1_ASAP7_75t_L g684 ( .A(n_676), .B(n_667), .C(n_673), .D(n_658), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_678), .A2(n_632), .B1(n_629), .B2(n_642), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_682), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_683), .B(n_680), .C(n_648), .Y(n_687) );
OR3x2_ASAP7_75t_L g688 ( .A(n_684), .B(n_679), .C(n_677), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_686), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_687), .B(n_685), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_688), .B1(n_646), .B2(n_674), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_691), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_692), .Y(n_693) );
AOI221xp5_ASAP7_75t_SL g694 ( .A1(n_693), .A2(n_221), .B1(n_596), .B2(n_689), .C(n_691), .Y(n_694) );
endmodule