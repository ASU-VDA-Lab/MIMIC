module real_jpeg_4417_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_1),
.B(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_4),
.B(n_34),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_5),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_9),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_90),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_134),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_13),
.Y(n_118)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_14),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_14),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_14),
.B(n_34),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_123),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_51),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_30),
.C(n_33),
.Y(n_80)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_31),
.Y(n_131)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_35),
.Y(n_189)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_38),
.A2(n_39),
.B1(n_51),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.C(n_49),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_40),
.A2(n_41),
.B1(n_49),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_45),
.B(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_49),
.Y(n_210)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_78),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_103),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.C(n_97),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_98),
.Y(n_139)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_109),
.B1(n_121),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_116),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_138),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_125),
.B(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_128),
.B(n_138),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_132),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_130),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_135),
.Y(n_184)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_212),
.B(n_216),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_198),
.B(n_211),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_181),
.B(n_197),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_164),
.B(n_180),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_160),
.B(n_163),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_155),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_196),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_196),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_185),
.C(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_206),
.C(n_207),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_205),
.C(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);


endmodule