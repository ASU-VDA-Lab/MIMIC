module fake_jpeg_2914_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_103),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_83),
.C(n_76),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_80),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_67),
.B1(n_55),
.B2(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_105),
.B1(n_61),
.B2(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_57),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_57),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_53),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_82),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_67),
.B1(n_65),
.B2(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_64),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_91),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_119),
.C(n_123),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_118),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_82),
.B1(n_53),
.B2(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_66),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_51),
.B(n_54),
.Y(n_119)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_56),
.B1(n_44),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_58),
.B(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_0),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_136),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_97),
.B1(n_100),
.B2(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_134),
.B1(n_141),
.B2(n_7),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_41),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_11),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_143),
.B1(n_121),
.B2(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_151),
.B1(n_137),
.B2(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_34),
.C(n_32),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_31),
.B(n_29),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_28),
.C(n_26),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_21),
.C(n_19),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_11),
.CI(n_12),
.CON(n_167),
.SN(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_130),
.B(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_129),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_171),
.B1(n_172),
.B2(n_148),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_162),
.B(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_168),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_155),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_175),
.B(n_179),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_163),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_180),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_150),
.C(n_154),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_164),
.B1(n_160),
.B2(n_167),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_183),
.B(n_164),
.C(n_184),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_182),
.C(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_13),
.C(n_14),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_15),
.C(n_16),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_17),
.Y(n_193)
);


endmodule