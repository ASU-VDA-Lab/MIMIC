module fake_jpeg_14154_n_132 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_29),
.B(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_45),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_14),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_25),
.B1(n_24),
.B2(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_16),
.Y(n_54)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_22),
.B(n_5),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_7),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_23),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_33),
.B(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_70),
.B1(n_59),
.B2(n_61),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_62),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_17),
.B(n_24),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_71),
.C(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_25),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_41),
.B1(n_54),
.B2(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_56),
.B1(n_60),
.B2(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_75),
.B1(n_55),
.B2(n_53),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_56),
.B1(n_86),
.B2(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_85),
.B1(n_78),
.B2(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_86),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_111),
.B1(n_106),
.B2(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_83),
.B1(n_78),
.B2(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_99),
.B1(n_98),
.B2(n_100),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_91),
.B(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_96),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_113),
.B1(n_112),
.B2(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_112),
.B1(n_107),
.B2(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_97),
.B1(n_119),
.B2(n_117),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_117),
.B(n_120),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_122),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_129),
.B(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_120),
.Y(n_132)
);


endmodule