module fake_jpeg_28920_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx24_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_17),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_42),
.B1(n_31),
.B2(n_30),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_10),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_14),
.B1(n_22),
.B2(n_15),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_61),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_30),
.B(n_13),
.C(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_60),
.B1(n_34),
.B2(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_32),
.B1(n_15),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_40),
.B1(n_29),
.B2(n_37),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_30),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_29),
.B1(n_31),
.B2(n_14),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_86),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_69),
.B(n_70),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_71),
.B(n_1),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_58),
.B1(n_50),
.B2(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_67),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_56),
.B1(n_63),
.B2(n_55),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_75),
.B(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_56),
.B1(n_63),
.B2(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_79),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_48),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_65),
.C(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_76),
.B1(n_79),
.B2(n_77),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_81),
.A3(n_82),
.B1(n_10),
.B2(n_9),
.C1(n_73),
.C2(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_0),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_95),
.C(n_93),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_103),
.B1(n_107),
.B2(n_88),
.C(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_86),
.B1(n_93),
.B2(n_87),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_105),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_77),
.B(n_2),
.Y(n_107)
);

AOI211xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_107),
.B(n_100),
.C(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_90),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_112),
.B(n_3),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_93),
.B1(n_96),
.B2(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_115),
.B1(n_106),
.B2(n_4),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_99),
.C(n_102),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_120),
.C(n_5),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_86),
.C(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_115),
.C(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_114),
.B1(n_110),
.B2(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_6),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.C(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_3),
.C(n_5),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_3),
.B(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_124),
.C(n_6),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_7),
.Y(n_137)
);


endmodule