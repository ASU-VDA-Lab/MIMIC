module fake_netlist_6_2344_n_1724 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1724);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1724;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_22),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_38),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_72),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_20),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_33),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_11),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_19),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_89),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_47),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_54),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_96),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_56),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_93),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_53),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_26),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_28),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_1),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_32),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_77),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_98),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_49),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_17),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_90),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_17),
.Y(n_206)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_62),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_54),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_38),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_19),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_33),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_29),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_120),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_86),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_102),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_138),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_15),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_63),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_132),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_135),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_139),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_34),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_30),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_105),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

BUFx2_ASAP7_75t_SL g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_142),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_34),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_131),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_49),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_36),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_79),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_68),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_134),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_149),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_51),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_22),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_7),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_67),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_136),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_121),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_82),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_21),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_150),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_117),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_58),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_125),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_16),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_152),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_111),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_31),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_27),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_85),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_56),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_14),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_88),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_51),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_115),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_55),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_65),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_42),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_151),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_108),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_119),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_29),
.Y(n_293)
);

BUFx2_ASAP7_75t_SL g294 ( 
.A(n_41),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_104),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_106),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_124),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_122),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_55),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_123),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_100),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_112),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_14),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_107),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_168),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_179),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_179),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_170),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_179),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_169),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_179),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_153),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_169),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_190),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_177),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_179),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_160),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_155),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_193),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_179),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_179),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_213),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_213),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_213),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_213),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_257),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_295),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_292),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_260),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_197),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_155),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_159),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_265),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_184),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_208),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_209),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_209),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_230),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_215),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_237),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_159),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_237),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_223),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_228),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_249),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_249),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_162),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_292),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_275),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_275),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_162),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_307),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_277),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_232),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_299),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_235),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_177),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_363),
.B(n_368),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

OR2x6_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_207),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_329),
.Y(n_389)
);

BUFx8_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_366),
.B(n_238),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_338),
.B(n_198),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_370),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_313),
.B(n_197),
.Y(n_406)
);

BUFx12f_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_316),
.B(n_198),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_197),
.Y(n_412)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_346),
.B(n_271),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_311),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_271),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_319),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_347),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_324),
.Y(n_424)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_368),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_348),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_324),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_325),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_326),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_321),
.B(n_202),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_351),
.B(n_276),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_337),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_306),
.B1(n_308),
.B2(n_276),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_406),
.A2(n_306),
.B1(n_365),
.B2(n_342),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_349),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_377),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_421),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_356),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_419),
.B(n_360),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_387),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_361),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_428),
.B(n_341),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_434),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_400),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_396),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_399),
.A2(n_194),
.B1(n_241),
.B2(n_303),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_380),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

AO22x1_ASAP7_75t_L g477 ( 
.A1(n_420),
.A2(n_274),
.B1(n_247),
.B2(n_250),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g478 ( 
.A1(n_435),
.A2(n_240),
.B1(n_251),
.B2(n_278),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_428),
.B(n_353),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_428),
.B(n_373),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_410),
.B(n_199),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_403),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_428),
.B(n_376),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_380),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_410),
.A2(n_172),
.B1(n_164),
.B2(n_175),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_420),
.B(n_437),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_403),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_428),
.B(n_343),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_407),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_422),
.B(n_229),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_315),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_380),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_398),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_428),
.B(n_156),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_422),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_255),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_429),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_382),
.B(n_234),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_382),
.B(n_294),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_380),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_322),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_433),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_400),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_264),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_R g527 ( 
.A(n_384),
.B(n_443),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_428),
.B(n_156),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_439),
.B(n_330),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_385),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_407),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_418),
.B(n_420),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_380),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_385),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_388),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_305),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_435),
.A2(n_382),
.B1(n_400),
.B2(n_413),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_380),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_416),
.B(n_218),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_380),
.B(n_242),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_384),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_382),
.A2(n_204),
.B1(n_231),
.B2(n_224),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_437),
.A2(n_288),
.B1(n_186),
.B2(n_212),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_382),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_395),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_428),
.B(n_157),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_381),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_390),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_381),
.B(n_281),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_397),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_381),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_395),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_384),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_412),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_389),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_413),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_437),
.A2(n_263),
.B1(n_273),
.B2(n_244),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_381),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_398),
.B(n_355),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_381),
.B(n_283),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_389),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_381),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_412),
.B(n_244),
.Y(n_574)
);

AO22x1_ASAP7_75t_L g575 ( 
.A1(n_437),
.A2(n_183),
.B1(n_178),
.B2(n_166),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_397),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_381),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_381),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_386),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_386),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_391),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_386),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_386),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_386),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_386),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_391),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_394),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_386),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_386),
.B(n_285),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_393),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_382),
.B(n_332),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_447),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_493),
.B(n_382),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_447),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_493),
.B(n_393),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_454),
.B(n_413),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_287),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_445),
.A2(n_413),
.B1(n_425),
.B2(n_335),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_459),
.B(n_393),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_570),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_540),
.B(n_390),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_459),
.B(n_393),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_470),
.B(n_425),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_447),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_470),
.B(n_443),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_464),
.B(n_393),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_445),
.A2(n_417),
.B(n_437),
.C(n_161),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_448),
.B(n_425),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_393),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_466),
.B(n_393),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_455),
.B(n_425),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_456),
.A2(n_256),
.B1(n_412),
.B2(n_167),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_466),
.B(n_393),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_503),
.B(n_390),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_456),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_468),
.B(n_405),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_450),
.B(n_405),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_487),
.B(n_509),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_574),
.B(n_218),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_449),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_488),
.B(n_379),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_457),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_574),
.A2(n_256),
.B1(n_412),
.B2(n_182),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_535),
.B(n_451),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_570),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_527),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_529),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_449),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_523),
.B(n_425),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_502),
.B(n_405),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_458),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_542),
.B(n_405),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_523),
.B(n_425),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_542),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_507),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_489),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_458),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_506),
.B(n_390),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_574),
.A2(n_412),
.B1(n_252),
.B2(n_188),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_554),
.B(n_166),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_545),
.B(n_405),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_550),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_506),
.B(n_390),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_550),
.B(n_405),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_506),
.B(n_405),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_463),
.A2(n_553),
.B1(n_517),
.B2(n_516),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_506),
.B(n_432),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_548),
.B(n_443),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_551),
.A2(n_217),
.B(n_266),
.C(n_225),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_549),
.B(n_379),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_458),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_565),
.B(n_432),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_565),
.B(n_432),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_560),
.A2(n_417),
.B(n_432),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_572),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_530),
.B(n_432),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

BUFx4f_ASAP7_75t_L g664 ( 
.A(n_517),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_461),
.B(n_431),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_548),
.B(n_431),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_563),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_553),
.A2(n_517),
.B1(n_516),
.B2(n_480),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_516),
.A2(n_154),
.B1(n_219),
.B2(n_216),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_561),
.B(n_157),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_431),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_446),
.B(n_436),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_581),
.B(n_432),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_530),
.B(n_163),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_494),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_513),
.B(n_163),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_586),
.B(n_587),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_574),
.A2(n_205),
.B1(n_293),
.B2(n_282),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_586),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_530),
.B(n_171),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_587),
.B(n_432),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_473),
.B(n_476),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_532),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_460),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_574),
.A2(n_218),
.B1(n_239),
.B2(n_246),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_574),
.A2(n_516),
.B1(n_472),
.B2(n_492),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_SL g688 ( 
.A(n_566),
.B(n_218),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_507),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_516),
.A2(n_218),
.B1(n_239),
.B2(n_246),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_460),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_585),
.A2(n_404),
.B(n_394),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_476),
.B(n_432),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_530),
.B(n_239),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_526),
.B(n_171),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_566),
.B(n_239),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_482),
.B(n_401),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_482),
.B(n_401),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_483),
.B(n_239),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_537),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_537),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_483),
.B(n_246),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_496),
.B(n_402),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_567),
.A2(n_246),
.B1(n_203),
.B2(n_165),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_539),
.B(n_173),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_496),
.B(n_402),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_521),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_462),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_507),
.Y(n_709)
);

OAI21xp33_ASAP7_75t_L g710 ( 
.A1(n_444),
.A2(n_270),
.B(n_227),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_499),
.B(n_510),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_499),
.B(n_510),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_512),
.B(n_404),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_477),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_462),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_512),
.B(n_408),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_462),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_518),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_465),
.B(n_173),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_552),
.B(n_201),
.C(n_279),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_538),
.Y(n_721)
);

OAI221xp5_ASAP7_75t_L g722 ( 
.A1(n_544),
.A2(n_296),
.B1(n_302),
.B2(n_158),
.C(n_272),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_525),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_562),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_553),
.A2(n_269),
.B1(n_267),
.B2(n_262),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_525),
.B(n_408),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_546),
.B(n_246),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_525),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_534),
.B(n_409),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_478),
.B(n_497),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_481),
.B(n_174),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_531),
.Y(n_732)
);

BUFx5_ASAP7_75t_L g733 ( 
.A(n_515),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_534),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_553),
.A2(n_269),
.B1(n_187),
.B2(n_185),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_534),
.B(n_409),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_575),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_491),
.B(n_411),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_SL g739 ( 
.A(n_490),
.B(n_178),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_471),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_517),
.A2(n_291),
.B1(n_289),
.B2(n_270),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_491),
.B(n_411),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_491),
.B(n_415),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_515),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_471),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_591),
.B(n_195),
.C(n_192),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_189),
.C(n_280),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_579),
.B(n_174),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_517),
.B(n_176),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_511),
.B(n_176),
.Y(n_750)
);

AO221x1_ASAP7_75t_L g751 ( 
.A1(n_491),
.A2(n_590),
.B1(n_520),
.B2(n_541),
.C(n_583),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_579),
.B(n_436),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_579),
.B(n_180),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_477),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_520),
.B(n_415),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_557),
.B(n_183),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_621),
.A2(n_555),
.B1(n_528),
.B2(n_558),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_692),
.A2(n_589),
.B(n_571),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_730),
.A2(n_522),
.B1(n_524),
.B2(n_467),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_730),
.B(n_584),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_639),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_621),
.B(n_590),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_752),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_679),
.A2(n_498),
.B1(n_484),
.B2(n_533),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_597),
.A2(n_590),
.B1(n_573),
.B2(n_556),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_667),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_597),
.A2(n_590),
.B1(n_573),
.B2(n_556),
.Y(n_767)
);

NOR2x2_ASAP7_75t_L g768 ( 
.A(n_679),
.B(n_227),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_666),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_665),
.B(n_180),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_752),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_584),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_611),
.B(n_520),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_672),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_655),
.A2(n_522),
.B1(n_524),
.B2(n_467),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_653),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_655),
.A2(n_452),
.B1(n_453),
.B2(n_469),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_611),
.B(n_520),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_634),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_707),
.B(n_541),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_710),
.A2(n_268),
.B(n_261),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_601),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_614),
.B(n_584),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_690),
.A2(n_741),
.B1(n_626),
.B2(n_618),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_638),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_607),
.B(n_629),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_639),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_684),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_614),
.A2(n_588),
.B(n_583),
.C(n_580),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_700),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_625),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_701),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_640),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_626),
.B(n_588),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_594),
.B(n_588),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_583),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_677),
.B(n_583),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_639),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_639),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_721),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_651),
.B(n_605),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_593),
.A2(n_573),
.B1(n_580),
.B2(n_556),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_604),
.B(n_609),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_628),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_695),
.B(n_541),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_689),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_687),
.B(n_541),
.Y(n_808)
);

BUFx4f_ASAP7_75t_SL g809 ( 
.A(n_676),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_695),
.A2(n_580),
.B(n_573),
.C(n_556),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_705),
.B(n_580),
.Y(n_811)
);

AND2x2_ASAP7_75t_SL g812 ( 
.A(n_690),
.B(n_505),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_705),
.B(n_452),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_724),
.Y(n_814)
);

BUFx4f_ASAP7_75t_L g815 ( 
.A(n_714),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_689),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_660),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_741),
.A2(n_686),
.B1(n_751),
.B2(n_704),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_754),
.Y(n_819)
);

AND3x1_ASAP7_75t_L g820 ( 
.A(n_746),
.B(n_359),
.C(n_355),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_661),
.B(n_438),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_644),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_SL g823 ( 
.A(n_747),
.B(n_268),
.C(n_261),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_670),
.B(n_469),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_689),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_680),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_673),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_732),
.B(n_505),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_683),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_624),
.B(n_181),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_739),
.B(n_181),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_686),
.A2(n_485),
.B1(n_253),
.B2(n_254),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_737),
.B(n_258),
.C(n_248),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_678),
.B(n_485),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_689),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_709),
.B(n_438),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_592),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_709),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_687),
.B(n_649),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_756),
.Y(n_840)
);

NOR2x1p5_ASAP7_75t_L g841 ( 
.A(n_720),
.B(n_253),
.Y(n_841)
);

AND2x6_ASAP7_75t_L g842 ( 
.A(n_632),
.B(n_518),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_627),
.B(n_471),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_704),
.A2(n_254),
.B1(n_475),
.B2(n_479),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_748),
.A2(n_508),
.B(n_475),
.C(n_479),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_620),
.B(n_475),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_711),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_596),
.B(n_479),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_712),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_649),
.B(n_518),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_709),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_712),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_649),
.B(n_518),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_719),
.B(n_543),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_744),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_615),
.B(n_357),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_709),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_649),
.B(n_518),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_664),
.A2(n_284),
.B1(n_196),
.B2(n_210),
.Y(n_859)
);

AO22x1_ASAP7_75t_L g860 ( 
.A1(n_749),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_860)
);

BUFx12f_ASAP7_75t_SL g861 ( 
.A(n_723),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_728),
.A2(n_505),
.B1(n_578),
.B2(n_577),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_649),
.B(n_518),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_664),
.A2(n_233),
.B1(n_236),
.B2(n_243),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_595),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_723),
.B(n_357),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_671),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_719),
.A2(n_486),
.B(n_495),
.C(n_500),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_599),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_606),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_R g871 ( 
.A(n_632),
.B(n_185),
.Y(n_871)
);

NOR2x1p5_ASAP7_75t_L g872 ( 
.A(n_734),
.B(n_286),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_617),
.A2(n_505),
.B1(n_578),
.B2(n_577),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_723),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_617),
.A2(n_569),
.B1(n_578),
.B2(n_577),
.Y(n_875)
);

NAND2x1_ASAP7_75t_L g876 ( 
.A(n_723),
.B(n_536),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_633),
.A2(n_519),
.B(n_500),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_646),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_615),
.A2(n_486),
.B1(n_495),
.B2(n_500),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_649),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_733),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_637),
.B(n_486),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_718),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_623),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_637),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_697),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_731),
.B(n_569),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_643),
.A2(n_725),
.B1(n_735),
.B2(n_749),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_643),
.B(n_495),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_631),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_698),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_635),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_726),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_748),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_753),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_641),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_733),
.B(n_536),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_750),
.A2(n_508),
.B(n_501),
.C(n_504),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_718),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_656),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_602),
.B(n_642),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_L g903 ( 
.A(n_733),
.B(n_536),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_750),
.A2(n_514),
.B1(n_508),
.B2(n_501),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_753),
.B(n_569),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_663),
.Y(n_906)
);

NOR2xp67_ASAP7_75t_L g907 ( 
.A(n_722),
.B(n_543),
.Y(n_907)
);

BUFx8_ASAP7_75t_L g908 ( 
.A(n_685),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_733),
.B(n_501),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_602),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_729),
.B(n_290),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_706),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_691),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_642),
.B(n_359),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_713),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_708),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_SL g917 ( 
.A(n_669),
.B(n_248),
.C(n_245),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_647),
.B(n_362),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_715),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_717),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_647),
.B(n_362),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_733),
.B(n_736),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_610),
.B(n_364),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_622),
.A2(n_519),
.B1(n_514),
.B2(n_504),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_733),
.B(n_504),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_598),
.A2(n_578),
.B1(n_577),
.B2(n_569),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_600),
.B(n_514),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_716),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_603),
.B(n_536),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_608),
.B(n_536),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_612),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_659),
.A2(n_658),
.B(n_613),
.C(n_616),
.Y(n_932)
);

BUFx6f_ASAP7_75t_SL g933 ( 
.A(n_654),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_696),
.B(n_187),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_740),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_619),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_657),
.B(n_519),
.Y(n_937)
);

OR2x2_ASAP7_75t_SL g938 ( 
.A(n_674),
.B(n_364),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_794),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_851),
.B(n_718),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_903),
.A2(n_662),
.B(n_652),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_826),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_827),
.B(n_774),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_785),
.A2(n_839),
.B1(n_881),
.B2(n_812),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_894),
.A2(n_682),
.B(n_645),
.C(n_648),
.Y(n_945)
);

BUFx5_ASAP7_75t_L g946 ( 
.A(n_842),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_783),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_888),
.A2(n_802),
.B1(n_785),
.B2(n_869),
.Y(n_948)
);

NOR2xp67_ASAP7_75t_SL g949 ( 
.A(n_851),
.B(n_718),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_761),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_839),
.A2(n_878),
.B1(n_847),
.B2(n_829),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_864),
.A2(n_681),
.B(n_675),
.C(n_699),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_SL g953 ( 
.A1(n_764),
.A2(n_226),
.B1(n_245),
.B2(n_258),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_881),
.A2(n_650),
.B(n_652),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_792),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_770),
.B(n_745),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_773),
.A2(n_662),
.B(n_650),
.Y(n_957)
);

O2A1O1Ixp5_ASAP7_75t_L g958 ( 
.A1(n_784),
.A2(n_694),
.B(n_688),
.C(n_699),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_776),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_778),
.A2(n_694),
.B(n_636),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_886),
.B(n_755),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_SL g962 ( 
.A1(n_828),
.A2(n_781),
.B(n_887),
.C(n_905),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_855),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_891),
.B(n_738),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_787),
.B(n_742),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_898),
.B(n_743),
.Y(n_966)
);

AO32x1_ASAP7_75t_L g967 ( 
.A1(n_910),
.A2(n_367),
.A3(n_369),
.B1(n_372),
.B2(n_377),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_779),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_761),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_912),
.A2(n_693),
.B(n_702),
.C(n_727),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_780),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_786),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_809),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_851),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_761),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_880),
.A2(n_582),
.B(n_702),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_880),
.A2(n_582),
.B(n_576),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_812),
.A2(n_226),
.B1(n_259),
.B2(n_262),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_769),
.B(n_259),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_819),
.B(n_267),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_818),
.B(n_367),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_864),
.A2(n_833),
.B(n_760),
.C(n_915),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_783),
.B(n_301),
.Y(n_983)
);

OR2x6_ASAP7_75t_SL g984 ( 
.A(n_911),
.B(n_297),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_817),
.B(n_372),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_928),
.B(n_427),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_815),
.B(n_297),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_SL g988 ( 
.A1(n_859),
.A2(n_374),
.B(n_375),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_815),
.B(n_298),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_L g990 ( 
.A(n_833),
.B(n_300),
.C(n_301),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_760),
.A2(n_427),
.B(n_423),
.C(n_576),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_893),
.B(n_423),
.Y(n_992)
);

CKINVDCx8_ASAP7_75t_R g993 ( 
.A(n_761),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_808),
.A2(n_543),
.B(n_576),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_805),
.B(n_300),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_908),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_893),
.B(n_582),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_802),
.A2(n_568),
.B1(n_559),
.B2(n_547),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_867),
.B(n_582),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_807),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_822),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_758),
.A2(n_582),
.B(n_568),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_818),
.A2(n_582),
.B1(n_568),
.B2(n_559),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_559),
.B1(n_547),
.B2(n_441),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_922),
.A2(n_547),
.B(n_474),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_931),
.B(n_441),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_931),
.B(n_441),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_883),
.A2(n_474),
.B(n_442),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_763),
.B(n_101),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_896),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_895),
.A2(n_905),
.B(n_887),
.C(n_849),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_782),
.A2(n_790),
.B(n_781),
.C(n_808),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_801),
.A2(n_375),
.B(n_374),
.C(n_441),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_896),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_883),
.A2(n_474),
.B(n_442),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_861),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_859),
.B(n_474),
.Y(n_1017)
);

INVx8_ASAP7_75t_L g1018 ( 
.A(n_802),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_885),
.B(n_442),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_802),
.A2(n_442),
.B1(n_144),
.B2(n_143),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_442),
.B(n_140),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_920),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_900),
.A2(n_442),
.B(n_126),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_807),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_840),
.B(n_0),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_852),
.A2(n_757),
.B(n_889),
.C(n_856),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_766),
.B(n_442),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_908),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_830),
.A2(n_0),
.B(n_2),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_814),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_821),
.B(n_841),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_823),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_830),
.A2(n_3),
.B(n_5),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_821),
.B(n_3),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_828),
.B(n_6),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_SL g1036 ( 
.A(n_807),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_860),
.B(n_6),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_813),
.A2(n_99),
.B(n_95),
.C(n_94),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_823),
.A2(n_8),
.B(n_9),
.C(n_12),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_854),
.A2(n_442),
.B(n_9),
.C(n_18),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_843),
.A2(n_87),
.B(n_80),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_866),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_866),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_902),
.B(n_78),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_771),
.A2(n_8),
.B1(n_18),
.B2(n_20),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_848),
.A2(n_73),
.B(n_71),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_902),
.B(n_61),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_872),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_918),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_936),
.B(n_23),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_762),
.B(n_25),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_920),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_810),
.A2(n_31),
.B(n_32),
.C(n_37),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_902),
.A2(n_59),
.B1(n_40),
.B2(n_41),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_831),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_846),
.A2(n_897),
.B(n_925),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_871),
.B(n_37),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_820),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_807),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_897),
.A2(n_42),
.B(n_43),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_909),
.A2(n_882),
.B(n_863),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_899),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_899),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1063)
);

BUFx5_ASAP7_75t_L g1064 ( 
.A(n_842),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_768),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_918),
.A2(n_921),
.B(n_811),
.C(n_798),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_824),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_831),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_804),
.B(n_48),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_789),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_836),
.B(n_50),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_797),
.A2(n_50),
.B1(n_52),
.B2(n_806),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_837),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_921),
.A2(n_795),
.B(n_791),
.C(n_793),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_795),
.A2(n_775),
.B1(n_873),
.B2(n_875),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_816),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_951),
.B(n_834),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_965),
.B(n_938),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_948),
.A2(n_832),
.B1(n_879),
.B2(n_775),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1002),
.A2(n_796),
.B(n_877),
.Y(n_1080)
);

O2A1O1Ixp5_ASAP7_75t_SL g1081 ( 
.A1(n_1072),
.A2(n_796),
.B(n_930),
.C(n_929),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_939),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1042),
.B(n_917),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_SL g1084 ( 
.A(n_974),
.B(n_914),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1066),
.A2(n_932),
.B(n_850),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1005),
.A2(n_845),
.B(n_862),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1075),
.A2(n_850),
.B(n_853),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_951),
.B(n_836),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_974),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_973),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_977),
.A2(n_1056),
.B(n_1061),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1067),
.B(n_759),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1026),
.A2(n_1012),
.B(n_944),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_982),
.A2(n_917),
.B(n_907),
.C(n_803),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_962),
.A2(n_853),
.B(n_858),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_941),
.A2(n_858),
.B(n_863),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1037),
.B(n_871),
.C(n_934),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_976),
.A2(n_930),
.B(n_929),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1011),
.A2(n_868),
.A3(n_937),
.B(n_927),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_957),
.A2(n_926),
.B(n_914),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_981),
.A2(n_832),
.B1(n_879),
.B2(n_759),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_994),
.A2(n_954),
.B(n_960),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_952),
.A2(n_765),
.B(n_767),
.C(n_935),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1003),
.A2(n_876),
.B(n_777),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_949),
.B(n_825),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1034),
.B(n_923),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_942),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1058),
.B(n_923),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_857),
.B(n_799),
.C(n_800),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_991),
.A2(n_777),
.B(n_904),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_975),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1051),
.A2(n_914),
.B(n_923),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_955),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_961),
.B(n_964),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1006),
.A2(n_825),
.B(n_788),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_966),
.B(n_799),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_959),
.B(n_933),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1074),
.A2(n_884),
.B(n_916),
.C(n_913),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1007),
.A2(n_788),
.B(n_838),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1029),
.B(n_844),
.C(n_904),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1000),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_958),
.A2(n_924),
.B(n_857),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_970),
.A2(n_874),
.B(n_816),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_945),
.A2(n_772),
.B(n_924),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_986),
.B(n_800),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1044),
.A2(n_1047),
.B1(n_963),
.B2(n_1030),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_940),
.A2(n_874),
.B(n_816),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1001),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1031),
.B(n_870),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_947),
.Y(n_1130)
);

OAI22x1_ASAP7_75t_L g1131 ( 
.A1(n_1032),
.A2(n_919),
.B1(n_906),
.B2(n_901),
.Y(n_1131)
);

AOI211x1_ASAP7_75t_L g1132 ( 
.A1(n_1033),
.A2(n_772),
.B(n_844),
.C(n_934),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1065),
.B(n_892),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_998),
.A2(n_772),
.B(n_842),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_998),
.A2(n_890),
.B(n_865),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1040),
.A2(n_772),
.A3(n_842),
.B(n_835),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1038),
.A2(n_842),
.B(n_838),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1068),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1004),
.A2(n_835),
.B(n_838),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_979),
.B(n_874),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_997),
.A2(n_835),
.B(n_838),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_990),
.A2(n_1053),
.B(n_1050),
.C(n_1062),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_1036),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1046),
.A2(n_1008),
.B(n_1015),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1063),
.A2(n_1060),
.B(n_1039),
.C(n_1071),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_996),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1028),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1017),
.A2(n_1041),
.B(n_1020),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1016),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1018),
.A2(n_956),
.B(n_992),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_968),
.B(n_972),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_971),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1069),
.A2(n_999),
.B(n_1018),
.C(n_1070),
.Y(n_1153)
);

OAI22x1_ASAP7_75t_L g1154 ( 
.A1(n_1057),
.A2(n_1055),
.B1(n_1025),
.B2(n_980),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_985),
.B(n_983),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1073),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1010),
.B(n_1014),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1018),
.A2(n_1009),
.B(n_1049),
.C(n_988),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1001),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1048),
.B(n_1043),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1022),
.B(n_1052),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_950),
.B(n_969),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_950),
.B(n_969),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_995),
.B(n_943),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_953),
.B(n_993),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1009),
.A2(n_1047),
.B(n_1044),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1044),
.B(n_1047),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1013),
.A2(n_1021),
.B(n_1023),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1019),
.A2(n_1027),
.B(n_1054),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_987),
.A2(n_989),
.B(n_978),
.C(n_975),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_967),
.A2(n_1076),
.A3(n_1000),
.B(n_946),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_975),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_946),
.A2(n_1064),
.B(n_967),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_967),
.A2(n_946),
.B(n_1064),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1076),
.B(n_1024),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_946),
.B(n_1064),
.Y(n_1176)
);

AND3x4_ASAP7_75t_L g1177 ( 
.A(n_984),
.B(n_1045),
.C(n_1024),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1059),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1064),
.B(n_946),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1059),
.B(n_1064),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1059),
.B(n_629),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_1075),
.A2(n_617),
.B(n_611),
.C(n_614),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_951),
.B(n_621),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_944),
.A2(n_1054),
.B1(n_1075),
.B2(n_1072),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1026),
.A2(n_1066),
.B(n_1011),
.C(n_1017),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1002),
.A2(n_1005),
.B(n_977),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_942),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1031),
.A2(n_322),
.B1(n_330),
.B2(n_320),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1042),
.B(n_629),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_942),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_951),
.B(n_621),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1002),
.A2(n_1005),
.B(n_977),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_951),
.A2(n_1063),
.B(n_1062),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_939),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1002),
.A2(n_1005),
.B(n_977),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_947),
.Y(n_1201)
);

AO21x1_ASAP7_75t_L g1202 ( 
.A1(n_1075),
.A2(n_944),
.B(n_982),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_982),
.A2(n_730),
.B(n_655),
.C(n_621),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_942),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1075),
.A2(n_944),
.A3(n_899),
.B(n_1066),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_951),
.B(n_621),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1031),
.B(n_1048),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_982),
.A2(n_730),
.B(n_655),
.C(n_621),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_959),
.B(n_461),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1066),
.A2(n_903),
.B(n_881),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_993),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_951),
.B(n_621),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1107),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1091),
.A2(n_1144),
.B(n_1123),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1113),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1130),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1203),
.A2(n_1208),
.B1(n_1114),
.B2(n_1164),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1167),
.B(n_1152),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1202),
.A2(n_1184),
.B1(n_1079),
.B2(n_1101),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1167),
.B(n_1166),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1135),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1156),
.B(n_1106),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1078),
.B(n_1130),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1101),
.A2(n_1155),
.B1(n_1192),
.B2(n_1206),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1093),
.A2(n_1182),
.B(n_1102),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1086),
.A2(n_1098),
.B(n_1080),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1096),
.A2(n_1085),
.B(n_1122),
.Y(n_1228)
);

AND2x6_ASAP7_75t_L g1229 ( 
.A(n_1176),
.B(n_1179),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1190),
.B(n_1129),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1108),
.B(n_1083),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1187),
.B(n_1191),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1183),
.A2(n_1212),
.B1(n_1206),
.B2(n_1079),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_1196),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1188),
.A2(n_1195),
.B(n_1210),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1090),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1204),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1151),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1197),
.A2(n_1200),
.B(n_1199),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1142),
.A2(n_1145),
.B(n_1183),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1212),
.A2(n_1134),
.B(n_1124),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1151),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1158),
.A2(n_1094),
.B(n_1153),
.C(n_1124),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1084),
.A2(n_1194),
.B(n_1150),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1157),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_1100),
.A3(n_1095),
.B(n_1087),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1120),
.A2(n_1077),
.B(n_1093),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1104),
.A2(n_1148),
.B(n_1109),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1184),
.A2(n_1177),
.B1(n_1097),
.B2(n_1126),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1189),
.A2(n_1117),
.B1(n_1133),
.B2(n_1088),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1185),
.A2(n_1077),
.B(n_1148),
.Y(n_1251)
);

OAI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1170),
.A2(n_1209),
.B1(n_1165),
.B2(n_1168),
.C(n_1149),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1103),
.A2(n_1081),
.B(n_1088),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1111),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1201),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1134),
.A2(n_1110),
.B1(n_1092),
.B2(n_1132),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1092),
.A2(n_1179),
.B(n_1176),
.C(n_1137),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1137),
.A2(n_1173),
.B(n_1168),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1207),
.B(n_1160),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1140),
.B(n_1181),
.C(n_1160),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1154),
.A2(n_1131),
.B1(n_1207),
.B2(n_1125),
.C(n_1116),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1147),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1112),
.A2(n_1139),
.B(n_1169),
.Y(n_1263)
);

NAND2x1p5_ASAP7_75t_L g1264 ( 
.A(n_1089),
.B(n_1111),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1157),
.B(n_1161),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1211),
.A2(n_1159),
.B1(n_1128),
.B2(n_1082),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1118),
.A2(n_1141),
.B(n_1119),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1211),
.A2(n_1105),
.B1(n_1143),
.B2(n_1089),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1162),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1211),
.B(n_1143),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1172),
.B(n_1178),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1127),
.B(n_1180),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1162),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_R g1274 ( 
.A(n_1146),
.B(n_1138),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1111),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1163),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1111),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1089),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1175),
.A2(n_1121),
.B(n_1099),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1099),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1205),
.A2(n_1136),
.A3(n_1171),
.B(n_1175),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1205),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1121),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1186),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1171),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1171),
.A2(n_1174),
.B(n_1173),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1167),
.B(n_1207),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1107),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1107),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1078),
.B(n_1130),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1101),
.A2(n_435),
.B1(n_770),
.B2(n_1079),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1107),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1114),
.B(n_707),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1166),
.B(n_1018),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1089),
.B(n_1111),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1202),
.A2(n_888),
.B1(n_730),
.B2(n_655),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1166),
.B(n_1018),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1203),
.A2(n_948),
.B1(n_1208),
.B2(n_679),
.Y(n_1304)
);

AND2x2_ASAP7_75t_SL g1305 ( 
.A(n_1167),
.B(n_948),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1107),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1307)
);

OAI221xp5_ASAP7_75t_L g1308 ( 
.A1(n_1203),
.A2(n_435),
.B1(n_1208),
.B2(n_655),
.C(n_732),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1196),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1310)
);

XNOR2xp5_ASAP7_75t_L g1311 ( 
.A(n_1189),
.B(n_489),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1167),
.B(n_1044),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1166),
.B(n_1018),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1090),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1090),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1088),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1211),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1138),
.B(n_461),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1203),
.A2(n_1208),
.B(n_1101),
.C(n_730),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1089),
.B(n_1111),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1196),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1107),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1089),
.B(n_1111),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1203),
.A2(n_1208),
.B(n_1101),
.C(n_730),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1130),
.Y(n_1333)
);

BUFx8_ASAP7_75t_L g1334 ( 
.A(n_1147),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1138),
.B(n_461),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1211),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1167),
.B(n_1044),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1078),
.B(n_1130),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1186),
.A2(n_1198),
.B(n_1193),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1202),
.A2(n_1208),
.A3(n_1203),
.B(n_1174),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1304),
.A2(n_1332),
.B(n_1326),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1230),
.B(n_1231),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1301),
.A2(n_1249),
.B1(n_1308),
.B2(n_1305),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1326),
.A2(n_1332),
.B(n_1240),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1292),
.A2(n_1218),
.B(n_1301),
.C(n_1252),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1235),
.A2(n_1239),
.B(n_1251),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1223),
.B(n_1305),
.Y(n_1347)
);

AND2x6_ASAP7_75t_L g1348 ( 
.A(n_1221),
.B(n_1282),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1217),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1281),
.Y(n_1350)
);

CKINVDCx12_ASAP7_75t_R g1351 ( 
.A(n_1274),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1254),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1249),
.A2(n_1292),
.B1(n_1220),
.B2(n_1250),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1216),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_L g1355 ( 
.A(n_1224),
.B(n_1291),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1260),
.A2(n_1338),
.B1(n_1337),
.B2(n_1316),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1316),
.A2(n_1337),
.B1(n_1219),
.B2(n_1333),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1323),
.B(n_1247),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1264),
.A2(n_1331),
.B(n_1298),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1288),
.B(n_1259),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1271),
.B(n_1232),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1225),
.B(n_1251),
.C(n_1233),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1235),
.A2(n_1239),
.B(n_1243),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1269),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1272),
.A2(n_1257),
.B(n_1253),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1264),
.A2(n_1298),
.B(n_1331),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1266),
.A2(n_1261),
.B1(n_1311),
.B2(n_1255),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1237),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1232),
.B(n_1290),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1261),
.A2(n_1244),
.B(n_1241),
.C(n_1268),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1236),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1238),
.A2(n_1257),
.B(n_1272),
.C(n_1293),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1242),
.B(n_1245),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1266),
.A2(n_1256),
.B1(n_1321),
.B2(n_1322),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1256),
.A2(n_1336),
.B1(n_1324),
.B2(n_1270),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1213),
.B(n_1289),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1324),
.A2(n_1336),
.B1(n_1270),
.B2(n_1296),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1273),
.B(n_1276),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1281),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1327),
.A2(n_1254),
.B(n_1275),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1267),
.A2(n_1296),
.B(n_1318),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1330),
.B(n_1306),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1265),
.B(n_1284),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1284),
.B(n_1234),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1229),
.B(n_1325),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1277),
.B(n_1309),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1309),
.B(n_1329),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1303),
.A2(n_1318),
.B(n_1283),
.C(n_1335),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1229),
.B(n_1329),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_SL g1390 ( 
.A1(n_1280),
.A2(n_1222),
.B(n_1286),
.C(n_1340),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1340),
.B(n_1226),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1303),
.A2(n_1267),
.B(n_1226),
.C(n_1327),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1267),
.A2(n_1226),
.B(n_1263),
.C(n_1248),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1254),
.A2(n_1275),
.B1(n_1278),
.B2(n_1262),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1340),
.B(n_1246),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1275),
.A2(n_1278),
.B1(n_1262),
.B2(n_1258),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1229),
.B(n_1340),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1215),
.A2(n_1339),
.B(n_1214),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1229),
.B(n_1246),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1258),
.A2(n_1248),
.B1(n_1263),
.B2(n_1286),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1246),
.B(n_1229),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1263),
.Y(n_1402)
);

NOR2xp67_ASAP7_75t_L g1403 ( 
.A(n_1287),
.B(n_1334),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1246),
.B(n_1258),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1248),
.B(n_1228),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1285),
.B(n_1227),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1294),
.A2(n_1297),
.B(n_1299),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1334),
.A2(n_1300),
.B1(n_1302),
.B2(n_1307),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1310),
.A2(n_1312),
.B(n_1313),
.C(n_1314),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1315),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1317),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1319),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1320),
.A2(n_1292),
.B(n_1203),
.C(n_1208),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1328),
.B(n_1230),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1235),
.A2(n_1208),
.B(n_1203),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1301),
.A2(n_1208),
.B(n_1203),
.C(n_1251),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1279),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1235),
.A2(n_1208),
.B(n_1203),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1301),
.A2(n_948),
.B1(n_1249),
.B2(n_1177),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1218),
.B(n_1295),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1253),
.A2(n_1239),
.B(n_1235),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1301),
.A2(n_948),
.B1(n_1249),
.B2(n_1177),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1224),
.B(n_1291),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1253),
.A2(n_1239),
.B(n_1235),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1345),
.A2(n_1416),
.B(n_1415),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1358),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1401),
.B(n_1391),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1346),
.A2(n_1363),
.B(n_1418),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1417),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1402),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1393),
.A2(n_1398),
.B(n_1407),
.Y(n_1431)
);

BUFx2_ASAP7_75t_SL g1432 ( 
.A(n_1403),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1350),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1391),
.B(n_1397),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_SL g1436 ( 
.A(n_1343),
.B(n_1419),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1350),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1399),
.B(n_1395),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1354),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1404),
.B(n_1400),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1344),
.B(n_1341),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1358),
.B(n_1414),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1379),
.B(n_1405),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1368),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1365),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1341),
.B(n_1392),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1411),
.Y(n_1450)
);

NAND2x1_ASAP7_75t_L g1451 ( 
.A(n_1348),
.B(n_1344),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1408),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1376),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1390),
.B(n_1410),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1355),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1390),
.B(n_1410),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1388),
.B(n_1370),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1412),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1372),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1412),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1382),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1369),
.B(n_1413),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1373),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1378),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1364),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1430),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1442),
.B(n_1389),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1429),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1430),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1436),
.A2(n_1422),
.B1(n_1353),
.B2(n_1367),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1451),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

AOI211xp5_ASAP7_75t_L g1473 ( 
.A1(n_1425),
.A2(n_1374),
.B(n_1420),
.C(n_1362),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1426),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1437),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1436),
.B(n_1385),
.Y(n_1476)
);

OAI222xp33_ASAP7_75t_L g1477 ( 
.A1(n_1457),
.A2(n_1356),
.B1(n_1347),
.B2(n_1357),
.C1(n_1375),
.C2(n_1361),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1455),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1427),
.B(n_1383),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1442),
.B(n_1349),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1465),
.Y(n_1481)
);

OAI21xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1443),
.A2(n_1366),
.B(n_1359),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1426),
.B(n_1396),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1425),
.B(n_1371),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1342),
.Y(n_1485)
);

NOR2x1_ASAP7_75t_L g1486 ( 
.A(n_1443),
.B(n_1366),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1434),
.B(n_1409),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1462),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1457),
.A2(n_1384),
.B1(n_1386),
.B2(n_1360),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1455),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1471),
.B(n_1447),
.Y(n_1491)
);

NAND4xp75_ASAP7_75t_L g1492 ( 
.A(n_1486),
.B(n_1459),
.C(n_1387),
.D(n_1435),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1478),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1480),
.B(n_1444),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1470),
.A2(n_1457),
.B1(n_1449),
.B2(n_1451),
.C(n_1452),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1475),
.Y(n_1496)
);

AO31x2_ASAP7_75t_L g1497 ( 
.A1(n_1468),
.A2(n_1433),
.A3(n_1460),
.B(n_1450),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1473),
.B(n_1457),
.C(n_1453),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1481),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1488),
.B(n_1474),
.Y(n_1501)
);

OAI332xp33_ASAP7_75t_L g1502 ( 
.A1(n_1484),
.A2(n_1459),
.A3(n_1464),
.B1(n_1458),
.B2(n_1445),
.B3(n_1463),
.C1(n_1456),
.C2(n_1454),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1481),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1457),
.C(n_1453),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1485),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1484),
.A2(n_1457),
.B1(n_1449),
.B2(n_1452),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1447),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1465),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1470),
.A2(n_1462),
.B1(n_1444),
.B2(n_1446),
.C(n_1461),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1490),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1486),
.B(n_1449),
.C(n_1462),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1469),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_R g1513 ( 
.A(n_1476),
.B(n_1449),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1488),
.A2(n_1431),
.B(n_1439),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1469),
.Y(n_1515)
);

AOI21xp33_ASAP7_75t_L g1516 ( 
.A1(n_1482),
.A2(n_1449),
.B(n_1451),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1472),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1489),
.A2(n_1449),
.B1(n_1476),
.B2(n_1485),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1467),
.B(n_1444),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1490),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1482),
.A2(n_1428),
.B(n_1359),
.Y(n_1521)
);

NOR2x1_ASAP7_75t_L g1522 ( 
.A(n_1467),
.B(n_1458),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1471),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1479),
.B(n_1440),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1485),
.Y(n_1525)
);

OAI211xp5_ASAP7_75t_L g1526 ( 
.A1(n_1489),
.A2(n_1448),
.B(n_1438),
.C(n_1439),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1521),
.A2(n_1439),
.B(n_1438),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_L g1528 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1471),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1497),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1517),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1487),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1496),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1500),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1500),
.Y(n_1538)
);

INVx4_ASAP7_75t_SL g1539 ( 
.A(n_1497),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_SL g1540 ( 
.A(n_1492),
.B(n_1471),
.Y(n_1540)
);

OAI31xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1498),
.A2(n_1487),
.A3(n_1377),
.B(n_1394),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1523),
.B(n_1471),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1468),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1504),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1497),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1516),
.A2(n_1438),
.B(n_1515),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1533),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1530),
.B(n_1519),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1523),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1543),
.Y(n_1553)
);

INVx4_ASAP7_75t_SL g1554 ( 
.A(n_1529),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1528),
.B(n_1491),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1549),
.B(n_1491),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1547),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1547),
.B(n_1508),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1549),
.B(n_1507),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_L g1560 ( 
.A(n_1534),
.B(n_1502),
.C(n_1495),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1546),
.B(n_1471),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1541),
.B(n_1506),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1531),
.B(n_1505),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1530),
.B(n_1525),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1543),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1546),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1549),
.B(n_1539),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1549),
.B(n_1514),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1499),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1536),
.B(n_1509),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1529),
.A2(n_1518),
.B1(n_1428),
.B2(n_1471),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1530),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1549),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1535),
.B(n_1494),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1510),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1535),
.B(n_1524),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1537),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1520),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1549),
.B(n_1514),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1537),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1544),
.B(n_1512),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1542),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1527),
.B(n_1483),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1550),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1553),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1541),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1550),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1554),
.B(n_1545),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1557),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1571),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1546),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1571),
.Y(n_1601)
);

OAI32xp33_ASAP7_75t_L g1602 ( 
.A1(n_1564),
.A2(n_1513),
.A3(n_1543),
.B1(n_1503),
.B2(n_1540),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1557),
.B(n_1558),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1558),
.B(n_1576),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1576),
.B(n_1527),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1581),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1568),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_1546),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.B(n_1527),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1527),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1554),
.B(n_1546),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1553),
.B(n_1544),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1579),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1567),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1554),
.B(n_1493),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1527),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1562),
.B(n_1563),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1526),
.C(n_1477),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1562),
.B(n_1546),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1581),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1551),
.B(n_1527),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1563),
.B(n_1546),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1613),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1583),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1617),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1615),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1620),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1598),
.A2(n_1575),
.B1(n_1573),
.B2(n_1529),
.C(n_1577),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1606),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1621),
.A2(n_1529),
.B1(n_1555),
.B2(n_1565),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1574),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1618),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1620),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1592),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1612),
.B(n_1555),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1592),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1623),
.B(n_1574),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1595),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1595),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1578),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1596),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1616),
.A2(n_1529),
.B1(n_1555),
.B2(n_1565),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1624),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1624),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1641),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1632),
.B(n_1622),
.Y(n_1653)
);

AOI21xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1638),
.A2(n_1602),
.B(n_1604),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1604),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1643),
.Y(n_1656)
);

OA21x2_ASAP7_75t_SL g1657 ( 
.A1(n_1631),
.A2(n_1614),
.B(n_1612),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1633),
.A2(n_1602),
.B(n_1577),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1636),
.A2(n_1529),
.B1(n_1597),
.B2(n_1614),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1629),
.A2(n_1529),
.B1(n_1597),
.B2(n_1614),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1643),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1627),
.B(n_1600),
.Y(n_1662)
);

OAI322xp33_ASAP7_75t_L g1663 ( 
.A1(n_1630),
.A2(n_1588),
.A3(n_1609),
.B1(n_1610),
.B2(n_1605),
.C1(n_1619),
.C2(n_1625),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1629),
.A2(n_1552),
.B(n_1611),
.C(n_1608),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1628),
.A2(n_1601),
.B1(n_1599),
.B2(n_1600),
.C(n_1608),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1637),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1582),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1648),
.A2(n_1552),
.B(n_1611),
.C(n_1569),
.Y(n_1668)
);

O2A1O1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1650),
.B(n_1651),
.C(n_1634),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1641),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1639),
.A2(n_1646),
.B1(n_1637),
.B2(n_1651),
.C(n_1634),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1666),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1666),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1662),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1658),
.A2(n_1639),
.B1(n_1641),
.B2(n_1645),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1662),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1670),
.B(n_1647),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1656),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1661),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1653),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1659),
.A2(n_1540),
.B1(n_1622),
.B2(n_1626),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1654),
.C(n_1669),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1652),
.B1(n_1667),
.B2(n_1665),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_L g1684 ( 
.A(n_1676),
.B(n_1655),
.Y(n_1684)
);

NAND4xp25_ASAP7_75t_L g1685 ( 
.A(n_1677),
.B(n_1657),
.C(n_1671),
.D(n_1664),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_L g1686 ( 
.A(n_1672),
.B(n_1668),
.C(n_1660),
.Y(n_1686)
);

O2A1O1Ixp5_ASAP7_75t_L g1687 ( 
.A1(n_1676),
.A2(n_1663),
.B(n_1607),
.C(n_1596),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1673),
.A2(n_1644),
.B1(n_1642),
.B2(n_1640),
.C(n_1646),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1680),
.B(n_1626),
.C(n_1607),
.D(n_1612),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1674),
.B(n_1552),
.C(n_1556),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_L g1691 ( 
.A1(n_1682),
.A2(n_1683),
.B(n_1685),
.C(n_1684),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1687),
.A2(n_1679),
.B(n_1678),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1689),
.B(n_1568),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1688),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1686),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1690),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1693),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1694),
.B(n_1681),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1692),
.B(n_1579),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1691),
.B(n_1568),
.C(n_1569),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1693),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1696),
.A2(n_1568),
.B1(n_1561),
.B2(n_1609),
.C(n_1610),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1701),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1699),
.B(n_1582),
.Y(n_1704)
);

OAI322xp33_ASAP7_75t_L g1705 ( 
.A1(n_1698),
.A2(n_1605),
.A3(n_1619),
.B1(n_1625),
.B2(n_1568),
.C1(n_1588),
.C2(n_1569),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1697),
.B(n_1586),
.Y(n_1706)
);

NOR3xp33_ASAP7_75t_L g1707 ( 
.A(n_1703),
.B(n_1700),
.C(n_1351),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1704),
.B(n_1586),
.Y(n_1708)
);

AO22x2_ASAP7_75t_L g1709 ( 
.A1(n_1706),
.A2(n_1570),
.B1(n_1584),
.B2(n_1591),
.Y(n_1709)
);

NAND4xp75_ASAP7_75t_L g1710 ( 
.A(n_1708),
.B(n_1705),
.C(n_1702),
.D(n_1570),
.Y(n_1710)
);

AOI222xp33_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1709),
.B1(n_1707),
.B2(n_1570),
.C1(n_1584),
.C2(n_1556),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1493),
.B(n_1587),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1712),
.Y(n_1713)
);

OAI22x1_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1561),
.B1(n_1559),
.B2(n_1556),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1546),
.Y(n_1715)
);

OAI222xp33_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1561),
.B1(n_1587),
.B2(n_1590),
.C1(n_1591),
.C2(n_1584),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1351),
.B1(n_1590),
.B2(n_1591),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1716),
.A2(n_1561),
.B1(n_1559),
.B2(n_1540),
.Y(n_1718)
);

AOI31xp67_ASAP7_75t_L g1719 ( 
.A1(n_1717),
.A2(n_1590),
.A3(n_1587),
.B(n_1586),
.Y(n_1719)
);

AOI22x1_ASAP7_75t_L g1720 ( 
.A1(n_1718),
.A2(n_1589),
.B1(n_1585),
.B2(n_1559),
.Y(n_1720)
);

OA22x2_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1589),
.B1(n_1585),
.B2(n_1586),
.Y(n_1721)
);

AOI22x1_ASAP7_75t_L g1722 ( 
.A1(n_1719),
.A2(n_1432),
.B1(n_1578),
.B2(n_1352),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1721),
.A2(n_1722),
.B1(n_1544),
.B2(n_1532),
.C(n_1548),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1380),
.B(n_1544),
.C(n_1352),
.Y(n_1724)
);


endmodule